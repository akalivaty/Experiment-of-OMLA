

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585;

  XNOR2_X1 U322 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U323 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U324 ( .A(n429), .B(KEYINPUT48), .ZN(n430) );
  XNOR2_X1 U325 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U326 ( .A(n431), .B(n430), .ZN(n536) );
  XNOR2_X1 U327 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U328 ( .A(n395), .B(n394), .ZN(n424) );
  XNOR2_X1 U329 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U330 ( .A(n459), .B(G176GAT), .ZN(n460) );
  XNOR2_X1 U331 ( .A(n461), .B(n460), .ZN(G1349GAT) );
  XOR2_X1 U332 ( .A(KEYINPUT0), .B(KEYINPUT83), .Z(n291) );
  XNOR2_X1 U333 ( .A(KEYINPUT82), .B(G127GAT), .ZN(n290) );
  XNOR2_X1 U334 ( .A(n291), .B(n290), .ZN(n292) );
  XOR2_X1 U335 ( .A(G113GAT), .B(n292), .Z(n310) );
  XOR2_X1 U336 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n294) );
  XNOR2_X1 U337 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n293) );
  XNOR2_X1 U338 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U339 ( .A(G169GAT), .B(n295), .Z(n338) );
  XNOR2_X1 U340 ( .A(n310), .B(n338), .ZN(n306) );
  XOR2_X1 U341 ( .A(G43GAT), .B(G134GAT), .Z(n408) );
  XOR2_X1 U342 ( .A(KEYINPUT84), .B(KEYINPUT20), .Z(n297) );
  XNOR2_X1 U343 ( .A(G190GAT), .B(KEYINPUT85), .ZN(n296) );
  XNOR2_X1 U344 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U345 ( .A(n408), .B(n298), .Z(n300) );
  NAND2_X1 U346 ( .A1(G227GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U347 ( .A(n300), .B(n299), .ZN(n302) );
  XNOR2_X1 U348 ( .A(G99GAT), .B(G71GAT), .ZN(n301) );
  XNOR2_X1 U349 ( .A(n301), .B(G120GAT), .ZN(n388) );
  XOR2_X1 U350 ( .A(n302), .B(n388), .Z(n304) );
  XNOR2_X1 U351 ( .A(G15GAT), .B(G176GAT), .ZN(n303) );
  XNOR2_X1 U352 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U353 ( .A(n306), .B(n305), .ZN(n467) );
  XNOR2_X1 U354 ( .A(G148GAT), .B(G85GAT), .ZN(n307) );
  XNOR2_X1 U355 ( .A(n307), .B(G57GAT), .ZN(n387) );
  XOR2_X1 U356 ( .A(G29GAT), .B(KEYINPUT75), .Z(n403) );
  XOR2_X1 U357 ( .A(n387), .B(n403), .Z(n309) );
  NAND2_X1 U358 ( .A1(G225GAT), .A2(G233GAT), .ZN(n308) );
  XNOR2_X1 U359 ( .A(n309), .B(n308), .ZN(n312) );
  INV_X1 U360 ( .A(n310), .ZN(n311) );
  XNOR2_X1 U361 ( .A(n312), .B(n311), .ZN(n329) );
  XOR2_X1 U362 ( .A(KEYINPUT4), .B(KEYINPUT94), .Z(n314) );
  XNOR2_X1 U363 ( .A(KEYINPUT96), .B(KEYINPUT1), .ZN(n313) );
  XNOR2_X1 U364 ( .A(n314), .B(n313), .ZN(n318) );
  XOR2_X1 U365 ( .A(KEYINPUT5), .B(G162GAT), .Z(n316) );
  XNOR2_X1 U366 ( .A(G120GAT), .B(G134GAT), .ZN(n315) );
  XNOR2_X1 U367 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U368 ( .A(n318), .B(n317), .Z(n327) );
  XNOR2_X1 U369 ( .A(KEYINPUT90), .B(KEYINPUT91), .ZN(n319) );
  XNOR2_X1 U370 ( .A(n319), .B(KEYINPUT2), .ZN(n320) );
  XOR2_X1 U371 ( .A(n320), .B(KEYINPUT3), .Z(n322) );
  XNOR2_X1 U372 ( .A(G141GAT), .B(G155GAT), .ZN(n321) );
  XNOR2_X1 U373 ( .A(n322), .B(n321), .ZN(n449) );
  XOR2_X1 U374 ( .A(KEYINPUT95), .B(KEYINPUT6), .Z(n324) );
  XNOR2_X1 U375 ( .A(G1GAT), .B(KEYINPUT93), .ZN(n323) );
  XNOR2_X1 U376 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U377 ( .A(n449), .B(n325), .ZN(n326) );
  XNOR2_X1 U378 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U379 ( .A(n329), .B(n328), .ZN(n476) );
  XNOR2_X1 U380 ( .A(KEYINPUT97), .B(n476), .ZN(n524) );
  XOR2_X1 U381 ( .A(G36GAT), .B(G190GAT), .Z(n404) );
  XOR2_X1 U382 ( .A(G64GAT), .B(G92GAT), .Z(n331) );
  XNOR2_X1 U383 ( .A(G176GAT), .B(G204GAT), .ZN(n330) );
  XNOR2_X1 U384 ( .A(n331), .B(n330), .ZN(n380) );
  XOR2_X1 U385 ( .A(n404), .B(n380), .Z(n333) );
  NAND2_X1 U386 ( .A1(G226GAT), .A2(G233GAT), .ZN(n332) );
  XNOR2_X1 U387 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U388 ( .A(n334), .B(KEYINPUT99), .Z(n336) );
  XOR2_X1 U389 ( .A(G8GAT), .B(KEYINPUT77), .Z(n345) );
  XNOR2_X1 U390 ( .A(n345), .B(KEYINPUT98), .ZN(n335) );
  XNOR2_X1 U391 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U392 ( .A(n338), .B(n337), .ZN(n343) );
  XOR2_X1 U393 ( .A(KEYINPUT89), .B(KEYINPUT21), .Z(n340) );
  XNOR2_X1 U394 ( .A(G197GAT), .B(G211GAT), .ZN(n339) );
  XNOR2_X1 U395 ( .A(n340), .B(n339), .ZN(n342) );
  XOR2_X1 U396 ( .A(G218GAT), .B(KEYINPUT88), .Z(n341) );
  XNOR2_X1 U397 ( .A(n342), .B(n341), .ZN(n452) );
  XNOR2_X1 U398 ( .A(n343), .B(n452), .ZN(n527) );
  XNOR2_X1 U399 ( .A(n527), .B(KEYINPUT122), .ZN(n432) );
  XNOR2_X1 U400 ( .A(G22GAT), .B(G15GAT), .ZN(n344) );
  XNOR2_X1 U401 ( .A(n344), .B(G1GAT), .ZN(n366) );
  XOR2_X1 U402 ( .A(n366), .B(n345), .Z(n347) );
  NAND2_X1 U403 ( .A1(G231GAT), .A2(G233GAT), .ZN(n346) );
  XNOR2_X1 U404 ( .A(n347), .B(n346), .ZN(n363) );
  XOR2_X1 U405 ( .A(KEYINPUT15), .B(KEYINPUT79), .Z(n349) );
  XNOR2_X1 U406 ( .A(G64GAT), .B(KEYINPUT80), .ZN(n348) );
  XNOR2_X1 U407 ( .A(n349), .B(n348), .ZN(n361) );
  XOR2_X1 U408 ( .A(G78GAT), .B(G155GAT), .Z(n351) );
  XNOR2_X1 U409 ( .A(G127GAT), .B(G211GAT), .ZN(n350) );
  XNOR2_X1 U410 ( .A(n351), .B(n350), .ZN(n359) );
  XOR2_X1 U411 ( .A(KEYINPUT78), .B(KEYINPUT81), .Z(n353) );
  XNOR2_X1 U412 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(n352) );
  XNOR2_X1 U413 ( .A(n353), .B(n352), .ZN(n357) );
  XOR2_X1 U414 ( .A(KEYINPUT13), .B(G57GAT), .Z(n355) );
  XNOR2_X1 U415 ( .A(G183GAT), .B(G71GAT), .ZN(n354) );
  XNOR2_X1 U416 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U417 ( .A(n357), .B(n356), .Z(n358) );
  XNOR2_X1 U418 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U419 ( .A(n361), .B(n360), .Z(n362) );
  XNOR2_X1 U420 ( .A(n363), .B(n362), .ZN(n565) );
  XOR2_X1 U421 ( .A(G141GAT), .B(G197GAT), .Z(n365) );
  XNOR2_X1 U422 ( .A(G50GAT), .B(G29GAT), .ZN(n364) );
  XNOR2_X1 U423 ( .A(n365), .B(n364), .ZN(n379) );
  XOR2_X1 U424 ( .A(n366), .B(G36GAT), .Z(n368) );
  XOR2_X1 U425 ( .A(KEYINPUT8), .B(KEYINPUT7), .Z(n416) );
  XNOR2_X1 U426 ( .A(G43GAT), .B(n416), .ZN(n367) );
  XNOR2_X1 U427 ( .A(n368), .B(n367), .ZN(n372) );
  XOR2_X1 U428 ( .A(KEYINPUT67), .B(KEYINPUT30), .Z(n370) );
  NAND2_X1 U429 ( .A1(G229GAT), .A2(G233GAT), .ZN(n369) );
  XNOR2_X1 U430 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U431 ( .A(n372), .B(n371), .Z(n377) );
  XOR2_X1 U432 ( .A(KEYINPUT68), .B(G8GAT), .Z(n374) );
  XNOR2_X1 U433 ( .A(G169GAT), .B(G113GAT), .ZN(n373) );
  XNOR2_X1 U434 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U435 ( .A(n375), .B(KEYINPUT29), .ZN(n376) );
  XNOR2_X1 U436 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U437 ( .A(n379), .B(n378), .Z(n573) );
  XNOR2_X1 U438 ( .A(n380), .B(KEYINPUT73), .ZN(n382) );
  XOR2_X1 U439 ( .A(G106GAT), .B(G78GAT), .Z(n445) );
  XOR2_X1 U440 ( .A(n445), .B(KEYINPUT70), .Z(n381) );
  XNOR2_X1 U441 ( .A(n382), .B(n381), .ZN(n386) );
  XOR2_X1 U442 ( .A(KEYINPUT31), .B(KEYINPUT13), .Z(n384) );
  NAND2_X1 U443 ( .A1(G230GAT), .A2(G233GAT), .ZN(n383) );
  XOR2_X1 U444 ( .A(n384), .B(n383), .Z(n385) );
  XNOR2_X1 U445 ( .A(n386), .B(n385), .ZN(n395) );
  XNOR2_X1 U446 ( .A(n388), .B(n387), .ZN(n393) );
  XOR2_X1 U447 ( .A(KEYINPUT33), .B(KEYINPUT71), .Z(n390) );
  XNOR2_X1 U448 ( .A(KEYINPUT69), .B(KEYINPUT32), .ZN(n389) );
  XNOR2_X1 U449 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U450 ( .A(n391), .B(KEYINPUT72), .ZN(n392) );
  NAND2_X1 U451 ( .A1(n424), .A2(KEYINPUT65), .ZN(n397) );
  OR2_X1 U452 ( .A1(n424), .A2(KEYINPUT65), .ZN(n396) );
  NAND2_X1 U453 ( .A1(n397), .A2(n396), .ZN(n398) );
  XNOR2_X1 U454 ( .A(n398), .B(KEYINPUT41), .ZN(n555) );
  NOR2_X1 U455 ( .A1(n573), .A2(n555), .ZN(n399) );
  XNOR2_X1 U456 ( .A(n399), .B(KEYINPUT46), .ZN(n400) );
  NOR2_X1 U457 ( .A1(n565), .A2(n400), .ZN(n421) );
  XOR2_X1 U458 ( .A(KEYINPUT66), .B(KEYINPUT76), .Z(n402) );
  XNOR2_X1 U459 ( .A(G106GAT), .B(KEYINPUT9), .ZN(n401) );
  XNOR2_X1 U460 ( .A(n402), .B(n401), .ZN(n420) );
  XOR2_X1 U461 ( .A(n404), .B(n403), .Z(n406) );
  XNOR2_X1 U462 ( .A(G99GAT), .B(G218GAT), .ZN(n405) );
  XNOR2_X1 U463 ( .A(n406), .B(n405), .ZN(n412) );
  XNOR2_X1 U464 ( .A(G50GAT), .B(KEYINPUT74), .ZN(n407) );
  XNOR2_X1 U465 ( .A(n407), .B(G162GAT), .ZN(n444) );
  XOR2_X1 U466 ( .A(n444), .B(n408), .Z(n410) );
  NAND2_X1 U467 ( .A1(G232GAT), .A2(G233GAT), .ZN(n409) );
  XNOR2_X1 U468 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U469 ( .A(n412), .B(n411), .Z(n418) );
  XOR2_X1 U470 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n414) );
  XNOR2_X1 U471 ( .A(G85GAT), .B(G92GAT), .ZN(n413) );
  XNOR2_X1 U472 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U473 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U474 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U475 ( .A(n420), .B(n419), .Z(n462) );
  NAND2_X1 U476 ( .A1(n421), .A2(n462), .ZN(n422) );
  XNOR2_X1 U477 ( .A(n422), .B(KEYINPUT47), .ZN(n428) );
  INV_X1 U478 ( .A(n573), .ZN(n562) );
  XNOR2_X1 U479 ( .A(KEYINPUT36), .B(n462), .ZN(n583) );
  INV_X1 U480 ( .A(n565), .ZN(n580) );
  NOR2_X1 U481 ( .A1(n583), .A2(n580), .ZN(n423) );
  XNOR2_X1 U482 ( .A(KEYINPUT45), .B(n423), .ZN(n425) );
  NAND2_X1 U483 ( .A1(n425), .A2(n424), .ZN(n426) );
  NOR2_X1 U484 ( .A1(n562), .A2(n426), .ZN(n427) );
  NOR2_X1 U485 ( .A1(n428), .A2(n427), .ZN(n431) );
  INV_X1 U486 ( .A(KEYINPUT64), .ZN(n429) );
  AND2_X1 U487 ( .A1(n432), .A2(n536), .ZN(n436) );
  INV_X1 U488 ( .A(KEYINPUT123), .ZN(n434) );
  INV_X1 U489 ( .A(KEYINPUT54), .ZN(n433) );
  NOR2_X1 U490 ( .A1(n524), .A2(n437), .ZN(n572) );
  XOR2_X1 U491 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n439) );
  XNOR2_X1 U492 ( .A(G22GAT), .B(KEYINPUT92), .ZN(n438) );
  XNOR2_X1 U493 ( .A(n439), .B(n438), .ZN(n443) );
  XOR2_X1 U494 ( .A(G148GAT), .B(G204GAT), .Z(n441) );
  XNOR2_X1 U495 ( .A(KEYINPUT22), .B(KEYINPUT87), .ZN(n440) );
  XNOR2_X1 U496 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U497 ( .A(n443), .B(n442), .Z(n451) );
  XOR2_X1 U498 ( .A(n445), .B(n444), .Z(n447) );
  NAND2_X1 U499 ( .A1(G228GAT), .A2(G233GAT), .ZN(n446) );
  XNOR2_X1 U500 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U501 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U502 ( .A(n451), .B(n450), .ZN(n453) );
  XNOR2_X1 U503 ( .A(n453), .B(n452), .ZN(n472) );
  NAND2_X1 U504 ( .A1(n572), .A2(n472), .ZN(n457) );
  XOR2_X1 U505 ( .A(KEYINPUT125), .B(KEYINPUT55), .Z(n455) );
  INV_X1 U506 ( .A(KEYINPUT124), .ZN(n454) );
  NOR2_X1 U507 ( .A1(n467), .A2(n458), .ZN(n568) );
  XNOR2_X1 U508 ( .A(n555), .B(KEYINPUT111), .ZN(n541) );
  NAND2_X1 U509 ( .A1(n568), .A2(n541), .ZN(n461) );
  XOR2_X1 U510 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n459) );
  NAND2_X1 U511 ( .A1(n424), .A2(n562), .ZN(n494) );
  INV_X1 U512 ( .A(n462), .ZN(n567) );
  NOR2_X1 U513 ( .A1(n567), .A2(n580), .ZN(n463) );
  XNOR2_X1 U514 ( .A(n463), .B(KEYINPUT16), .ZN(n481) );
  XNOR2_X1 U515 ( .A(KEYINPUT27), .B(n527), .ZN(n470) );
  NAND2_X1 U516 ( .A1(n470), .A2(n524), .ZN(n464) );
  XOR2_X1 U517 ( .A(KEYINPUT100), .B(n464), .Z(n551) );
  XNOR2_X1 U518 ( .A(n472), .B(KEYINPUT28), .ZN(n488) );
  NAND2_X1 U519 ( .A1(n551), .A2(n488), .ZN(n539) );
  XOR2_X1 U520 ( .A(n467), .B(KEYINPUT86), .Z(n465) );
  NOR2_X1 U521 ( .A1(n539), .A2(n465), .ZN(n466) );
  XNOR2_X1 U522 ( .A(KEYINPUT101), .B(n466), .ZN(n480) );
  INV_X1 U523 ( .A(n467), .ZN(n537) );
  NOR2_X1 U524 ( .A1(n472), .A2(n537), .ZN(n469) );
  XNOR2_X1 U525 ( .A(KEYINPUT102), .B(KEYINPUT26), .ZN(n468) );
  XNOR2_X1 U526 ( .A(n469), .B(n468), .ZN(n571) );
  NAND2_X1 U527 ( .A1(n571), .A2(n470), .ZN(n475) );
  NAND2_X1 U528 ( .A1(n537), .A2(n527), .ZN(n471) );
  NAND2_X1 U529 ( .A1(n472), .A2(n471), .ZN(n473) );
  XOR2_X1 U530 ( .A(KEYINPUT25), .B(n473), .Z(n474) );
  NAND2_X1 U531 ( .A1(n475), .A2(n474), .ZN(n477) );
  NAND2_X1 U532 ( .A1(n477), .A2(n476), .ZN(n478) );
  XOR2_X1 U533 ( .A(KEYINPUT103), .B(n478), .Z(n479) );
  NAND2_X1 U534 ( .A1(n480), .A2(n479), .ZN(n491) );
  NAND2_X1 U535 ( .A1(n481), .A2(n491), .ZN(n509) );
  NOR2_X1 U536 ( .A1(n494), .A2(n509), .ZN(n489) );
  NAND2_X1 U537 ( .A1(n489), .A2(n524), .ZN(n482) );
  XNOR2_X1 U538 ( .A(n482), .B(KEYINPUT34), .ZN(n483) );
  XNOR2_X1 U539 ( .A(G1GAT), .B(n483), .ZN(G1324GAT) );
  NAND2_X1 U540 ( .A1(n527), .A2(n489), .ZN(n484) );
  XNOR2_X1 U541 ( .A(n484), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U542 ( .A(KEYINPUT35), .B(KEYINPUT104), .Z(n486) );
  NAND2_X1 U543 ( .A1(n489), .A2(n537), .ZN(n485) );
  XNOR2_X1 U544 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U545 ( .A(G15GAT), .B(n487), .ZN(G1326GAT) );
  INV_X1 U546 ( .A(n488), .ZN(n530) );
  NAND2_X1 U547 ( .A1(n489), .A2(n530), .ZN(n490) );
  XNOR2_X1 U548 ( .A(n490), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U549 ( .A1(n580), .A2(n491), .ZN(n492) );
  NOR2_X1 U550 ( .A1(n583), .A2(n492), .ZN(n493) );
  XNOR2_X1 U551 ( .A(KEYINPUT37), .B(n493), .ZN(n522) );
  NOR2_X1 U552 ( .A1(n494), .A2(n522), .ZN(n495) );
  XNOR2_X1 U553 ( .A(n495), .B(KEYINPUT38), .ZN(n504) );
  NAND2_X1 U554 ( .A1(n504), .A2(n524), .ZN(n498) );
  XNOR2_X1 U555 ( .A(G29GAT), .B(KEYINPUT105), .ZN(n496) );
  XNOR2_X1 U556 ( .A(n496), .B(KEYINPUT39), .ZN(n497) );
  XNOR2_X1 U557 ( .A(n498), .B(n497), .ZN(G1328GAT) );
  NAND2_X1 U558 ( .A1(n504), .A2(n527), .ZN(n499) );
  XNOR2_X1 U559 ( .A(n499), .B(KEYINPUT106), .ZN(n500) );
  XNOR2_X1 U560 ( .A(G36GAT), .B(n500), .ZN(G1329GAT) );
  XOR2_X1 U561 ( .A(KEYINPUT40), .B(KEYINPUT107), .Z(n502) );
  NAND2_X1 U562 ( .A1(n504), .A2(n537), .ZN(n501) );
  XNOR2_X1 U563 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U564 ( .A(G43GAT), .B(n503), .ZN(G1330GAT) );
  XOR2_X1 U565 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n506) );
  NAND2_X1 U566 ( .A1(n530), .A2(n504), .ZN(n505) );
  XNOR2_X1 U567 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U568 ( .A(G50GAT), .B(n507), .ZN(G1331GAT) );
  XOR2_X1 U569 ( .A(KEYINPUT114), .B(KEYINPUT113), .Z(n511) );
  NAND2_X1 U570 ( .A1(n541), .A2(n573), .ZN(n508) );
  XNOR2_X1 U571 ( .A(n508), .B(KEYINPUT112), .ZN(n523) );
  NOR2_X1 U572 ( .A1(n523), .A2(n509), .ZN(n518) );
  NAND2_X1 U573 ( .A1(n518), .A2(n524), .ZN(n510) );
  XNOR2_X1 U574 ( .A(n511), .B(n510), .ZN(n513) );
  XOR2_X1 U575 ( .A(G57GAT), .B(KEYINPUT42), .Z(n512) );
  XNOR2_X1 U576 ( .A(n513), .B(n512), .ZN(n514) );
  XOR2_X1 U577 ( .A(KEYINPUT110), .B(n514), .Z(G1332GAT) );
  NAND2_X1 U578 ( .A1(n527), .A2(n518), .ZN(n515) );
  XNOR2_X1 U579 ( .A(n515), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U580 ( .A(G71GAT), .B(KEYINPUT115), .Z(n517) );
  NAND2_X1 U581 ( .A1(n518), .A2(n537), .ZN(n516) );
  XNOR2_X1 U582 ( .A(n517), .B(n516), .ZN(G1334GAT) );
  XOR2_X1 U583 ( .A(KEYINPUT43), .B(KEYINPUT116), .Z(n520) );
  NAND2_X1 U584 ( .A1(n518), .A2(n530), .ZN(n519) );
  XNOR2_X1 U585 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U586 ( .A(G78GAT), .B(n521), .ZN(G1335GAT) );
  XOR2_X1 U587 ( .A(G85GAT), .B(KEYINPUT117), .Z(n526) );
  NOR2_X1 U588 ( .A1(n523), .A2(n522), .ZN(n531) );
  NAND2_X1 U589 ( .A1(n531), .A2(n524), .ZN(n525) );
  XNOR2_X1 U590 ( .A(n526), .B(n525), .ZN(G1336GAT) );
  NAND2_X1 U591 ( .A1(n527), .A2(n531), .ZN(n528) );
  XNOR2_X1 U592 ( .A(n528), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U593 ( .A1(n537), .A2(n531), .ZN(n529) );
  XNOR2_X1 U594 ( .A(n529), .B(G99GAT), .ZN(G1338GAT) );
  XNOR2_X1 U595 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n535) );
  XOR2_X1 U596 ( .A(KEYINPUT119), .B(KEYINPUT118), .Z(n533) );
  NAND2_X1 U597 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U598 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U599 ( .A(n535), .B(n534), .ZN(G1339GAT) );
  NAND2_X1 U600 ( .A1(n537), .A2(n536), .ZN(n538) );
  NOR2_X1 U601 ( .A1(n539), .A2(n538), .ZN(n548) );
  NAND2_X1 U602 ( .A1(n562), .A2(n548), .ZN(n540) );
  XNOR2_X1 U603 ( .A(n540), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT120), .B(KEYINPUT49), .Z(n543) );
  NAND2_X1 U605 ( .A1(n548), .A2(n541), .ZN(n542) );
  XNOR2_X1 U606 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U607 ( .A(G120GAT), .B(n544), .ZN(G1341GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT121), .B(KEYINPUT50), .Z(n546) );
  NAND2_X1 U609 ( .A1(n548), .A2(n565), .ZN(n545) );
  XNOR2_X1 U610 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U611 ( .A(G127GAT), .B(n547), .ZN(G1342GAT) );
  XOR2_X1 U612 ( .A(G134GAT), .B(KEYINPUT51), .Z(n550) );
  NAND2_X1 U613 ( .A1(n548), .A2(n567), .ZN(n549) );
  XNOR2_X1 U614 ( .A(n550), .B(n549), .ZN(G1343GAT) );
  AND2_X1 U615 ( .A1(n571), .A2(n551), .ZN(n552) );
  NAND2_X1 U616 ( .A1(n536), .A2(n552), .ZN(n554) );
  INV_X1 U617 ( .A(n554), .ZN(n560) );
  NAND2_X1 U618 ( .A1(n560), .A2(n562), .ZN(n553) );
  XNOR2_X1 U619 ( .A(G141GAT), .B(n553), .ZN(G1344GAT) );
  NOR2_X1 U620 ( .A1(n555), .A2(n554), .ZN(n557) );
  XNOR2_X1 U621 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U623 ( .A(G148GAT), .B(n558), .ZN(G1345GAT) );
  NAND2_X1 U624 ( .A1(n560), .A2(n565), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n559), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U626 ( .A1(n567), .A2(n560), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n561), .B(G162GAT), .ZN(G1347GAT) );
  XNOR2_X1 U628 ( .A(G169GAT), .B(KEYINPUT126), .ZN(n564) );
  NAND2_X1 U629 ( .A1(n568), .A2(n562), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(G1348GAT) );
  NAND2_X1 U631 ( .A1(n568), .A2(n565), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n566), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U633 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n570) );
  NAND2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(G1351GAT) );
  NAND2_X1 U636 ( .A1(n572), .A2(n571), .ZN(n582) );
  NOR2_X1 U637 ( .A1(n582), .A2(n573), .ZN(n577) );
  XOR2_X1 U638 ( .A(KEYINPUT60), .B(KEYINPUT127), .Z(n575) );
  XNOR2_X1 U639 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n577), .B(n576), .ZN(G1352GAT) );
  NOR2_X1 U642 ( .A1(n424), .A2(n582), .ZN(n579) );
  XNOR2_X1 U643 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1353GAT) );
  NOR2_X1 U645 ( .A1(n580), .A2(n582), .ZN(n581) );
  XOR2_X1 U646 ( .A(G211GAT), .B(n581), .Z(G1354GAT) );
  NOR2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U648 ( .A(KEYINPUT62), .B(n584), .Z(n585) );
  XNOR2_X1 U649 ( .A(G218GAT), .B(n585), .ZN(G1355GAT) );
endmodule

