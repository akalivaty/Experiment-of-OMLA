//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 0 1 0 0 1 1 1 1 0 1 0 0 0 1 0 1 1 1 0 1 1 1 0 1 1 1 0 0 1 0 1 0 1 1 0 1 0 1 1 0 0 0 1 1 0 0 0 1 0 1 0 0 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:06 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1274, new_n1275, new_n1276, new_n1277, new_n1278, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  INV_X1    g0003(.A(G97), .ZN(new_n204));
  INV_X1    g0004(.A(G107), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT64), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n202), .A2(G50), .ZN(new_n216));
  XNOR2_X1  g0016(.A(KEYINPUT65), .B(G20), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  OR3_X1    g0018(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n220));
  INV_X1    g0020(.A(G50), .ZN(new_n221));
  INV_X1    g0021(.A(G226), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  XOR2_X1   g0023(.A(KEYINPUT66), .B(G238), .Z(new_n224));
  AOI21_X1  g0024(.A(new_n223), .B1(G68), .B2(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n226), .A2(KEYINPUT67), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n229));
  INV_X1    g0029(.A(KEYINPUT67), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n228), .B(new_n229), .C1(new_n225), .C2(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n211), .B1(new_n227), .B2(new_n231), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n215), .B(new_n219), .C1(KEYINPUT1), .C2(new_n232), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n233), .B1(KEYINPUT1), .B2(new_n232), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G264), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XOR2_X1   g0043(.A(G107), .B(G116), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G68), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  NOR2_X1   g0049(.A1(G20), .A2(G33), .ZN(new_n250));
  INV_X1    g0050(.A(G68), .ZN(new_n251));
  AOI22_X1  g0051(.A1(new_n250), .A2(G50), .B1(G20), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n217), .A2(G33), .ZN(new_n253));
  INV_X1    g0053(.A(G77), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n218), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT11), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n258), .A2(new_n259), .ZN(new_n262));
  INV_X1    g0062(.A(G13), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n263), .A2(G1), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G20), .ZN(new_n265));
  NOR3_X1   g0065(.A1(new_n265), .A2(KEYINPUT12), .A3(G68), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT12), .ZN(new_n267));
  NOR3_X1   g0067(.A1(new_n263), .A2(new_n209), .A3(G1), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n267), .B1(new_n268), .B2(new_n251), .ZN(new_n269));
  INV_X1    g0069(.A(new_n257), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n208), .A2(G20), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  OAI22_X1  g0072(.A1(new_n266), .A2(new_n269), .B1(new_n272), .B2(new_n251), .ZN(new_n273));
  NOR3_X1   g0073(.A1(new_n261), .A2(new_n262), .A3(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G169), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT70), .ZN(new_n277));
  INV_X1    g0077(.A(G1698), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(KEYINPUT70), .A2(G1698), .ZN(new_n280));
  AND2_X1   g0080(.A1(KEYINPUT3), .A2(G33), .ZN(new_n281));
  NOR2_X1   g0081(.A1(KEYINPUT3), .A2(G33), .ZN(new_n282));
  OAI211_X1 g0082(.A(new_n279), .B(new_n280), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G226), .ZN(new_n285));
  OR2_X1    g0085(.A1(KEYINPUT3), .A2(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(KEYINPUT3), .A2(G33), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n278), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  AOI22_X1  g0088(.A1(new_n288), .A2(G232), .B1(G33), .B2(G97), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n285), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n218), .B1(G33), .B2(G41), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT13), .ZN(new_n293));
  INV_X1    g0093(.A(G45), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(KEYINPUT68), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT68), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G45), .ZN(new_n297));
  INV_X1    g0097(.A(G41), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n295), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G274), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n300), .A2(G1), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT69), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n299), .A2(KEYINPUT69), .A3(new_n301), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G33), .ZN(new_n307));
  OAI211_X1 g0107(.A(G1), .B(G13), .C1(new_n307), .C2(new_n298), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(G238), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n292), .A2(new_n293), .A3(new_n306), .A4(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n306), .A2(new_n312), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n308), .B1(new_n285), .B2(new_n289), .ZN(new_n315));
  OAI21_X1  g0115(.A(KEYINPUT13), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n276), .B1(new_n313), .B2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT14), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n313), .A2(new_n316), .ZN(new_n319));
  INV_X1    g0119(.A(G179), .ZN(new_n320));
  OAI22_X1  g0120(.A1(new_n317), .A2(new_n318), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  AND2_X1   g0121(.A1(new_n317), .A2(new_n318), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n275), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n319), .A2(G200), .ZN(new_n324));
  INV_X1    g0124(.A(G190), .ZN(new_n325));
  OAI211_X1 g0125(.A(new_n324), .B(new_n274), .C1(new_n325), .C2(new_n319), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n209), .A2(KEYINPUT65), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT65), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(G20), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(G77), .ZN(new_n331));
  INV_X1    g0131(.A(new_n250), .ZN(new_n332));
  XNOR2_X1  g0132(.A(KEYINPUT8), .B(G58), .ZN(new_n333));
  XNOR2_X1  g0133(.A(KEYINPUT15), .B(G87), .ZN(new_n334));
  OAI221_X1 g0134(.A(new_n331), .B1(new_n332), .B2(new_n333), .C1(new_n253), .C2(new_n334), .ZN(new_n335));
  AND2_X1   g0135(.A1(new_n335), .A2(new_n257), .ZN(new_n336));
  INV_X1    g0136(.A(new_n272), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(G77), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n338), .B1(G77), .B2(new_n265), .ZN(new_n339));
  OR2_X1    g0139(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n311), .A2(G244), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n306), .A2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT74), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n284), .A2(new_n343), .A3(G232), .ZN(new_n344));
  INV_X1    g0144(.A(G232), .ZN(new_n345));
  OAI21_X1  g0145(.A(KEYINPUT74), .B1(new_n283), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT72), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n288), .A2(new_n348), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n348), .B(G1698), .C1(new_n281), .C2(new_n282), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n224), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n281), .A2(new_n282), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(G107), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n347), .A2(new_n352), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n342), .B1(new_n355), .B2(new_n291), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n340), .B1(new_n356), .B2(G190), .ZN(new_n357));
  AOI22_X1  g0157(.A1(new_n344), .A2(new_n346), .B1(G107), .B2(new_n353), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n308), .B1(new_n358), .B2(new_n352), .ZN(new_n359));
  OAI21_X1  g0159(.A(G200), .B1(new_n359), .B2(new_n342), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(KEYINPUT75), .B1(new_n356), .B2(G169), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n356), .A2(new_n320), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n336), .A2(new_n339), .ZN(new_n365));
  AOI211_X1 g0165(.A(G179), .B(new_n342), .C1(new_n355), .C2(new_n291), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n365), .B1(new_n366), .B2(KEYINPUT75), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n323), .A2(new_n326), .A3(new_n361), .A4(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n279), .A2(G223), .A3(new_n280), .ZN(new_n371));
  NAND2_X1  g0171(.A1(G226), .A2(G1698), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n353), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(G87), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n307), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n291), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  AND3_X1   g0176(.A1(new_n308), .A2(G232), .A3(new_n309), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  AND4_X1   g0178(.A1(new_n320), .A2(new_n306), .A3(new_n376), .A4(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n377), .B1(new_n304), .B2(new_n305), .ZN(new_n380));
  AOI21_X1  g0180(.A(G169), .B1(new_n380), .B2(new_n376), .ZN(new_n381));
  OAI21_X1  g0181(.A(KEYINPUT78), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT78), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n380), .A2(new_n320), .A3(new_n376), .ZN(new_n384));
  AND3_X1   g0184(.A1(new_n306), .A2(new_n376), .A3(new_n378), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n383), .B(new_n384), .C1(new_n385), .C2(G169), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n382), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(KEYINPUT73), .A2(G58), .ZN(new_n388));
  XNOR2_X1  g0188(.A(new_n388), .B(KEYINPUT8), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n389), .A2(KEYINPUT77), .A3(new_n271), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n268), .A2(new_n257), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(KEYINPUT77), .B1(new_n389), .B2(new_n271), .ZN(new_n393));
  OAI22_X1  g0193(.A1(new_n392), .A2(new_n393), .B1(new_n265), .B2(new_n389), .ZN(new_n394));
  AND2_X1   g0194(.A1(G58), .A2(G68), .ZN(new_n395));
  OR2_X1    g0195(.A1(new_n395), .A2(new_n201), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n396), .A2(G20), .B1(G159), .B2(new_n250), .ZN(new_n397));
  NOR3_X1   g0197(.A1(new_n281), .A2(new_n282), .A3(G20), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT7), .ZN(new_n399));
  OAI21_X1  g0199(.A(G68), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  AND3_X1   g0200(.A1(new_n353), .A2(new_n217), .A3(new_n399), .ZN(new_n401));
  OAI211_X1 g0201(.A(KEYINPUT16), .B(new_n397), .C1(new_n400), .C2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(KEYINPUT76), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n395), .A2(new_n201), .ZN(new_n404));
  INV_X1    g0204(.A(G159), .ZN(new_n405));
  OAI22_X1  g0205(.A1(new_n404), .A2(new_n209), .B1(new_n405), .B2(new_n332), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n286), .A2(new_n209), .A3(new_n287), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n251), .B1(new_n407), .B2(KEYINPUT7), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n353), .A2(new_n217), .A3(new_n399), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n406), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT76), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n410), .A2(new_n411), .A3(KEYINPUT16), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n403), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n286), .A2(new_n287), .ZN(new_n414));
  OAI21_X1  g0214(.A(KEYINPUT7), .B1(new_n414), .B2(new_n330), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n398), .A2(new_n399), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n397), .B1(new_n417), .B2(new_n251), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT16), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n270), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n394), .B1(new_n413), .B2(new_n420), .ZN(new_n421));
  OAI21_X1  g0221(.A(KEYINPUT18), .B1(new_n387), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n413), .A2(new_n420), .ZN(new_n423));
  INV_X1    g0223(.A(new_n394), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT18), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n425), .A2(new_n426), .A3(new_n382), .A4(new_n386), .ZN(new_n427));
  AND3_X1   g0227(.A1(new_n380), .A2(G190), .A3(new_n376), .ZN(new_n428));
  INV_X1    g0228(.A(G200), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n429), .B1(new_n380), .B2(new_n376), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n423), .A2(new_n431), .A3(new_n424), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT17), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n421), .A2(KEYINPUT17), .A3(new_n431), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n422), .A2(new_n427), .A3(new_n434), .A4(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT79), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n284), .A2(KEYINPUT71), .A3(G222), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT71), .ZN(new_n440));
  INV_X1    g0240(.A(G222), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n440), .B1(new_n283), .B2(new_n441), .ZN(new_n442));
  AOI22_X1  g0242(.A1(new_n439), .A2(new_n442), .B1(G77), .B2(new_n353), .ZN(new_n443));
  OAI21_X1  g0243(.A(G223), .B1(new_n349), .B2(new_n351), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n308), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n306), .B1(new_n222), .B2(new_n310), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n276), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT8), .ZN(new_n448));
  XNOR2_X1  g0248(.A(new_n388), .B(new_n448), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n253), .A2(new_n449), .ZN(new_n450));
  OAI21_X1  g0250(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n451));
  INV_X1    g0251(.A(G150), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n451), .B1(new_n452), .B2(new_n332), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n257), .B1(new_n450), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n337), .A2(G50), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n454), .B(new_n455), .C1(G50), .C2(new_n265), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n447), .A2(new_n456), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n445), .A2(new_n446), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n457), .B1(new_n320), .B2(new_n458), .ZN(new_n459));
  XNOR2_X1  g0259(.A(new_n456), .B(KEYINPUT9), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n458), .A2(G190), .ZN(new_n461));
  OAI21_X1  g0261(.A(G200), .B1(new_n445), .B2(new_n446), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(KEYINPUT10), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT10), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n460), .A2(new_n461), .A3(new_n465), .A4(new_n462), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n459), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n370), .A2(new_n437), .A3(new_n438), .A4(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n437), .ZN(new_n469));
  OAI21_X1  g0269(.A(KEYINPUT79), .B1(new_n469), .B2(new_n369), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n414), .A2(G264), .A3(G1698), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n353), .A2(G303), .ZN(new_n473));
  INV_X1    g0273(.A(G257), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n472), .B(new_n473), .C1(new_n474), .C2(new_n283), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(new_n291), .ZN(new_n476));
  OR2_X1    g0276(.A1(KEYINPUT5), .A2(G41), .ZN(new_n477));
  NAND2_X1  g0277(.A1(KEYINPUT5), .A2(G41), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n208), .A2(G45), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n482), .A2(G270), .A3(new_n308), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n291), .A2(new_n300), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n480), .B1(new_n477), .B2(new_n478), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AND2_X1   g0286(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n476), .A2(new_n487), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n265), .A2(G116), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n208), .A2(G33), .ZN(new_n490));
  AND3_X1   g0290(.A1(new_n270), .A2(new_n265), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n489), .B1(new_n491), .B2(G116), .ZN(new_n492));
  NAND2_X1  g0292(.A1(G33), .A2(G283), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n307), .A2(G97), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n217), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(G116), .ZN(new_n496));
  AOI22_X1  g0296(.A1(new_n256), .A2(new_n218), .B1(G20), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT20), .ZN(new_n499));
  OR2_X1    g0299(.A1(new_n499), .A2(KEYINPUT85), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(KEYINPUT85), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n498), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n495), .A2(KEYINPUT85), .A3(new_n499), .A4(new_n497), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n492), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n488), .A2(new_n504), .A3(G169), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT21), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AND3_X1   g0307(.A1(new_n492), .A2(new_n502), .A3(new_n503), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n476), .A2(new_n487), .A3(G190), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n483), .A2(new_n486), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n510), .B1(new_n291), .B2(new_n475), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n508), .B(new_n509), .C1(new_n429), .C2(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n276), .B1(new_n476), .B2(new_n487), .ZN(new_n513));
  AOI22_X1  g0313(.A1(new_n513), .A2(KEYINPUT21), .B1(new_n511), .B2(G179), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n507), .B(new_n512), .C1(new_n514), .C2(new_n508), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT86), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n488), .A2(KEYINPUT21), .A3(G169), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n511), .A2(G179), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n504), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n521), .A2(KEYINPUT86), .A3(new_n507), .A4(new_n512), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n517), .A2(new_n522), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n288), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT4), .ZN(new_n525));
  OAI21_X1  g0325(.A(G244), .B1(new_n281), .B2(new_n282), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n279), .A2(new_n280), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  AND2_X1   g0328(.A1(new_n279), .A2(new_n280), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n529), .A2(KEYINPUT4), .A3(G244), .A4(new_n414), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n524), .B(new_n528), .C1(new_n530), .C2(KEYINPUT80), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT80), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n526), .A2(new_n527), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n532), .B1(new_n533), .B2(KEYINPUT4), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n291), .B1(new_n531), .B2(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n291), .B1(new_n481), .B2(new_n479), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(G257), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n486), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n535), .A2(new_n320), .A3(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT82), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n535), .A2(new_n539), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n276), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n530), .A2(KEYINPUT80), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n533), .A2(new_n532), .A3(KEYINPUT4), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n545), .A2(new_n546), .A3(new_n528), .A4(new_n524), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n538), .B1(new_n547), .B2(new_n291), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n548), .A2(KEYINPUT82), .A3(new_n320), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n417), .A2(new_n205), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT6), .ZN(new_n551));
  NOR3_X1   g0351(.A1(new_n551), .A2(new_n204), .A3(G107), .ZN(new_n552));
  XNOR2_X1  g0352(.A(G97), .B(G107), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n552), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  OAI22_X1  g0354(.A1(new_n554), .A2(new_n217), .B1(new_n254), .B2(new_n332), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n257), .B1(new_n550), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n265), .A2(G97), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n557), .B1(new_n491), .B2(G97), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n542), .A2(new_n544), .A3(new_n549), .A4(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n535), .A2(G190), .A3(new_n539), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(KEYINPUT81), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n543), .A2(G200), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT81), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n548), .A2(new_n564), .A3(G190), .ZN(new_n565));
  INV_X1    g0365(.A(new_n559), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n562), .A2(new_n563), .A3(new_n565), .A4(new_n566), .ZN(new_n567));
  AND2_X1   g0367(.A1(new_n560), .A2(new_n567), .ZN(new_n568));
  OAI211_X1 g0368(.A(G257), .B(G1698), .C1(new_n281), .C2(new_n282), .ZN(new_n569));
  NAND2_X1  g0369(.A1(G33), .A2(G294), .ZN(new_n570));
  INV_X1    g0370(.A(G250), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n569), .B(new_n570), .C1(new_n283), .C2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n291), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n536), .A2(G264), .B1(new_n484), .B2(new_n485), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(G169), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT89), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n482), .A2(G264), .A3(new_n308), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(KEYINPUT90), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT90), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n536), .A2(new_n581), .A3(G264), .ZN(new_n582));
  AOI22_X1  g0382(.A1(new_n580), .A2(new_n582), .B1(new_n291), .B2(new_n572), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n583), .A2(G179), .A3(new_n486), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n575), .A2(KEYINPUT89), .A3(G169), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n578), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n374), .A2(KEYINPUT87), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n414), .A2(new_n217), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(KEYINPUT22), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT22), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n414), .A2(new_n217), .A3(new_n590), .A4(new_n587), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  AND2_X1   g0392(.A1(KEYINPUT88), .A2(KEYINPUT23), .ZN(new_n593));
  NOR2_X1   g0393(.A1(KEYINPUT88), .A2(KEYINPUT23), .ZN(new_n594));
  OAI22_X1  g0394(.A1(new_n593), .A2(new_n594), .B1(new_n209), .B2(G107), .ZN(new_n595));
  NAND2_X1  g0395(.A1(G33), .A2(G116), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n595), .B1(G20), .B2(new_n596), .ZN(new_n597));
  NOR3_X1   g0397(.A1(new_n217), .A2(KEYINPUT23), .A3(G107), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT24), .ZN(new_n600));
  AND3_X1   g0400(.A1(new_n592), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n600), .B1(new_n592), .B2(new_n599), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n257), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(KEYINPUT25), .B1(new_n268), .B2(new_n205), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n268), .A2(KEYINPUT25), .A3(new_n205), .ZN(new_n606));
  AOI22_X1  g0406(.A1(G107), .A2(new_n491), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n586), .A2(new_n608), .ZN(new_n609));
  AOI21_X1  g0409(.A(G200), .B1(new_n583), .B2(new_n486), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n575), .A2(G190), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n603), .B(new_n607), .C1(new_n610), .C2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT19), .ZN(new_n614));
  NOR3_X1   g0414(.A1(new_n614), .A2(new_n307), .A3(new_n204), .ZN(new_n615));
  OAI22_X1  g0415(.A1(new_n615), .A2(new_n330), .B1(G87), .B2(new_n206), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n327), .A2(new_n329), .A3(G33), .A4(G97), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n614), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n414), .A2(new_n217), .A3(G68), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n616), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n620), .A2(new_n257), .B1(new_n268), .B2(new_n334), .ZN(new_n621));
  INV_X1    g0421(.A(new_n334), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n491), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(KEYINPUT83), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n481), .A2(G274), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n480), .A2(G250), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n626), .B1(new_n291), .B2(new_n627), .ZN(new_n628));
  OAI211_X1 g0428(.A(G244), .B(G1698), .C1(new_n281), .C2(new_n282), .ZN(new_n629));
  INV_X1    g0429(.A(G238), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n596), .B(new_n629), .C1(new_n283), .C2(new_n630), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n628), .B1(new_n631), .B2(new_n291), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(G179), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n633), .B1(new_n276), .B2(new_n632), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT83), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n621), .A2(new_n635), .A3(new_n623), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n625), .A2(new_n634), .A3(new_n636), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n632), .A2(new_n429), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n632), .A2(G190), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n391), .A2(new_n490), .ZN(new_n641));
  OAI21_X1  g0441(.A(KEYINPUT84), .B1(new_n641), .B2(new_n374), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT84), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n491), .A2(new_n643), .A3(G87), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n639), .A2(new_n640), .A3(new_n621), .A4(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n637), .A2(new_n646), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n613), .A2(new_n647), .ZN(new_n648));
  AND4_X1   g0448(.A1(new_n471), .A2(new_n523), .A3(new_n568), .A4(new_n648), .ZN(G372));
  AND2_X1   g0449(.A1(new_n422), .A2(new_n427), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n323), .A2(new_n368), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n326), .A2(new_n434), .A3(new_n435), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n650), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n464), .A2(new_n466), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n459), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n471), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n507), .B1(new_n514), .B2(new_n508), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(new_n609), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n634), .A2(new_n624), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n646), .A2(new_n660), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n568), .A2(new_n612), .A3(new_n659), .A4(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n559), .B1(new_n548), .B2(G169), .ZN(new_n663));
  AOI21_X1  g0463(.A(KEYINPUT82), .B1(new_n548), .B2(new_n320), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT26), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n665), .A2(new_n661), .A3(new_n666), .A4(new_n549), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n665), .A2(new_n549), .A3(new_n646), .A4(new_n637), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(KEYINPUT26), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n662), .A2(new_n660), .A3(new_n667), .A4(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n655), .B1(new_n656), .B2(new_n671), .ZN(G369));
  NAND2_X1  g0472(.A1(new_n217), .A2(new_n264), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(G213), .A3(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(G343), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n657), .A2(new_n679), .ZN(new_n680));
  OAI22_X1  g0480(.A1(new_n613), .A2(new_n680), .B1(new_n609), .B2(new_n678), .ZN(new_n681));
  XOR2_X1   g0481(.A(new_n681), .B(KEYINPUT92), .Z(new_n682));
  NAND2_X1  g0482(.A1(new_n678), .A2(new_n504), .ZN(new_n683));
  XOR2_X1   g0483(.A(new_n683), .B(KEYINPUT91), .Z(new_n684));
  NAND2_X1  g0484(.A1(new_n523), .A2(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n685), .B1(new_n658), .B2(new_n684), .ZN(new_n686));
  INV_X1    g0486(.A(new_n613), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n608), .A2(new_n678), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g0489(.A(KEYINPUT89), .B1(new_n575), .B2(G169), .ZN(new_n690));
  AOI211_X1 g0490(.A(new_n577), .B(new_n276), .C1(new_n573), .C2(new_n574), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AOI22_X1  g0492(.A1(new_n692), .A2(new_n584), .B1(new_n603), .B2(new_n607), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(new_n678), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n689), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n686), .A2(G330), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n682), .A2(new_n696), .ZN(G399));
  INV_X1    g0497(.A(new_n212), .ZN(new_n698));
  OR3_X1    g0498(.A1(new_n698), .A2(KEYINPUT93), .A3(G41), .ZN(new_n699));
  OAI21_X1  g0499(.A(KEYINPUT93), .B1(new_n698), .B2(G41), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NOR3_X1   g0501(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n702));
  AND3_X1   g0502(.A1(new_n701), .A2(G1), .A3(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n216), .ZN(new_n704));
  INV_X1    g0504(.A(new_n701), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n703), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  XOR2_X1   g0506(.A(new_n706), .B(KEYINPUT28), .Z(new_n707));
  NAND2_X1  g0507(.A1(new_n670), .A2(new_n679), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT29), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(KEYINPUT94), .B1(new_n668), .B2(new_n666), .ZN(new_n711));
  OAI211_X1 g0511(.A(KEYINPUT94), .B(new_n666), .C1(new_n560), .C2(new_n647), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n665), .A2(new_n661), .A3(KEYINPUT26), .A4(new_n549), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  OAI211_X1 g0515(.A(new_n612), .B(new_n661), .C1(new_n693), .C2(new_n657), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n560), .A2(new_n567), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n660), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  OAI211_X1 g0518(.A(KEYINPUT29), .B(new_n679), .C1(new_n715), .C2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n710), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(G330), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n648), .A2(new_n523), .A3(new_n568), .A4(new_n679), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT30), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n511), .A2(new_n583), .A3(G179), .A4(new_n632), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n723), .B1(new_n724), .B2(new_n543), .ZN(new_n725));
  NOR3_X1   g0525(.A1(new_n511), .A2(G179), .A3(new_n632), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n583), .A2(new_n486), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n726), .A2(new_n543), .A3(new_n727), .ZN(new_n728));
  AND2_X1   g0528(.A1(new_n583), .A2(new_n632), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n488), .A2(new_n320), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n729), .A2(new_n730), .A3(new_n548), .A4(KEYINPUT30), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n725), .A2(new_n728), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(new_n678), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(KEYINPUT31), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT31), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n732), .A2(new_n735), .A3(new_n678), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n721), .B1(new_n722), .B2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n720), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n707), .B1(new_n741), .B2(G1), .ZN(G364));
  NOR2_X1   g0542(.A1(new_n330), .A2(new_n263), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G45), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(G1), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n705), .A2(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n746), .B1(new_n686), .B2(G330), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n747), .B1(G330), .B2(new_n686), .ZN(new_n748));
  NOR2_X1   g0548(.A1(G13), .A2(G33), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(G20), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n218), .B1(G20), .B2(new_n276), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n212), .A2(new_n414), .ZN(new_n754));
  INV_X1    g0554(.A(G355), .ZN(new_n755));
  OAI22_X1  g0555(.A1(new_n754), .A2(new_n755), .B1(G116), .B2(new_n212), .ZN(new_n756));
  XOR2_X1   g0556(.A(new_n756), .B(KEYINPUT95), .Z(new_n757));
  AND2_X1   g0557(.A1(new_n295), .A2(new_n297), .ZN(new_n758));
  AND2_X1   g0558(.A1(new_n704), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n698), .A2(new_n414), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AOI211_X1 g0561(.A(new_n759), .B(new_n761), .C1(G45), .C2(new_n248), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n753), .B1(new_n757), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(new_n746), .ZN(new_n764));
  NOR2_X1   g0564(.A1(G179), .A2(G200), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(G190), .ZN(new_n766));
  AND2_X1   g0566(.A1(new_n330), .A2(new_n766), .ZN(new_n767));
  XOR2_X1   g0567(.A(new_n767), .B(KEYINPUT97), .Z(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(new_n204), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n217), .A2(new_n320), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n771), .A2(new_n325), .A3(new_n429), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n770), .B1(G77), .B2(new_n773), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n771), .A2(G190), .A3(G200), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n771), .A2(new_n325), .A3(G200), .ZN(new_n776));
  OAI221_X1 g0576(.A(new_n774), .B1(new_n221), .B2(new_n775), .C1(new_n251), .C2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n429), .A2(G179), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n217), .A2(new_n779), .A3(G190), .ZN(new_n780));
  OR2_X1    g0580(.A1(new_n780), .A2(KEYINPUT96), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(KEYINPUT96), .ZN(new_n782));
  AND2_X1   g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(G107), .ZN(new_n784));
  NOR3_X1   g0584(.A1(new_n779), .A2(new_n209), .A3(new_n325), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n414), .B1(new_n786), .B2(new_n374), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n771), .A2(G190), .A3(new_n429), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n787), .B1(G58), .B2(new_n789), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n330), .A2(new_n325), .A3(new_n765), .ZN(new_n791));
  OAI21_X1  g0591(.A(KEYINPUT32), .B1(new_n791), .B2(new_n405), .ZN(new_n792));
  OR3_X1    g0592(.A1(new_n791), .A2(KEYINPUT32), .A3(new_n405), .ZN(new_n793));
  NAND4_X1  g0593(.A1(new_n784), .A2(new_n790), .A3(new_n792), .A4(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n776), .ZN(new_n795));
  XNOR2_X1  g0595(.A(KEYINPUT33), .B(G317), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(G311), .ZN(new_n798));
  XNOR2_X1  g0598(.A(KEYINPUT98), .B(G326), .ZN(new_n799));
  OAI221_X1 g0599(.A(new_n797), .B1(new_n798), .B2(new_n772), .C1(new_n775), .C2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(G294), .ZN(new_n801));
  INV_X1    g0601(.A(G303), .ZN(new_n802));
  OAI221_X1 g0602(.A(new_n353), .B1(new_n767), .B2(new_n801), .C1(new_n786), .C2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n791), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n803), .B1(G329), .B2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(G322), .ZN(new_n806));
  INV_X1    g0606(.A(G283), .ZN(new_n807));
  INV_X1    g0607(.A(new_n783), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n805), .B1(new_n806), .B2(new_n788), .C1(new_n807), .C2(new_n808), .ZN(new_n809));
  OAI22_X1  g0609(.A1(new_n777), .A2(new_n794), .B1(new_n800), .B2(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n764), .B1(new_n810), .B2(new_n752), .ZN(new_n811));
  INV_X1    g0611(.A(new_n751), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n811), .B1(new_n686), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n748), .A2(new_n813), .ZN(G396));
  NAND3_X1  g0614(.A1(new_n364), .A2(new_n367), .A3(new_n679), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n276), .B1(new_n359), .B2(new_n342), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n366), .B1(KEYINPUT75), .B2(new_n816), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n356), .A2(KEYINPUT75), .A3(new_n320), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n818), .A2(new_n340), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n365), .A2(new_n679), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n821), .B1(new_n357), .B2(new_n360), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n815), .B1(new_n820), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n708), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n821), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n361), .A2(new_n825), .B1(new_n364), .B2(new_n367), .ZN(new_n826));
  INV_X1    g0626(.A(new_n815), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n560), .A2(new_n647), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n667), .B1(new_n829), .B2(new_n666), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n828), .B(new_n679), .C1(new_n718), .C2(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n824), .A2(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n746), .B1(new_n832), .B2(new_n739), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n833), .B1(new_n739), .B2(new_n832), .ZN(new_n834));
  INV_X1    g0634(.A(new_n746), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n752), .A2(new_n749), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n835), .B1(new_n254), .B2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n775), .ZN(new_n838));
  AOI22_X1  g0638(.A1(G294), .A2(new_n789), .B1(new_n838), .B2(G303), .ZN(new_n839));
  XOR2_X1   g0639(.A(KEYINPUT99), .B(G283), .Z(new_n840));
  OAI221_X1 g0640(.A(new_n839), .B1(new_n496), .B2(new_n772), .C1(new_n776), .C2(new_n840), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n808), .A2(new_n374), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n353), .B1(new_n798), .B2(new_n791), .C1(new_n786), .C2(new_n205), .ZN(new_n843));
  NOR4_X1   g0643(.A1(new_n841), .A2(new_n842), .A3(new_n770), .A4(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(G137), .ZN(new_n845));
  OAI22_X1  g0645(.A1(new_n845), .A2(new_n775), .B1(new_n776), .B2(new_n452), .ZN(new_n846));
  XNOR2_X1  g0646(.A(new_n846), .B(KEYINPUT100), .ZN(new_n847));
  INV_X1    g0647(.A(G143), .ZN(new_n848));
  OAI221_X1 g0648(.A(new_n847), .B1(new_n848), .B2(new_n788), .C1(new_n405), .C2(new_n772), .ZN(new_n849));
  XNOR2_X1  g0649(.A(new_n849), .B(KEYINPUT34), .ZN(new_n850));
  INV_X1    g0650(.A(new_n767), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(G58), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n353), .B1(new_n785), .B2(G50), .ZN(new_n853));
  INV_X1    g0653(.A(G132), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n852), .B(new_n853), .C1(new_n854), .C2(new_n791), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n855), .B1(new_n783), .B2(G68), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n844), .B1(new_n850), .B2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n752), .ZN(new_n858));
  OAI221_X1 g0658(.A(new_n837), .B1(new_n750), .B2(new_n828), .C1(new_n857), .C2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n834), .A2(new_n859), .ZN(G384));
  NOR3_X1   g0660(.A1(new_n217), .A2(new_n496), .A3(new_n218), .ZN(new_n861));
  XOR2_X1   g0661(.A(new_n554), .B(KEYINPUT101), .Z(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT35), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n861), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n865), .B1(new_n864), .B2(new_n863), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n866), .B(KEYINPUT102), .ZN(new_n867));
  XNOR2_X1  g0667(.A(new_n867), .B(KEYINPUT36), .ZN(new_n868));
  OR3_X1    g0668(.A1(new_n216), .A2(new_n254), .A3(new_n395), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n221), .A2(G68), .ZN(new_n870));
  AOI211_X1 g0670(.A(new_n208), .B(G13), .C1(new_n869), .C2(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n722), .A2(new_n737), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT107), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n722), .A2(new_n737), .A3(KEYINPUT107), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT106), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n421), .A2(new_n676), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n425), .A2(new_n382), .A3(new_n386), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT37), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n881), .A2(new_n882), .A3(new_n883), .A4(new_n432), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n432), .B1(new_n387), .B2(new_n421), .ZN(new_n885));
  OAI21_X1  g0685(.A(KEYINPUT37), .B1(new_n885), .B2(new_n880), .ZN(new_n886));
  AOI22_X1  g0686(.A1(new_n884), .A2(new_n886), .B1(new_n436), .B2(new_n880), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n879), .B1(new_n887), .B2(KEYINPUT38), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n886), .A2(new_n884), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n436), .A2(new_n880), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT38), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n891), .A2(KEYINPUT106), .A3(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT104), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n397), .B1(new_n400), .B2(new_n401), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n270), .B1(new_n895), .B2(new_n419), .ZN(new_n896));
  AOI22_X1  g0696(.A1(new_n894), .A2(new_n896), .B1(new_n403), .B2(new_n412), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n257), .B1(new_n410), .B2(KEYINPUT16), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(KEYINPUT104), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n394), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n432), .B1(new_n900), .B2(new_n676), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n900), .A2(new_n387), .ZN(new_n902));
  OAI21_X1  g0702(.A(KEYINPUT37), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n900), .A2(new_n676), .ZN(new_n904));
  AOI22_X1  g0704(.A1(new_n903), .A2(new_n884), .B1(new_n436), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(KEYINPUT38), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n888), .A2(new_n893), .A3(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n274), .A2(new_n679), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n323), .A2(new_n326), .A3(new_n909), .ZN(new_n910));
  OR2_X1    g0710(.A1(new_n321), .A2(new_n322), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n908), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n823), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n878), .A2(new_n907), .A3(new_n913), .ZN(new_n914));
  AND2_X1   g0714(.A1(new_n914), .A2(KEYINPUT40), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n903), .A2(new_n884), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n436), .A2(new_n904), .ZN(new_n917));
  AOI21_X1  g0717(.A(KEYINPUT38), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n906), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT40), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n878), .A2(new_n920), .A3(new_n921), .A4(new_n913), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n471), .B(new_n878), .C1(new_n915), .C2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n914), .A2(KEYINPUT40), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n925), .B(new_n922), .C1(new_n656), .C2(new_n877), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n924), .A2(G330), .A3(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT39), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n907), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n911), .A2(new_n275), .A3(new_n679), .ZN(new_n930));
  XOR2_X1   g0730(.A(new_n930), .B(KEYINPUT105), .Z(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n919), .A2(KEYINPUT39), .A3(new_n906), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n929), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n910), .A2(new_n912), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n831), .A2(KEYINPUT103), .A3(new_n815), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(KEYINPUT103), .B1(new_n831), .B2(new_n815), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n920), .B(new_n935), .C1(new_n937), .C2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(new_n676), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n650), .A2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n934), .A2(new_n939), .A3(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n710), .A2(new_n471), .A3(new_n719), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(new_n655), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n943), .B(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n927), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n208), .B2(new_n743), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n927), .A2(new_n946), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n872), .B1(new_n948), .B2(new_n949), .ZN(G367));
  OAI221_X1 g0750(.A(new_n753), .B1(new_n212), .B2(new_n334), .C1(new_n761), .C2(new_n241), .ZN(new_n951));
  AND2_X1   g0751(.A1(new_n746), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n621), .A2(new_n645), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(new_n678), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n661), .A2(new_n954), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n660), .A2(new_n954), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n785), .A2(G116), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT46), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n958), .A2(new_n959), .B1(new_n205), .B2(new_n767), .ZN(new_n960));
  AOI211_X1 g0760(.A(new_n414), .B(new_n960), .C1(new_n959), .C2(new_n958), .ZN(new_n961));
  INV_X1    g0761(.A(new_n780), .ZN(new_n962));
  INV_X1    g0762(.A(G317), .ZN(new_n963));
  OAI221_X1 g0763(.A(new_n961), .B1(new_n204), .B2(new_n962), .C1(new_n963), .C2(new_n791), .ZN(new_n964));
  INV_X1    g0764(.A(new_n840), .ZN(new_n965));
  AOI22_X1  g0765(.A1(G311), .A2(new_n838), .B1(new_n773), .B2(new_n965), .ZN(new_n966));
  OAI221_X1 g0766(.A(new_n966), .B1(new_n801), .B2(new_n776), .C1(new_n802), .C2(new_n788), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n768), .A2(G68), .ZN(new_n968));
  OAI221_X1 g0768(.A(new_n968), .B1(new_n221), .B2(new_n772), .C1(new_n405), .C2(new_n776), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n353), .B1(new_n785), .B2(G58), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n970), .B1(new_n845), .B2(new_n791), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n971), .B1(G77), .B2(new_n780), .ZN(new_n972));
  OAI221_X1 g0772(.A(new_n972), .B1(new_n848), .B2(new_n775), .C1(new_n452), .C2(new_n788), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n964), .A2(new_n967), .B1(new_n969), .B2(new_n973), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n974), .B(KEYINPUT47), .Z(new_n975));
  OAI221_X1 g0775(.A(new_n952), .B1(new_n812), .B2(new_n957), .C1(new_n975), .C2(new_n858), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n701), .B(KEYINPUT41), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n686), .A2(G330), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n613), .A2(new_n680), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(new_n680), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n982), .B1(new_n695), .B2(new_n983), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n980), .B(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n986), .A2(new_n739), .A3(new_n720), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT44), .ZN(new_n988));
  OAI211_X1 g0788(.A(new_n560), .B(new_n567), .C1(new_n566), .C2(new_n679), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n665), .A2(new_n549), .A3(new_n678), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n988), .B1(new_n682), .B2(new_n991), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n681), .B(KEYINPUT92), .ZN(new_n993));
  AND2_X1   g0793(.A1(new_n989), .A2(new_n990), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n993), .A2(KEYINPUT44), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n992), .A2(new_n995), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n682), .A2(KEYINPUT45), .A3(new_n991), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT45), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(new_n993), .B2(new_n994), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n996), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT110), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n1001), .A2(new_n1002), .A3(new_n696), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n696), .A2(new_n1002), .ZN(new_n1004));
  OR2_X1    g0804(.A1(new_n696), .A2(new_n1002), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n996), .A2(new_n1000), .A3(new_n1004), .A4(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n987), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n979), .B1(new_n1007), .B2(new_n740), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n745), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n696), .A2(new_n994), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n991), .A2(new_n981), .ZN(new_n1013));
  AND2_X1   g0813(.A1(new_n1013), .A2(KEYINPUT42), .ZN(new_n1014));
  OR2_X1    g0814(.A1(new_n989), .A2(new_n609), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n678), .B1(new_n1015), .B2(new_n560), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n1013), .A2(KEYINPUT42), .ZN(new_n1017));
  NOR3_X1   g0817(.A1(new_n1014), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n957), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(KEYINPUT108), .B(KEYINPUT43), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1018), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n957), .A2(KEYINPUT43), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1021), .B1(new_n1018), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT109), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1023), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1027), .B1(new_n1023), .B2(new_n1026), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1012), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1030), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1032), .A2(new_n1011), .A3(new_n1028), .ZN(new_n1033));
  AND2_X1   g0833(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n977), .B1(new_n1010), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n1035), .ZN(G387));
  NAND2_X1  g0836(.A1(new_n740), .A2(new_n985), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n987), .A2(new_n705), .A3(new_n1037), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n689), .A2(new_n694), .A3(new_n751), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n760), .B1(new_n238), .B2(new_n758), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1040), .B1(new_n702), .B2(new_n754), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n333), .A2(G50), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT50), .ZN(new_n1043));
  AOI21_X1  g0843(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1043), .A2(new_n702), .A3(new_n1044), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n1041), .A2(new_n1045), .B1(new_n205), .B2(new_n698), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n753), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n746), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(G50), .A2(new_n789), .B1(new_n795), .B2(new_n389), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(new_n251), .B2(new_n772), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n804), .A2(G150), .B1(new_n785), .B2(G77), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT111), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n783), .A2(G97), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n768), .A2(new_n622), .ZN(new_n1054));
  NAND4_X1  g0854(.A1(new_n1052), .A2(new_n1053), .A3(new_n414), .A4(new_n1054), .ZN(new_n1055));
  OAI21_X1  g0855(.A(KEYINPUT112), .B1(new_n775), .B2(new_n405), .ZN(new_n1056));
  OR3_X1    g0856(.A1(new_n775), .A2(KEYINPUT112), .A3(new_n405), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n1050), .B(new_n1055), .C1(new_n1056), .C2(new_n1057), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT113), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n414), .B1(new_n780), .B2(G116), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(G303), .A2(new_n773), .B1(new_n789), .B2(G317), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n1061), .B1(new_n798), .B2(new_n776), .C1(new_n806), .C2(new_n775), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT48), .ZN(new_n1063));
  OR2_X1    g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n851), .A2(new_n965), .B1(new_n785), .B2(G294), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1064), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT49), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n1060), .B1(new_n791), .B2(new_n799), .C1(new_n1067), .C2(new_n1068), .ZN(new_n1069));
  AND2_X1   g0869(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1059), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1048), .B1(new_n1071), .B2(new_n752), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n986), .A2(new_n745), .B1(new_n1039), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1038), .A2(new_n1073), .ZN(G393));
  NOR2_X1   g0874(.A1(new_n1007), .A2(new_n701), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1003), .A2(new_n987), .A3(new_n1006), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1009), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n994), .A2(new_n751), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n753), .B1(new_n204), .B2(new_n212), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(new_n760), .B2(new_n245), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n452), .A2(new_n775), .B1(new_n788), .B2(new_n405), .ZN(new_n1082));
  XOR2_X1   g0882(.A(new_n1082), .B(KEYINPUT51), .Z(new_n1083));
  NAND2_X1  g0883(.A1(new_n768), .A2(G77), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n353), .B1(new_n785), .B2(G68), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1084), .B(new_n1085), .C1(new_n848), .C2(new_n791), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n221), .A2(new_n776), .B1(new_n772), .B2(new_n333), .ZN(new_n1087));
  OR4_X1    g0887(.A1(new_n842), .A2(new_n1083), .A3(new_n1086), .A4(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n414), .B1(new_n785), .B2(new_n965), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n784), .B(new_n1089), .C1(new_n806), .C2(new_n791), .ZN(new_n1090));
  XOR2_X1   g0890(.A(new_n1090), .B(KEYINPUT115), .Z(new_n1091));
  OAI22_X1  g0891(.A1(new_n798), .A2(new_n788), .B1(new_n775), .B2(new_n963), .ZN(new_n1092));
  XOR2_X1   g0892(.A(KEYINPUT114), .B(KEYINPUT52), .Z(new_n1093));
  XNOR2_X1  g0893(.A(new_n1092), .B(new_n1093), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n776), .A2(new_n802), .B1(new_n496), .B2(new_n767), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n1095), .A2(KEYINPUT116), .B1(G294), .B2(new_n773), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1094), .B(new_n1096), .C1(KEYINPUT116), .C2(new_n1095), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1088), .B1(new_n1091), .B2(new_n1097), .ZN(new_n1098));
  AOI211_X1 g0898(.A(new_n835), .B(new_n1081), .C1(new_n1098), .C2(new_n752), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1078), .B1(new_n1079), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1077), .A2(new_n1100), .ZN(G390));
  NAND2_X1  g0901(.A1(new_n831), .A2(new_n815), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT103), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n936), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n738), .A2(new_n828), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n935), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n875), .A2(G330), .A3(new_n876), .A4(new_n913), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n875), .A2(G330), .A3(new_n828), .A4(new_n876), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(new_n1107), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n826), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n679), .B(new_n1113), .C1(new_n715), .C2(new_n718), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n873), .A2(new_n913), .A3(G330), .ZN(new_n1115));
  AND3_X1   g0915(.A1(new_n1114), .A2(new_n1115), .A3(new_n815), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n1105), .A2(new_n1110), .B1(new_n1112), .B2(new_n1116), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n471), .A2(G330), .A3(new_n875), .A4(new_n876), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1118), .A2(new_n944), .A3(new_n655), .ZN(new_n1119));
  OAI21_X1  g0919(.A(KEYINPUT117), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1110), .A2(new_n1105), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1112), .A2(new_n1116), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(KEYINPUT117), .ZN(new_n1124));
  AND3_X1   g0924(.A1(new_n1118), .A2(new_n944), .A3(new_n655), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1123), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1120), .A2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1107), .B1(new_n1104), .B2(new_n936), .ZN(new_n1128));
  AOI21_X1  g0928(.A(KEYINPUT38), .B1(new_n889), .B2(new_n890), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n1129), .A2(KEYINPUT106), .B1(KEYINPUT38), .B2(new_n905), .ZN(new_n1130));
  AOI21_X1  g0930(.A(KEYINPUT39), .B1(new_n1130), .B2(new_n888), .ZN(new_n1131));
  AND3_X1   g0931(.A1(new_n916), .A2(KEYINPUT38), .A3(new_n917), .ZN(new_n1132));
  NOR3_X1   g0932(.A1(new_n1132), .A2(new_n918), .A3(new_n928), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n1128), .A2(new_n932), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n907), .A2(new_n931), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1107), .B1(new_n1114), .B2(new_n815), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1134), .A2(new_n1138), .A3(new_n1115), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n877), .A2(new_n721), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n935), .B1(new_n937), .B2(new_n938), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n1141), .A2(new_n931), .B1(new_n929), .B2(new_n933), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n913), .B(new_n1140), .C1(new_n1142), .C2(new_n1137), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1127), .A2(new_n1139), .A3(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1115), .ZN(new_n1145));
  NOR3_X1   g0945(.A1(new_n1142), .A2(new_n1137), .A3(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1109), .B1(new_n1134), .B2(new_n1138), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1126), .B(new_n1120), .C1(new_n1146), .C2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1144), .A2(new_n1148), .A3(new_n705), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n749), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n785), .A2(G150), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n1152), .B(KEYINPUT53), .ZN(new_n1153));
  AND2_X1   g0953(.A1(new_n804), .A2(G125), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n962), .A2(new_n221), .ZN(new_n1155));
  NOR4_X1   g0955(.A1(new_n1153), .A2(new_n353), .A3(new_n1154), .A4(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n838), .A2(G128), .ZN(new_n1157));
  XOR2_X1   g0957(.A(KEYINPUT54), .B(G143), .Z(new_n1158));
  XNOR2_X1  g0958(.A(new_n1158), .B(KEYINPUT118), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n773), .A2(new_n1159), .B1(new_n795), .B2(G137), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n768), .A2(G159), .B1(G132), .B2(new_n789), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n1156), .A2(new_n1157), .A3(new_n1160), .A4(new_n1161), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(G107), .A2(new_n795), .B1(new_n838), .B2(G283), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1163), .B1(new_n204), .B2(new_n772), .ZN(new_n1164));
  XOR2_X1   g0964(.A(new_n1164), .B(KEYINPUT119), .Z(new_n1165));
  AOI21_X1  g0965(.A(new_n414), .B1(new_n785), .B2(G87), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n1166), .B(KEYINPUT120), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(G294), .B2(new_n804), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n783), .A2(G68), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n789), .A2(G116), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1168), .A2(new_n1169), .A3(new_n1084), .A4(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1162), .B1(new_n1165), .B2(new_n1171), .ZN(new_n1172));
  AND2_X1   g0972(.A1(new_n1172), .A2(new_n752), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n835), .B(new_n1173), .C1(new_n449), .C2(new_n836), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n1150), .A2(new_n745), .B1(new_n1151), .B2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1149), .A2(new_n1175), .ZN(G378));
  INV_X1    g0976(.A(KEYINPUT123), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n456), .A2(new_n940), .ZN(new_n1178));
  OR2_X1    g0978(.A1(new_n467), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n467), .A2(new_n1178), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1179), .A2(new_n1180), .A3(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1181), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n943), .A2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n721), .B1(new_n925), .B2(new_n922), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1185), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n934), .A2(new_n939), .A3(new_n942), .A4(new_n1188), .ZN(new_n1189));
  AND3_X1   g0989(.A1(new_n1186), .A2(new_n1187), .A3(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1187), .B1(new_n1186), .B2(new_n1189), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1177), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g0992(.A(G330), .B1(new_n915), .B2(new_n923), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1133), .B1(new_n928), .B2(new_n907), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n941), .B1(new_n1194), .B2(new_n932), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1188), .B1(new_n1195), .B2(new_n939), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1189), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1193), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1186), .A2(new_n1187), .A3(new_n1189), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1198), .A2(KEYINPUT123), .A3(new_n1199), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1192), .A2(new_n745), .A3(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n836), .A2(new_n221), .ZN(new_n1202));
  AND2_X1   g1002(.A1(new_n746), .A2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n968), .B1(new_n334), .B2(new_n772), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(G97), .A2(new_n795), .B1(new_n838), .B2(G116), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1205), .B1(new_n205), .B2(new_n788), .ZN(new_n1206));
  AOI211_X1 g1006(.A(G41), .B(new_n414), .C1(new_n785), .C2(G77), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n780), .A2(G58), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1207), .B(new_n1208), .C1(new_n807), .C2(new_n791), .ZN(new_n1209));
  NOR3_X1   g1009(.A1(new_n1204), .A2(new_n1206), .A3(new_n1209), .ZN(new_n1210));
  XOR2_X1   g1010(.A(new_n1210), .B(KEYINPUT121), .Z(new_n1211));
  OR2_X1    g1011(.A1(new_n1211), .A2(KEYINPUT58), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1211), .A2(KEYINPUT58), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n221), .B1(new_n281), .B2(G41), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(G125), .A2(new_n838), .B1(new_n795), .B2(G132), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n789), .A2(G128), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n1215), .B(new_n1216), .C1(new_n769), .C2(new_n452), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1159), .A2(new_n785), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1218), .B1(new_n845), .B2(new_n772), .ZN(new_n1219));
  OR3_X1    g1019(.A1(new_n1217), .A2(KEYINPUT59), .A3(new_n1219), .ZN(new_n1220));
  OAI21_X1  g1020(.A(KEYINPUT59), .B1(new_n1217), .B2(new_n1219), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n780), .A2(G159), .ZN(new_n1222));
  AOI211_X1 g1022(.A(G33), .B(G41), .C1(new_n804), .C2(G124), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1220), .A2(new_n1221), .A3(new_n1222), .A4(new_n1223), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .A4(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(KEYINPUT122), .B1(new_n1225), .B2(new_n752), .ZN(new_n1226));
  AND3_X1   g1026(.A1(new_n1225), .A2(KEYINPUT122), .A3(new_n752), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n1203), .B1(new_n1188), .B2(new_n750), .C1(new_n1226), .C2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1201), .A2(new_n1228), .ZN(new_n1229));
  XNOR2_X1  g1029(.A(new_n1119), .B(KEYINPUT124), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  NOR3_X1   g1031(.A1(new_n1117), .A2(KEYINPUT117), .A3(new_n1119), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1124), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1143), .A2(new_n1139), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1231), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1236), .A2(new_n1192), .A3(new_n1200), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT57), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  OAI21_X1  g1039(.A(KEYINPUT57), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n701), .B1(new_n1241), .B2(new_n1236), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1229), .B1(new_n1239), .B2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(G375));
  NOR2_X1   g1044(.A1(new_n935), .A2(new_n750), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n353), .B1(new_n786), .B2(new_n204), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1246), .B1(new_n804), .B2(G303), .ZN(new_n1247));
  OAI211_X1 g1047(.A(new_n1054), .B(new_n1247), .C1(new_n808), .C2(new_n254), .ZN(new_n1248));
  OAI22_X1  g1048(.A1(new_n205), .A2(new_n772), .B1(new_n776), .B2(new_n496), .ZN(new_n1249));
  OAI22_X1  g1049(.A1(new_n807), .A2(new_n788), .B1(new_n775), .B2(new_n801), .ZN(new_n1250));
  NOR3_X1   g1050(.A1(new_n1248), .A2(new_n1249), .A3(new_n1250), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n769), .A2(new_n221), .B1(new_n845), .B2(new_n788), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n795), .A2(new_n1159), .ZN(new_n1253));
  OAI221_X1 g1053(.A(new_n1253), .B1(new_n854), .B2(new_n775), .C1(new_n452), .C2(new_n772), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n353), .B1(new_n785), .B2(G159), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n804), .A2(G128), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1255), .A2(new_n1256), .A3(new_n1208), .ZN(new_n1257));
  NOR3_X1   g1057(.A1(new_n1252), .A2(new_n1254), .A3(new_n1257), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n752), .B1(new_n1251), .B2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n836), .A2(new_n251), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1259), .A2(new_n746), .A3(new_n1260), .ZN(new_n1261));
  OAI22_X1  g1061(.A1(new_n1117), .A2(new_n1009), .B1(new_n1245), .B2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1120), .A2(new_n1126), .A3(new_n1264), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1263), .B1(new_n1265), .B2(new_n978), .ZN(G381));
  INV_X1    g1066(.A(G378), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1243), .A2(new_n1267), .ZN(new_n1268));
  AND2_X1   g1068(.A1(new_n1077), .A2(new_n1100), .ZN(new_n1269));
  INV_X1    g1069(.A(G384), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(G393), .A2(G396), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1269), .A2(new_n1270), .A3(new_n1271), .ZN(new_n1272));
  OR4_X1    g1072(.A1(G387), .A2(new_n1268), .A3(G381), .A4(new_n1272), .ZN(G407));
  INV_X1    g1073(.A(G213), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1274), .A2(G343), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1268), .A2(new_n1276), .ZN(new_n1277));
  XNOR2_X1  g1077(.A(new_n1277), .B(KEYINPUT125), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1278), .A2(G213), .A3(G407), .ZN(G409));
  OAI21_X1  g1079(.A(new_n745), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1280));
  AND4_X1   g1080(.A1(new_n1149), .A2(new_n1175), .A3(new_n1228), .A4(new_n1280), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1236), .A2(new_n1192), .A3(new_n979), .A4(new_n1200), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1275), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT60), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1264), .A2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(new_n705), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1286), .B1(KEYINPUT60), .B2(new_n1265), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1270), .B1(new_n1287), .B2(new_n1262), .ZN(new_n1288));
  AND2_X1   g1088(.A1(new_n1265), .A2(KEYINPUT60), .ZN(new_n1289));
  OAI211_X1 g1089(.A(G384), .B(new_n1263), .C1(new_n1289), .C2(new_n1286), .ZN(new_n1290));
  AND2_X1   g1090(.A1(new_n1288), .A2(new_n1290), .ZN(new_n1291));
  OAI211_X1 g1091(.A(new_n1283), .B(new_n1291), .C1(new_n1243), .C2(new_n1267), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(KEYINPUT62), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT61), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1275), .A2(G2897), .ZN(new_n1295));
  AND3_X1   g1095(.A1(new_n1288), .A2(new_n1290), .A3(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1295), .B1(new_n1288), .B2(new_n1290), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1239), .A2(new_n1242), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1229), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1267), .B1(new_n1299), .B2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(new_n1276), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1298), .B1(new_n1301), .B2(new_n1303), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1230), .B1(new_n1150), .B2(new_n1127), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n705), .B1(new_n1240), .B2(new_n1305), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1306), .B1(new_n1238), .B2(new_n1237), .ZN(new_n1307));
  OAI21_X1  g1107(.A(G378), .B1(new_n1307), .B2(new_n1229), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT62), .ZN(new_n1309));
  NAND4_X1  g1109(.A1(new_n1308), .A2(new_n1309), .A3(new_n1283), .A4(new_n1291), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1293), .A2(new_n1294), .A3(new_n1304), .A4(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1312), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1269), .B1(new_n1313), .B2(new_n977), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1035), .A2(G390), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT127), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1317), .B1(new_n1035), .B2(G390), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1271), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT126), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(G393), .A2(G396), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1319), .A2(new_n1320), .A3(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1322), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1320), .B1(new_n1319), .B2(new_n1321), .ZN(new_n1324));
  NOR2_X1   g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1316), .B1(new_n1318), .B2(new_n1325), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1324), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1327), .A2(new_n1322), .ZN(new_n1328));
  NAND4_X1  g1128(.A1(new_n1328), .A2(new_n1314), .A3(new_n1315), .A4(new_n1317), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1326), .A2(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1311), .A2(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1308), .A2(new_n1283), .ZN(new_n1333));
  AOI21_X1  g1133(.A(KEYINPUT61), .B1(new_n1333), .B2(new_n1298), .ZN(new_n1334));
  INV_X1    g1134(.A(KEYINPUT63), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1292), .A2(new_n1335), .ZN(new_n1336));
  NAND4_X1  g1136(.A1(new_n1308), .A2(KEYINPUT63), .A3(new_n1283), .A4(new_n1291), .ZN(new_n1337));
  NAND4_X1  g1137(.A1(new_n1334), .A2(new_n1330), .A3(new_n1336), .A4(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1332), .A2(new_n1338), .ZN(G405));
  INV_X1    g1139(.A(new_n1291), .ZN(new_n1340));
  AND3_X1   g1140(.A1(new_n1330), .A2(new_n1268), .A3(new_n1308), .ZN(new_n1341));
  AOI21_X1  g1141(.A(new_n1330), .B1(new_n1268), .B2(new_n1308), .ZN(new_n1342));
  OAI21_X1  g1142(.A(new_n1340), .B1(new_n1341), .B2(new_n1342), .ZN(new_n1343));
  INV_X1    g1143(.A(new_n1268), .ZN(new_n1344));
  OAI21_X1  g1144(.A(new_n1331), .B1(new_n1344), .B2(new_n1301), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1330), .A2(new_n1268), .A3(new_n1308), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1345), .A2(new_n1291), .A3(new_n1346), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1343), .A2(new_n1347), .ZN(G402));
endmodule


