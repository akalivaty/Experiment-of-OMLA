

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U557 ( .A1(G2104), .A2(G2105), .ZN(n906) );
  INV_X2 U558 ( .A(n766), .ZN(n739) );
  NOR2_X2 U559 ( .A1(G2105), .A2(n559), .ZN(n573) );
  BUF_X2 U560 ( .A(n611), .Z(n523) );
  XNOR2_X1 U561 ( .A(KEYINPUT67), .B(n547), .ZN(n611) );
  NAND2_X1 U562 ( .A1(n718), .A2(n717), .ZN(n722) );
  INV_X1 U563 ( .A(KEYINPUT100), .ZN(n745) );
  INV_X1 U564 ( .A(KEYINPUT29), .ZN(n735) );
  NOR2_X1 U565 ( .A1(n722), .A2(n537), .ZN(n536) );
  NOR2_X1 U566 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U567 ( .A1(n800), .A2(n801), .ZN(n766) );
  AND2_X1 U568 ( .A1(n583), .A2(n530), .ZN(n800) );
  NOR2_X1 U569 ( .A1(n532), .A2(n531), .ZN(n530) );
  INV_X1 U570 ( .A(G40), .ZN(n531) );
  INV_X1 U571 ( .A(n584), .ZN(n532) );
  NOR2_X1 U572 ( .A1(G164), .A2(G1384), .ZN(n801) );
  AND2_X1 U573 ( .A1(G2105), .A2(n559), .ZN(n560) );
  NAND2_X1 U574 ( .A1(G114), .A2(n906), .ZN(n555) );
  XNOR2_X2 U575 ( .A(n544), .B(n543), .ZN(n612) );
  XOR2_X1 U576 ( .A(KEYINPUT31), .B(n756), .Z(n524) );
  XOR2_X1 U577 ( .A(n536), .B(KEYINPUT98), .Z(n525) );
  OR2_X1 U578 ( .A1(n799), .A2(n798), .ZN(n526) );
  NOR2_X1 U579 ( .A1(n786), .A2(n799), .ZN(n527) );
  NOR2_X1 U580 ( .A1(n838), .A2(n835), .ZN(n528) );
  AND2_X1 U581 ( .A1(n583), .A2(n584), .ZN(G160) );
  XNOR2_X1 U582 ( .A(n533), .B(KEYINPUT106), .ZN(n850) );
  NAND2_X1 U583 ( .A1(n534), .A2(n528), .ZN(n533) );
  NAND2_X1 U584 ( .A1(n535), .A2(n526), .ZN(n534) );
  XNOR2_X1 U585 ( .A(n794), .B(KEYINPUT105), .ZN(n535) );
  NAND2_X1 U586 ( .A1(n539), .A2(n538), .ZN(n537) );
  INV_X1 U587 ( .A(n1002), .ZN(n538) );
  INV_X1 U588 ( .A(n1010), .ZN(n539) );
  INV_X1 U589 ( .A(G2104), .ZN(n559) );
  AND2_X1 U590 ( .A1(n765), .A2(n759), .ZN(n761) );
  NOR2_X1 U591 ( .A1(KEYINPUT33), .A2(n527), .ZN(n540) );
  XOR2_X1 U592 ( .A(G651), .B(KEYINPUT66), .Z(n541) );
  INV_X1 U593 ( .A(KEYINPUT99), .ZN(n750) );
  XNOR2_X1 U594 ( .A(n750), .B(KEYINPUT30), .ZN(n751) );
  XNOR2_X1 U595 ( .A(n752), .B(n751), .ZN(n753) );
  XNOR2_X1 U596 ( .A(n746), .B(n745), .ZN(n755) );
  NOR2_X1 U597 ( .A1(G1966), .A2(n799), .ZN(n747) );
  INV_X1 U598 ( .A(KEYINPUT101), .ZN(n760) );
  NOR2_X1 U599 ( .A1(n540), .A2(n788), .ZN(n789) );
  AND2_X1 U600 ( .A1(n790), .A2(n789), .ZN(n791) );
  INV_X1 U601 ( .A(KEYINPUT13), .ZN(n601) );
  XNOR2_X1 U602 ( .A(n542), .B(KEYINPUT1), .ZN(n543) );
  XNOR2_X1 U603 ( .A(n602), .B(n601), .ZN(n603) );
  XOR2_X1 U604 ( .A(KEYINPUT15), .B(n620), .Z(n1002) );
  NOR2_X1 U605 ( .A1(G651), .A2(n667), .ZN(n677) );
  INV_X1 U606 ( .A(KEYINPUT9), .ZN(n551) );
  NOR2_X1 U607 ( .A1(n564), .A2(n563), .ZN(G164) );
  XOR2_X1 U608 ( .A(KEYINPUT0), .B(G543), .Z(n667) );
  NAND2_X1 U609 ( .A1(n677), .A2(G52), .ZN(n546) );
  NOR2_X1 U610 ( .A1(G543), .A2(n541), .ZN(n544) );
  INV_X1 U611 ( .A(KEYINPUT68), .ZN(n542) );
  NAND2_X1 U612 ( .A1(G64), .A2(n612), .ZN(n545) );
  NAND2_X1 U613 ( .A1(n546), .A2(n545), .ZN(n554) );
  OR2_X1 U614 ( .A1(n667), .A2(n541), .ZN(n547) );
  NAND2_X1 U615 ( .A1(n523), .A2(G77), .ZN(n548) );
  XOR2_X1 U616 ( .A(KEYINPUT69), .B(n548), .Z(n550) );
  NOR2_X2 U617 ( .A1(G651), .A2(G543), .ZN(n675) );
  NAND2_X1 U618 ( .A1(n675), .A2(G90), .ZN(n549) );
  NAND2_X1 U619 ( .A1(n550), .A2(n549), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n552), .B(n551), .ZN(n553) );
  NOR2_X1 U621 ( .A1(n554), .A2(n553), .ZN(G171) );
  INV_X1 U622 ( .A(G171), .ZN(G301) );
  NAND2_X1 U623 ( .A1(n573), .A2(G102), .ZN(n557) );
  XOR2_X1 U624 ( .A(KEYINPUT85), .B(n555), .Z(n556) );
  NAND2_X1 U625 ( .A1(n557), .A2(n556), .ZN(n564) );
  NOR2_X1 U626 ( .A1(G2104), .A2(G2105), .ZN(n558) );
  XOR2_X1 U627 ( .A(KEYINPUT17), .B(n558), .Z(n590) );
  NAND2_X1 U628 ( .A1(G138), .A2(n590), .ZN(n562) );
  XNOR2_X2 U629 ( .A(n560), .B(KEYINPUT64), .ZN(n907) );
  NAND2_X1 U630 ( .A1(G126), .A2(n907), .ZN(n561) );
  NAND2_X1 U631 ( .A1(n562), .A2(n561), .ZN(n563) );
  NAND2_X1 U632 ( .A1(G85), .A2(n675), .ZN(n566) );
  NAND2_X1 U633 ( .A1(G60), .A2(n612), .ZN(n565) );
  NAND2_X1 U634 ( .A1(n566), .A2(n565), .ZN(n570) );
  NAND2_X1 U635 ( .A1(G72), .A2(n523), .ZN(n568) );
  NAND2_X1 U636 ( .A1(G47), .A2(n677), .ZN(n567) );
  NAND2_X1 U637 ( .A1(n568), .A2(n567), .ZN(n569) );
  OR2_X1 U638 ( .A1(n570), .A2(n569), .ZN(G290) );
  NAND2_X1 U639 ( .A1(G113), .A2(n906), .ZN(n572) );
  NAND2_X1 U640 ( .A1(G137), .A2(n590), .ZN(n571) );
  AND2_X1 U641 ( .A1(n572), .A2(n571), .ZN(n584) );
  INV_X1 U642 ( .A(KEYINPUT23), .ZN(n575) );
  NAND2_X1 U643 ( .A1(n573), .A2(G101), .ZN(n574) );
  XNOR2_X1 U644 ( .A(n575), .B(n574), .ZN(n577) );
  NAND2_X1 U645 ( .A1(n907), .A2(G125), .ZN(n576) );
  NAND2_X1 U646 ( .A1(n577), .A2(n576), .ZN(n580) );
  INV_X1 U647 ( .A(n580), .ZN(n579) );
  INV_X1 U648 ( .A(KEYINPUT65), .ZN(n578) );
  NAND2_X1 U649 ( .A1(n579), .A2(n578), .ZN(n582) );
  NAND2_X1 U650 ( .A1(n580), .A2(KEYINPUT65), .ZN(n581) );
  NAND2_X1 U651 ( .A1(n582), .A2(n581), .ZN(n583) );
  AND2_X1 U652 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U653 ( .A1(G111), .A2(n906), .ZN(n586) );
  NAND2_X1 U654 ( .A1(G99), .A2(n573), .ZN(n585) );
  NAND2_X1 U655 ( .A1(n586), .A2(n585), .ZN(n589) );
  NAND2_X1 U656 ( .A1(n907), .A2(G123), .ZN(n587) );
  XOR2_X1 U657 ( .A(KEYINPUT18), .B(n587), .Z(n588) );
  NOR2_X1 U658 ( .A1(n589), .A2(n588), .ZN(n592) );
  BUF_X1 U659 ( .A(n590), .Z(n910) );
  NAND2_X1 U660 ( .A1(n910), .A2(G135), .ZN(n591) );
  NAND2_X1 U661 ( .A1(n592), .A2(n591), .ZN(n955) );
  XNOR2_X1 U662 ( .A(G2096), .B(n955), .ZN(n593) );
  OR2_X1 U663 ( .A1(G2100), .A2(n593), .ZN(G156) );
  INV_X1 U664 ( .A(G132), .ZN(G219) );
  INV_X1 U665 ( .A(G82), .ZN(G220) );
  XOR2_X1 U666 ( .A(KEYINPUT73), .B(KEYINPUT10), .Z(n595) );
  NAND2_X1 U667 ( .A1(G7), .A2(G661), .ZN(n594) );
  XNOR2_X1 U668 ( .A(n595), .B(n594), .ZN(G223) );
  INV_X1 U669 ( .A(G223), .ZN(n863) );
  NAND2_X1 U670 ( .A1(n863), .A2(G567), .ZN(n596) );
  XOR2_X1 U671 ( .A(KEYINPUT11), .B(n596), .Z(G234) );
  NAND2_X1 U672 ( .A1(G56), .A2(n612), .ZN(n597) );
  XOR2_X1 U673 ( .A(KEYINPUT14), .B(n597), .Z(n604) );
  NAND2_X1 U674 ( .A1(n675), .A2(G81), .ZN(n598) );
  XNOR2_X1 U675 ( .A(n598), .B(KEYINPUT12), .ZN(n600) );
  NAND2_X1 U676 ( .A1(G68), .A2(n523), .ZN(n599) );
  NAND2_X1 U677 ( .A1(n600), .A2(n599), .ZN(n602) );
  NOR2_X1 U678 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X1 U679 ( .A(n605), .B(KEYINPUT74), .ZN(n607) );
  NAND2_X1 U680 ( .A1(G43), .A2(n677), .ZN(n606) );
  NAND2_X2 U681 ( .A1(n607), .A2(n606), .ZN(n1010) );
  INV_X1 U682 ( .A(G860), .ZN(n653) );
  OR2_X1 U683 ( .A1(n1010), .A2(n653), .ZN(G153) );
  INV_X1 U684 ( .A(G868), .ZN(n695) );
  NOR2_X1 U685 ( .A1(KEYINPUT75), .A2(G171), .ZN(n608) );
  NOR2_X1 U686 ( .A1(KEYINPUT77), .A2(n608), .ZN(n609) );
  NOR2_X1 U687 ( .A1(n695), .A2(n609), .ZN(n625) );
  NAND2_X1 U688 ( .A1(G301), .A2(G868), .ZN(n610) );
  NAND2_X1 U689 ( .A1(n610), .A2(KEYINPUT75), .ZN(n623) );
  NAND2_X1 U690 ( .A1(n677), .A2(G54), .ZN(n619) );
  NAND2_X1 U691 ( .A1(G79), .A2(n523), .ZN(n614) );
  NAND2_X1 U692 ( .A1(G66), .A2(n612), .ZN(n613) );
  NAND2_X1 U693 ( .A1(n614), .A2(n613), .ZN(n617) );
  NAND2_X1 U694 ( .A1(n675), .A2(G92), .ZN(n615) );
  XOR2_X1 U695 ( .A(KEYINPUT76), .B(n615), .Z(n616) );
  NOR2_X1 U696 ( .A1(n617), .A2(n616), .ZN(n618) );
  NAND2_X1 U697 ( .A1(n619), .A2(n618), .ZN(n620) );
  NOR2_X1 U698 ( .A1(n538), .A2(KEYINPUT77), .ZN(n621) );
  NAND2_X1 U699 ( .A1(n695), .A2(n621), .ZN(n622) );
  NAND2_X1 U700 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U701 ( .A1(n625), .A2(n624), .ZN(n627) );
  NAND2_X1 U702 ( .A1(n538), .A2(KEYINPUT77), .ZN(n626) );
  NAND2_X1 U703 ( .A1(n627), .A2(n626), .ZN(G284) );
  NAND2_X1 U704 ( .A1(n677), .A2(G53), .ZN(n629) );
  NAND2_X1 U705 ( .A1(G65), .A2(n612), .ZN(n628) );
  NAND2_X1 U706 ( .A1(n629), .A2(n628), .ZN(n633) );
  NAND2_X1 U707 ( .A1(G91), .A2(n675), .ZN(n631) );
  NAND2_X1 U708 ( .A1(G78), .A2(n523), .ZN(n630) );
  NAND2_X1 U709 ( .A1(n631), .A2(n630), .ZN(n632) );
  NOR2_X1 U710 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U711 ( .A(n634), .B(KEYINPUT70), .ZN(n991) );
  XNOR2_X1 U712 ( .A(KEYINPUT71), .B(n991), .ZN(G299) );
  NAND2_X1 U713 ( .A1(n675), .A2(G89), .ZN(n635) );
  XNOR2_X1 U714 ( .A(n635), .B(KEYINPUT4), .ZN(n637) );
  NAND2_X1 U715 ( .A1(G76), .A2(n523), .ZN(n636) );
  NAND2_X1 U716 ( .A1(n637), .A2(n636), .ZN(n638) );
  XNOR2_X1 U717 ( .A(n638), .B(KEYINPUT5), .ZN(n643) );
  NAND2_X1 U718 ( .A1(n677), .A2(G51), .ZN(n640) );
  NAND2_X1 U719 ( .A1(G63), .A2(n612), .ZN(n639) );
  NAND2_X1 U720 ( .A1(n640), .A2(n639), .ZN(n641) );
  XOR2_X1 U721 ( .A(KEYINPUT6), .B(n641), .Z(n642) );
  NAND2_X1 U722 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U723 ( .A(n644), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U724 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NOR2_X1 U725 ( .A1(G299), .A2(G868), .ZN(n646) );
  NOR2_X1 U726 ( .A1(G286), .A2(n695), .ZN(n645) );
  NOR2_X1 U727 ( .A1(n646), .A2(n645), .ZN(G297) );
  NAND2_X1 U728 ( .A1(n653), .A2(G559), .ZN(n647) );
  NAND2_X1 U729 ( .A1(n647), .A2(n538), .ZN(n648) );
  XNOR2_X1 U730 ( .A(n648), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U731 ( .A1(G868), .A2(n1010), .ZN(n651) );
  NAND2_X1 U732 ( .A1(G868), .A2(n538), .ZN(n649) );
  NOR2_X1 U733 ( .A1(G559), .A2(n649), .ZN(n650) );
  NOR2_X1 U734 ( .A1(n651), .A2(n650), .ZN(G282) );
  NAND2_X1 U735 ( .A1(G559), .A2(n538), .ZN(n652) );
  XOR2_X1 U736 ( .A(n1010), .B(n652), .Z(n692) );
  NAND2_X1 U737 ( .A1(n653), .A2(n692), .ZN(n660) );
  NAND2_X1 U738 ( .A1(G93), .A2(n675), .ZN(n655) );
  NAND2_X1 U739 ( .A1(G80), .A2(n523), .ZN(n654) );
  NAND2_X1 U740 ( .A1(n655), .A2(n654), .ZN(n659) );
  NAND2_X1 U741 ( .A1(n677), .A2(G55), .ZN(n657) );
  NAND2_X1 U742 ( .A1(G67), .A2(n612), .ZN(n656) );
  NAND2_X1 U743 ( .A1(n657), .A2(n656), .ZN(n658) );
  NOR2_X1 U744 ( .A1(n659), .A2(n658), .ZN(n694) );
  XOR2_X1 U745 ( .A(n660), .B(n694), .Z(G145) );
  NAND2_X1 U746 ( .A1(G88), .A2(n675), .ZN(n662) );
  NAND2_X1 U747 ( .A1(G75), .A2(n523), .ZN(n661) );
  NAND2_X1 U748 ( .A1(n662), .A2(n661), .ZN(n666) );
  NAND2_X1 U749 ( .A1(n677), .A2(G50), .ZN(n664) );
  NAND2_X1 U750 ( .A1(G62), .A2(n612), .ZN(n663) );
  NAND2_X1 U751 ( .A1(n664), .A2(n663), .ZN(n665) );
  NOR2_X1 U752 ( .A1(n666), .A2(n665), .ZN(G166) );
  NAND2_X1 U753 ( .A1(G74), .A2(G651), .ZN(n672) );
  NAND2_X1 U754 ( .A1(G49), .A2(n677), .ZN(n669) );
  NAND2_X1 U755 ( .A1(G87), .A2(n667), .ZN(n668) );
  NAND2_X1 U756 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U757 ( .A1(n612), .A2(n670), .ZN(n671) );
  NAND2_X1 U758 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U759 ( .A(n673), .B(KEYINPUT78), .ZN(G288) );
  NAND2_X1 U760 ( .A1(G73), .A2(n523), .ZN(n674) );
  XNOR2_X1 U761 ( .A(n674), .B(KEYINPUT2), .ZN(n684) );
  NAND2_X1 U762 ( .A1(n675), .A2(G86), .ZN(n676) );
  XNOR2_X1 U763 ( .A(n676), .B(KEYINPUT80), .ZN(n679) );
  NAND2_X1 U764 ( .A1(G48), .A2(n677), .ZN(n678) );
  NAND2_X1 U765 ( .A1(n679), .A2(n678), .ZN(n682) );
  NAND2_X1 U766 ( .A1(G61), .A2(n612), .ZN(n680) );
  XNOR2_X1 U767 ( .A(KEYINPUT79), .B(n680), .ZN(n681) );
  NOR2_X1 U768 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U769 ( .A1(n684), .A2(n683), .ZN(n685) );
  XOR2_X1 U770 ( .A(KEYINPUT81), .B(n685), .Z(G305) );
  XNOR2_X1 U771 ( .A(n694), .B(KEYINPUT82), .ZN(n686) );
  XNOR2_X1 U772 ( .A(n686), .B(KEYINPUT19), .ZN(n687) );
  XNOR2_X1 U773 ( .A(n687), .B(G290), .ZN(n690) );
  XOR2_X1 U774 ( .A(G166), .B(G288), .Z(n688) );
  XNOR2_X1 U775 ( .A(G299), .B(n688), .ZN(n689) );
  XNOR2_X1 U776 ( .A(n690), .B(n689), .ZN(n691) );
  XNOR2_X1 U777 ( .A(n691), .B(G305), .ZN(n933) );
  XOR2_X1 U778 ( .A(n933), .B(n692), .Z(n693) );
  NOR2_X1 U779 ( .A1(n695), .A2(n693), .ZN(n697) );
  AND2_X1 U780 ( .A1(n695), .A2(n694), .ZN(n696) );
  NOR2_X1 U781 ( .A1(n697), .A2(n696), .ZN(G295) );
  NAND2_X1 U782 ( .A1(G2084), .A2(G2078), .ZN(n698) );
  XOR2_X1 U783 ( .A(KEYINPUT20), .B(n698), .Z(n699) );
  NAND2_X1 U784 ( .A1(G2090), .A2(n699), .ZN(n701) );
  XOR2_X1 U785 ( .A(KEYINPUT21), .B(KEYINPUT83), .Z(n700) );
  XNOR2_X1 U786 ( .A(n701), .B(n700), .ZN(n702) );
  NAND2_X1 U787 ( .A1(G2072), .A2(n702), .ZN(G158) );
  XOR2_X1 U788 ( .A(KEYINPUT72), .B(G57), .Z(G237) );
  XNOR2_X1 U789 ( .A(KEYINPUT84), .B(G44), .ZN(n703) );
  XNOR2_X1 U790 ( .A(n703), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U791 ( .A1(G108), .A2(G120), .ZN(n704) );
  NOR2_X1 U792 ( .A1(G237), .A2(n704), .ZN(n705) );
  NAND2_X1 U793 ( .A1(G69), .A2(n705), .ZN(n867) );
  NAND2_X1 U794 ( .A1(n867), .A2(G567), .ZN(n710) );
  NOR2_X1 U795 ( .A1(G220), .A2(G219), .ZN(n706) );
  XOR2_X1 U796 ( .A(KEYINPUT22), .B(n706), .Z(n707) );
  NOR2_X1 U797 ( .A1(G218), .A2(n707), .ZN(n708) );
  NAND2_X1 U798 ( .A1(G96), .A2(n708), .ZN(n868) );
  NAND2_X1 U799 ( .A1(n868), .A2(G2106), .ZN(n709) );
  NAND2_X1 U800 ( .A1(n710), .A2(n709), .ZN(n869) );
  NAND2_X1 U801 ( .A1(G483), .A2(G661), .ZN(n711) );
  NOR2_X1 U802 ( .A1(n869), .A2(n711), .ZN(n866) );
  NAND2_X1 U803 ( .A1(n866), .A2(G36), .ZN(G176) );
  XOR2_X1 U804 ( .A(KEYINPUT86), .B(G166), .Z(G303) );
  NAND2_X1 U805 ( .A1(n739), .A2(G1996), .ZN(n714) );
  INV_X1 U806 ( .A(n714), .ZN(n713) );
  INV_X1 U807 ( .A(KEYINPUT26), .ZN(n712) );
  NAND2_X1 U808 ( .A1(n713), .A2(n712), .ZN(n716) );
  NAND2_X1 U809 ( .A1(n714), .A2(KEYINPUT26), .ZN(n715) );
  NAND2_X1 U810 ( .A1(n716), .A2(n715), .ZN(n718) );
  NAND2_X1 U811 ( .A1(G1341), .A2(n766), .ZN(n717) );
  NAND2_X1 U812 ( .A1(G1348), .A2(n766), .ZN(n720) );
  XNOR2_X2 U813 ( .A(n739), .B(KEYINPUT96), .ZN(n737) );
  NAND2_X1 U814 ( .A1(G2067), .A2(n737), .ZN(n719) );
  NAND2_X1 U815 ( .A1(n720), .A2(n719), .ZN(n721) );
  NAND2_X1 U816 ( .A1(n525), .A2(n721), .ZN(n725) );
  OR2_X1 U817 ( .A1(n1010), .A2(n722), .ZN(n723) );
  NAND2_X1 U818 ( .A1(n723), .A2(n1002), .ZN(n724) );
  NAND2_X1 U819 ( .A1(n725), .A2(n724), .ZN(n730) );
  NAND2_X1 U820 ( .A1(G2072), .A2(n737), .ZN(n726) );
  XNOR2_X1 U821 ( .A(n726), .B(KEYINPUT27), .ZN(n728) );
  INV_X1 U822 ( .A(G1956), .ZN(n1024) );
  NOR2_X1 U823 ( .A1(n737), .A2(n1024), .ZN(n727) );
  NOR2_X1 U824 ( .A1(n728), .A2(n727), .ZN(n731) );
  NAND2_X1 U825 ( .A1(n731), .A2(n991), .ZN(n729) );
  NAND2_X1 U826 ( .A1(n730), .A2(n729), .ZN(n734) );
  NOR2_X1 U827 ( .A1(n731), .A2(n991), .ZN(n732) );
  XOR2_X1 U828 ( .A(n732), .B(KEYINPUT28), .Z(n733) );
  NAND2_X1 U829 ( .A1(n734), .A2(n733), .ZN(n736) );
  XNOR2_X1 U830 ( .A(n736), .B(n735), .ZN(n743) );
  XNOR2_X1 U831 ( .A(G2078), .B(KEYINPUT25), .ZN(n976) );
  NAND2_X1 U832 ( .A1(n976), .A2(n737), .ZN(n738) );
  XNOR2_X1 U833 ( .A(n738), .B(KEYINPUT97), .ZN(n741) );
  NOR2_X1 U834 ( .A1(n739), .A2(G1961), .ZN(n740) );
  NOR2_X1 U835 ( .A1(n741), .A2(n740), .ZN(n744) );
  OR2_X1 U836 ( .A1(n744), .A2(G301), .ZN(n742) );
  NAND2_X1 U837 ( .A1(n743), .A2(n742), .ZN(n757) );
  NAND2_X1 U838 ( .A1(G301), .A2(n744), .ZN(n746) );
  NOR2_X1 U839 ( .A1(G2084), .A2(n766), .ZN(n762) );
  INV_X1 U840 ( .A(KEYINPUT95), .ZN(n748) );
  NAND2_X1 U841 ( .A1(G8), .A2(n766), .ZN(n799) );
  XNOR2_X1 U842 ( .A(n748), .B(n747), .ZN(n758) );
  NOR2_X1 U843 ( .A1(n762), .A2(n758), .ZN(n749) );
  NAND2_X1 U844 ( .A1(G8), .A2(n749), .ZN(n752) );
  NOR2_X1 U845 ( .A1(G168), .A2(n753), .ZN(n754) );
  NAND2_X1 U846 ( .A1(n757), .A2(n524), .ZN(n765) );
  INV_X1 U847 ( .A(n758), .ZN(n759) );
  XNOR2_X1 U848 ( .A(n761), .B(n760), .ZN(n764) );
  NAND2_X1 U849 ( .A1(G8), .A2(n762), .ZN(n763) );
  NAND2_X1 U850 ( .A1(n764), .A2(n763), .ZN(n775) );
  NAND2_X1 U851 ( .A1(n765), .A2(G286), .ZN(n771) );
  NOR2_X1 U852 ( .A1(G1971), .A2(n799), .ZN(n768) );
  NOR2_X1 U853 ( .A1(G2090), .A2(n766), .ZN(n767) );
  NOR2_X1 U854 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U855 ( .A1(G303), .A2(n769), .ZN(n770) );
  NAND2_X1 U856 ( .A1(n771), .A2(n770), .ZN(n772) );
  NAND2_X1 U857 ( .A1(n772), .A2(G8), .ZN(n773) );
  XNOR2_X1 U858 ( .A(n773), .B(KEYINPUT32), .ZN(n774) );
  NAND2_X1 U859 ( .A1(n775), .A2(n774), .ZN(n776) );
  XNOR2_X1 U860 ( .A(n776), .B(KEYINPUT102), .ZN(n785) );
  NOR2_X1 U861 ( .A1(G2090), .A2(G303), .ZN(n777) );
  NAND2_X1 U862 ( .A1(G8), .A2(n777), .ZN(n778) );
  NAND2_X1 U863 ( .A1(n785), .A2(n778), .ZN(n779) );
  XNOR2_X1 U864 ( .A(n779), .B(KEYINPUT104), .ZN(n780) );
  NAND2_X1 U865 ( .A1(n780), .A2(n799), .ZN(n793) );
  XOR2_X1 U866 ( .A(G1981), .B(G305), .Z(n1007) );
  NOR2_X1 U867 ( .A1(G1976), .A2(G288), .ZN(n992) );
  NOR2_X1 U868 ( .A1(G303), .A2(G1971), .ZN(n997) );
  NOR2_X1 U869 ( .A1(n992), .A2(n997), .ZN(n781) );
  XOR2_X1 U870 ( .A(KEYINPUT103), .B(n781), .Z(n783) );
  INV_X1 U871 ( .A(KEYINPUT33), .ZN(n782) );
  AND2_X1 U872 ( .A1(n783), .A2(n782), .ZN(n784) );
  NAND2_X1 U873 ( .A1(n785), .A2(n784), .ZN(n790) );
  NAND2_X1 U874 ( .A1(G1976), .A2(G288), .ZN(n996) );
  INV_X1 U875 ( .A(n996), .ZN(n786) );
  NAND2_X1 U876 ( .A1(n992), .A2(KEYINPUT33), .ZN(n787) );
  NOR2_X1 U877 ( .A1(n787), .A2(n799), .ZN(n788) );
  NAND2_X1 U878 ( .A1(n1007), .A2(n791), .ZN(n792) );
  NAND2_X1 U879 ( .A1(n793), .A2(n792), .ZN(n794) );
  XNOR2_X1 U880 ( .A(KEYINPUT93), .B(KEYINPUT24), .ZN(n795) );
  XNOR2_X1 U881 ( .A(n795), .B(KEYINPUT94), .ZN(n797) );
  NOR2_X1 U882 ( .A1(G1981), .A2(G305), .ZN(n796) );
  XNOR2_X1 U883 ( .A(n797), .B(n796), .ZN(n798) );
  INV_X1 U884 ( .A(n800), .ZN(n802) );
  NOR2_X1 U885 ( .A1(n802), .A2(n801), .ZN(n803) );
  XNOR2_X1 U886 ( .A(n803), .B(KEYINPUT87), .ZN(n834) );
  INV_X1 U887 ( .A(n834), .ZN(n847) );
  NAND2_X1 U888 ( .A1(G131), .A2(n910), .ZN(n805) );
  NAND2_X1 U889 ( .A1(G119), .A2(n907), .ZN(n804) );
  NAND2_X1 U890 ( .A1(n805), .A2(n804), .ZN(n809) );
  NAND2_X1 U891 ( .A1(G107), .A2(n906), .ZN(n807) );
  NAND2_X1 U892 ( .A1(G95), .A2(n573), .ZN(n806) );
  NAND2_X1 U893 ( .A1(n807), .A2(n806), .ZN(n808) );
  NOR2_X1 U894 ( .A1(n809), .A2(n808), .ZN(n810) );
  XNOR2_X1 U895 ( .A(n810), .B(KEYINPUT89), .ZN(n919) );
  NAND2_X1 U896 ( .A1(G1991), .A2(n919), .ZN(n811) );
  XNOR2_X1 U897 ( .A(n811), .B(KEYINPUT90), .ZN(n821) );
  NAND2_X1 U898 ( .A1(G117), .A2(n906), .ZN(n813) );
  NAND2_X1 U899 ( .A1(G129), .A2(n907), .ZN(n812) );
  NAND2_X1 U900 ( .A1(n813), .A2(n812), .ZN(n816) );
  NAND2_X1 U901 ( .A1(n573), .A2(G105), .ZN(n814) );
  XOR2_X1 U902 ( .A(KEYINPUT38), .B(n814), .Z(n815) );
  NOR2_X1 U903 ( .A1(n816), .A2(n815), .ZN(n817) );
  XOR2_X1 U904 ( .A(KEYINPUT91), .B(n817), .Z(n819) );
  NAND2_X1 U905 ( .A1(n910), .A2(G141), .ZN(n818) );
  NAND2_X1 U906 ( .A1(n819), .A2(n818), .ZN(n928) );
  NAND2_X1 U907 ( .A1(G1996), .A2(n928), .ZN(n820) );
  NAND2_X1 U908 ( .A1(n821), .A2(n820), .ZN(n822) );
  XNOR2_X1 U909 ( .A(KEYINPUT92), .B(n822), .ZN(n965) );
  AND2_X1 U910 ( .A1(n847), .A2(n965), .ZN(n838) );
  XNOR2_X1 U911 ( .A(G1986), .B(G290), .ZN(n1004) );
  XNOR2_X1 U912 ( .A(G2067), .B(KEYINPUT37), .ZN(n844) );
  NAND2_X1 U913 ( .A1(G104), .A2(n573), .ZN(n824) );
  NAND2_X1 U914 ( .A1(G140), .A2(n910), .ZN(n823) );
  NAND2_X1 U915 ( .A1(n824), .A2(n823), .ZN(n825) );
  XNOR2_X1 U916 ( .A(KEYINPUT34), .B(n825), .ZN(n831) );
  NAND2_X1 U917 ( .A1(G116), .A2(n906), .ZN(n827) );
  NAND2_X1 U918 ( .A1(G128), .A2(n907), .ZN(n826) );
  NAND2_X1 U919 ( .A1(n827), .A2(n826), .ZN(n828) );
  XOR2_X1 U920 ( .A(KEYINPUT88), .B(n828), .Z(n829) );
  XNOR2_X1 U921 ( .A(KEYINPUT35), .B(n829), .ZN(n830) );
  NOR2_X1 U922 ( .A1(n831), .A2(n830), .ZN(n832) );
  XNOR2_X1 U923 ( .A(KEYINPUT36), .B(n832), .ZN(n918) );
  NOR2_X1 U924 ( .A1(n844), .A2(n918), .ZN(n952) );
  NOR2_X1 U925 ( .A1(n1004), .A2(n952), .ZN(n833) );
  NOR2_X1 U926 ( .A1(n834), .A2(n833), .ZN(n835) );
  XOR2_X1 U927 ( .A(KEYINPUT107), .B(KEYINPUT39), .Z(n841) );
  NOR2_X1 U928 ( .A1(G1996), .A2(n928), .ZN(n944) );
  NOR2_X1 U929 ( .A1(G1991), .A2(n919), .ZN(n958) );
  NOR2_X1 U930 ( .A1(G1986), .A2(G290), .ZN(n836) );
  NOR2_X1 U931 ( .A1(n958), .A2(n836), .ZN(n837) );
  NOR2_X1 U932 ( .A1(n838), .A2(n837), .ZN(n839) );
  NOR2_X1 U933 ( .A1(n944), .A2(n839), .ZN(n840) );
  XNOR2_X1 U934 ( .A(n841), .B(n840), .ZN(n843) );
  INV_X1 U935 ( .A(n952), .ZN(n842) );
  NAND2_X1 U936 ( .A1(n843), .A2(n842), .ZN(n845) );
  NAND2_X1 U937 ( .A1(n844), .A2(n918), .ZN(n953) );
  NAND2_X1 U938 ( .A1(n845), .A2(n953), .ZN(n846) );
  XNOR2_X1 U939 ( .A(KEYINPUT108), .B(n846), .ZN(n848) );
  NAND2_X1 U940 ( .A1(n848), .A2(n847), .ZN(n849) );
  NAND2_X1 U941 ( .A1(n850), .A2(n849), .ZN(n851) );
  XNOR2_X1 U942 ( .A(n851), .B(KEYINPUT40), .ZN(G329) );
  XNOR2_X1 U943 ( .A(G2446), .B(G2454), .ZN(n861) );
  XOR2_X1 U944 ( .A(G2430), .B(KEYINPUT110), .Z(n853) );
  XNOR2_X1 U945 ( .A(G2451), .B(G2443), .ZN(n852) );
  XNOR2_X1 U946 ( .A(n853), .B(n852), .ZN(n857) );
  XOR2_X1 U947 ( .A(G2427), .B(KEYINPUT109), .Z(n855) );
  XNOR2_X1 U948 ( .A(G1341), .B(G1348), .ZN(n854) );
  XNOR2_X1 U949 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U950 ( .A(n857), .B(n856), .Z(n859) );
  XNOR2_X1 U951 ( .A(G2438), .B(G2435), .ZN(n858) );
  XNOR2_X1 U952 ( .A(n859), .B(n858), .ZN(n860) );
  XNOR2_X1 U953 ( .A(n861), .B(n860), .ZN(n862) );
  NAND2_X1 U954 ( .A1(n862), .A2(G14), .ZN(n937) );
  XNOR2_X1 U955 ( .A(KEYINPUT111), .B(n937), .ZN(G401) );
  NAND2_X1 U956 ( .A1(G2106), .A2(n863), .ZN(G217) );
  AND2_X1 U957 ( .A1(G15), .A2(G2), .ZN(n864) );
  NAND2_X1 U958 ( .A1(G661), .A2(n864), .ZN(G259) );
  NAND2_X1 U959 ( .A1(G3), .A2(G1), .ZN(n865) );
  NAND2_X1 U960 ( .A1(n866), .A2(n865), .ZN(G188) );
  INV_X1 U962 ( .A(G120), .ZN(G236) );
  INV_X1 U963 ( .A(G108), .ZN(G238) );
  INV_X1 U964 ( .A(G96), .ZN(G221) );
  INV_X1 U965 ( .A(G69), .ZN(G235) );
  NOR2_X1 U966 ( .A1(n868), .A2(n867), .ZN(G325) );
  INV_X1 U967 ( .A(G325), .ZN(G261) );
  INV_X1 U968 ( .A(n869), .ZN(G319) );
  XOR2_X1 U969 ( .A(KEYINPUT113), .B(KEYINPUT112), .Z(n871) );
  XNOR2_X1 U970 ( .A(G2678), .B(KEYINPUT43), .ZN(n870) );
  XNOR2_X1 U971 ( .A(n871), .B(n870), .ZN(n875) );
  XOR2_X1 U972 ( .A(KEYINPUT42), .B(G2072), .Z(n873) );
  XNOR2_X1 U973 ( .A(G2067), .B(G2090), .ZN(n872) );
  XNOR2_X1 U974 ( .A(n873), .B(n872), .ZN(n874) );
  XOR2_X1 U975 ( .A(n875), .B(n874), .Z(n877) );
  XNOR2_X1 U976 ( .A(G2096), .B(G2100), .ZN(n876) );
  XNOR2_X1 U977 ( .A(n877), .B(n876), .ZN(n879) );
  XOR2_X1 U978 ( .A(G2084), .B(G2078), .Z(n878) );
  XNOR2_X1 U979 ( .A(n879), .B(n878), .ZN(G227) );
  XOR2_X1 U980 ( .A(G1976), .B(G1971), .Z(n881) );
  XNOR2_X1 U981 ( .A(G1986), .B(G1956), .ZN(n880) );
  XNOR2_X1 U982 ( .A(n881), .B(n880), .ZN(n882) );
  XOR2_X1 U983 ( .A(n882), .B(KEYINPUT41), .Z(n884) );
  XNOR2_X1 U984 ( .A(G1996), .B(G1991), .ZN(n883) );
  XNOR2_X1 U985 ( .A(n884), .B(n883), .ZN(n888) );
  XOR2_X1 U986 ( .A(G2474), .B(G1961), .Z(n886) );
  XNOR2_X1 U987 ( .A(G1981), .B(G1966), .ZN(n885) );
  XNOR2_X1 U988 ( .A(n886), .B(n885), .ZN(n887) );
  XNOR2_X1 U989 ( .A(n888), .B(n887), .ZN(G229) );
  NAND2_X1 U990 ( .A1(G112), .A2(n906), .ZN(n890) );
  NAND2_X1 U991 ( .A1(G100), .A2(n573), .ZN(n889) );
  NAND2_X1 U992 ( .A1(n890), .A2(n889), .ZN(n897) );
  NAND2_X1 U993 ( .A1(n907), .A2(G124), .ZN(n891) );
  XNOR2_X1 U994 ( .A(n891), .B(KEYINPUT114), .ZN(n892) );
  XNOR2_X1 U995 ( .A(KEYINPUT44), .B(n892), .ZN(n895) );
  NAND2_X1 U996 ( .A1(G136), .A2(n910), .ZN(n893) );
  XOR2_X1 U997 ( .A(KEYINPUT115), .B(n893), .Z(n894) );
  NAND2_X1 U998 ( .A1(n895), .A2(n894), .ZN(n896) );
  NOR2_X1 U999 ( .A1(n897), .A2(n896), .ZN(G162) );
  NAND2_X1 U1000 ( .A1(G115), .A2(n906), .ZN(n899) );
  NAND2_X1 U1001 ( .A1(G127), .A2(n907), .ZN(n898) );
  NAND2_X1 U1002 ( .A1(n899), .A2(n898), .ZN(n900) );
  XNOR2_X1 U1003 ( .A(n900), .B(KEYINPUT47), .ZN(n902) );
  NAND2_X1 U1004 ( .A1(G103), .A2(n573), .ZN(n901) );
  NAND2_X1 U1005 ( .A1(n902), .A2(n901), .ZN(n905) );
  NAND2_X1 U1006 ( .A1(n910), .A2(G139), .ZN(n903) );
  XOR2_X1 U1007 ( .A(KEYINPUT116), .B(n903), .Z(n904) );
  NOR2_X1 U1008 ( .A1(n905), .A2(n904), .ZN(n946) );
  NAND2_X1 U1009 ( .A1(G118), .A2(n906), .ZN(n909) );
  NAND2_X1 U1010 ( .A1(G130), .A2(n907), .ZN(n908) );
  NAND2_X1 U1011 ( .A1(n909), .A2(n908), .ZN(n915) );
  NAND2_X1 U1012 ( .A1(G106), .A2(n573), .ZN(n912) );
  NAND2_X1 U1013 ( .A1(G142), .A2(n910), .ZN(n911) );
  NAND2_X1 U1014 ( .A1(n912), .A2(n911), .ZN(n913) );
  XOR2_X1 U1015 ( .A(KEYINPUT45), .B(n913), .Z(n914) );
  NOR2_X1 U1016 ( .A1(n915), .A2(n914), .ZN(n916) );
  XOR2_X1 U1017 ( .A(n946), .B(n916), .Z(n917) );
  XNOR2_X1 U1018 ( .A(n918), .B(n917), .ZN(n922) );
  XNOR2_X1 U1019 ( .A(G162), .B(n919), .ZN(n920) );
  XNOR2_X1 U1020 ( .A(n920), .B(n955), .ZN(n921) );
  XOR2_X1 U1021 ( .A(n922), .B(n921), .Z(n927) );
  XOR2_X1 U1022 ( .A(KEYINPUT117), .B(KEYINPUT48), .Z(n924) );
  XNOR2_X1 U1023 ( .A(KEYINPUT118), .B(KEYINPUT46), .ZN(n923) );
  XNOR2_X1 U1024 ( .A(n924), .B(n923), .ZN(n925) );
  XNOR2_X1 U1025 ( .A(G164), .B(n925), .ZN(n926) );
  XNOR2_X1 U1026 ( .A(n927), .B(n926), .ZN(n930) );
  XOR2_X1 U1027 ( .A(n928), .B(G160), .Z(n929) );
  XNOR2_X1 U1028 ( .A(n930), .B(n929), .ZN(n931) );
  NOR2_X1 U1029 ( .A1(G37), .A2(n931), .ZN(G395) );
  XNOR2_X1 U1030 ( .A(G286), .B(G301), .ZN(n932) );
  XNOR2_X1 U1031 ( .A(n932), .B(n1002), .ZN(n935) );
  XOR2_X1 U1032 ( .A(n1010), .B(n933), .Z(n934) );
  XNOR2_X1 U1033 ( .A(n935), .B(n934), .ZN(n936) );
  NOR2_X1 U1034 ( .A1(G37), .A2(n936), .ZN(G397) );
  NAND2_X1 U1035 ( .A1(G319), .A2(n937), .ZN(n940) );
  NOR2_X1 U1036 ( .A1(G227), .A2(G229), .ZN(n938) );
  XNOR2_X1 U1037 ( .A(KEYINPUT49), .B(n938), .ZN(n939) );
  NOR2_X1 U1038 ( .A1(n940), .A2(n939), .ZN(n942) );
  NOR2_X1 U1039 ( .A1(G395), .A2(G397), .ZN(n941) );
  NAND2_X1 U1040 ( .A1(n942), .A2(n941), .ZN(G225) );
  INV_X1 U1041 ( .A(G225), .ZN(G308) );
  XOR2_X1 U1042 ( .A(G2090), .B(G162), .Z(n943) );
  NOR2_X1 U1043 ( .A1(n944), .A2(n943), .ZN(n945) );
  XOR2_X1 U1044 ( .A(KEYINPUT51), .B(n945), .Z(n963) );
  XNOR2_X1 U1045 ( .A(G2072), .B(n946), .ZN(n949) );
  XNOR2_X1 U1046 ( .A(G164), .B(G2078), .ZN(n947) );
  XNOR2_X1 U1047 ( .A(n947), .B(KEYINPUT120), .ZN(n948) );
  NAND2_X1 U1048 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1049 ( .A(n950), .B(KEYINPUT50), .ZN(n951) );
  NOR2_X1 U1050 ( .A1(n952), .A2(n951), .ZN(n954) );
  NAND2_X1 U1051 ( .A1(n954), .A2(n953), .ZN(n961) );
  XNOR2_X1 U1052 ( .A(G160), .B(G2084), .ZN(n956) );
  NAND2_X1 U1053 ( .A1(n956), .A2(n955), .ZN(n957) );
  NOR2_X1 U1054 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1055 ( .A(KEYINPUT119), .B(n959), .ZN(n960) );
  NOR2_X1 U1056 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1057 ( .A1(n963), .A2(n962), .ZN(n964) );
  NOR2_X1 U1058 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1059 ( .A(KEYINPUT52), .B(n966), .ZN(n967) );
  INV_X1 U1060 ( .A(KEYINPUT55), .ZN(n987) );
  NAND2_X1 U1061 ( .A1(n967), .A2(n987), .ZN(n968) );
  NAND2_X1 U1062 ( .A1(n968), .A2(G29), .ZN(n1050) );
  XNOR2_X1 U1063 ( .A(G2090), .B(G35), .ZN(n981) );
  XNOR2_X1 U1064 ( .A(G2067), .B(G26), .ZN(n970) );
  XNOR2_X1 U1065 ( .A(G33), .B(G2072), .ZN(n969) );
  NOR2_X1 U1066 ( .A1(n970), .A2(n969), .ZN(n975) );
  XOR2_X1 U1067 ( .A(G1991), .B(G25), .Z(n971) );
  NAND2_X1 U1068 ( .A1(n971), .A2(G28), .ZN(n973) );
  XNOR2_X1 U1069 ( .A(G32), .B(G1996), .ZN(n972) );
  NOR2_X1 U1070 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1071 ( .A1(n975), .A2(n974), .ZN(n978) );
  XOR2_X1 U1072 ( .A(G27), .B(n976), .Z(n977) );
  NOR2_X1 U1073 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1074 ( .A(KEYINPUT53), .B(n979), .ZN(n980) );
  NOR2_X1 U1075 ( .A1(n981), .A2(n980), .ZN(n982) );
  XOR2_X1 U1076 ( .A(KEYINPUT121), .B(n982), .Z(n985) );
  XOR2_X1 U1077 ( .A(KEYINPUT54), .B(G34), .Z(n983) );
  XNOR2_X1 U1078 ( .A(G2084), .B(n983), .ZN(n984) );
  NAND2_X1 U1079 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1080 ( .A(n987), .B(n986), .ZN(n989) );
  INV_X1 U1081 ( .A(G29), .ZN(n988) );
  NAND2_X1 U1082 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1083 ( .A1(G11), .A2(n990), .ZN(n1048) );
  XNOR2_X1 U1084 ( .A(G16), .B(KEYINPUT56), .ZN(n1018) );
  XOR2_X1 U1085 ( .A(n991), .B(G1956), .Z(n994) );
  XNOR2_X1 U1086 ( .A(n992), .B(KEYINPUT122), .ZN(n993) );
  NOR2_X1 U1087 ( .A1(n994), .A2(n993), .ZN(n1000) );
  NAND2_X1 U1088 ( .A1(G303), .A2(G1971), .ZN(n995) );
  NAND2_X1 U1089 ( .A1(n996), .A2(n995), .ZN(n998) );
  NOR2_X1 U1090 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1091 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1092 ( .A(KEYINPUT123), .B(n1001), .ZN(n1016) );
  XNOR2_X1 U1093 ( .A(G171), .B(G1961), .ZN(n1006) );
  XNOR2_X1 U1094 ( .A(G1348), .B(n1002), .ZN(n1003) );
  NOR2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1014) );
  XNOR2_X1 U1097 ( .A(G1966), .B(G168), .ZN(n1008) );
  NAND2_X1 U1098 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1099 ( .A(n1009), .B(KEYINPUT57), .ZN(n1012) );
  XOR2_X1 U1100 ( .A(G1341), .B(n1010), .Z(n1011) );
  NAND2_X1 U1101 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NOR2_X1 U1102 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1046) );
  INV_X1 U1105 ( .A(G16), .ZN(n1044) );
  XOR2_X1 U1106 ( .A(G1986), .B(G24), .Z(n1020) );
  XOR2_X1 U1107 ( .A(G1971), .B(G22), .Z(n1019) );
  NAND2_X1 U1108 ( .A1(n1020), .A2(n1019), .ZN(n1022) );
  XNOR2_X1 U1109 ( .A(G23), .B(G1976), .ZN(n1021) );
  NOR2_X1 U1110 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XOR2_X1 U1111 ( .A(KEYINPUT58), .B(n1023), .Z(n1041) );
  XNOR2_X1 U1112 ( .A(G1961), .B(G5), .ZN(n1038) );
  XOR2_X1 U1113 ( .A(G1981), .B(G6), .Z(n1026) );
  XNOR2_X1 U1114 ( .A(n1024), .B(G20), .ZN(n1025) );
  NAND2_X1 U1115 ( .A1(n1026), .A2(n1025), .ZN(n1032) );
  XOR2_X1 U1116 ( .A(G1341), .B(G19), .Z(n1030) );
  XNOR2_X1 U1117 ( .A(KEYINPUT59), .B(G4), .ZN(n1027) );
  XNOR2_X1 U1118 ( .A(n1027), .B(KEYINPUT124), .ZN(n1028) );
  XNOR2_X1 U1119 ( .A(G1348), .B(n1028), .ZN(n1029) );
  NAND2_X1 U1120 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NOR2_X1 U1121 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XOR2_X1 U1122 ( .A(KEYINPUT60), .B(n1033), .Z(n1035) );
  XNOR2_X1 U1123 ( .A(G1966), .B(G21), .ZN(n1034) );
  NOR2_X1 U1124 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  XNOR2_X1 U1125 ( .A(KEYINPUT125), .B(n1036), .ZN(n1037) );
  NOR2_X1 U1126 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  XOR2_X1 U1127 ( .A(KEYINPUT126), .B(n1039), .Z(n1040) );
  NOR2_X1 U1128 ( .A1(n1041), .A2(n1040), .ZN(n1042) );
  XNOR2_X1 U1129 ( .A(KEYINPUT61), .B(n1042), .ZN(n1043) );
  NAND2_X1 U1130 ( .A1(n1044), .A2(n1043), .ZN(n1045) );
  NAND2_X1 U1131 ( .A1(n1046), .A2(n1045), .ZN(n1047) );
  NOR2_X1 U1132 ( .A1(n1048), .A2(n1047), .ZN(n1049) );
  NAND2_X1 U1133 ( .A1(n1050), .A2(n1049), .ZN(n1051) );
  XOR2_X1 U1134 ( .A(KEYINPUT62), .B(n1051), .Z(G311) );
  INV_X1 U1135 ( .A(G311), .ZN(G150) );
endmodule

