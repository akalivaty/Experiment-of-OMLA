//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 1 0 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 1 0 0 0 1 1 1 0 0 0 0 1 1 1 1 1 1 0 0 0 0 1 0 0 1 1 1 0 1 0 1 0 0 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:46 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n586, new_n587, new_n588, new_n589,
    new_n590, new_n591, new_n592, new_n593, new_n594, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n620, new_n621, new_n622, new_n623, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n644, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949;
  INV_X1    g000(.A(KEYINPUT6), .ZN(new_n187));
  XNOR2_X1  g001(.A(G116), .B(G119), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(KEYINPUT5), .ZN(new_n189));
  INV_X1    g003(.A(G119), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G116), .ZN(new_n191));
  OAI211_X1 g005(.A(new_n189), .B(G113), .C1(KEYINPUT5), .C2(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT2), .B(G113), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(new_n188), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n192), .A2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT3), .ZN(new_n197));
  INV_X1    g011(.A(G104), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n197), .B1(new_n198), .B2(G107), .ZN(new_n199));
  INV_X1    g013(.A(G107), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n200), .A2(KEYINPUT3), .A3(G104), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n199), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G101), .ZN(new_n203));
  OAI21_X1  g017(.A(KEYINPUT71), .B1(new_n200), .B2(G104), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT71), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n205), .A2(new_n198), .A3(G107), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n202), .A2(new_n203), .A3(new_n204), .A4(new_n206), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n198), .A2(G107), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n200), .A2(G104), .ZN(new_n209));
  OAI21_X1  g023(.A(G101), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n207), .A2(new_n210), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n196), .A2(new_n211), .ZN(new_n212));
  AND3_X1   g026(.A1(new_n200), .A2(KEYINPUT3), .A3(G104), .ZN(new_n213));
  AOI21_X1  g027(.A(KEYINPUT3), .B1(new_n200), .B2(G104), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n204), .A2(new_n206), .ZN(new_n216));
  OAI21_X1  g030(.A(KEYINPUT72), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT72), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n202), .A2(new_n218), .A3(new_n204), .A4(new_n206), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n217), .A2(G101), .A3(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT73), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n207), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n217), .A2(new_n221), .A3(G101), .A4(new_n219), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n223), .A2(KEYINPUT4), .A3(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT4), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n217), .A2(new_n226), .A3(G101), .A4(new_n219), .ZN(new_n227));
  OR2_X1    g041(.A1(new_n194), .A2(new_n188), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(new_n195), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n212), .B1(new_n225), .B2(new_n231), .ZN(new_n232));
  XNOR2_X1  g046(.A(G110), .B(G122), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n187), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n233), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT75), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n235), .B1(new_n232), .B2(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n226), .B1(new_n220), .B2(new_n222), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n230), .B1(new_n238), .B2(new_n224), .ZN(new_n239));
  NOR3_X1   g053(.A1(new_n239), .A2(KEYINPUT75), .A3(new_n212), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n234), .B1(new_n237), .B2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G146), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G143), .ZN(new_n243));
  INV_X1    g057(.A(G143), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G146), .ZN(new_n245));
  AND2_X1   g059(.A1(KEYINPUT0), .A2(G128), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n243), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  XNOR2_X1  g061(.A(G143), .B(G146), .ZN(new_n248));
  XNOR2_X1  g062(.A(KEYINPUT0), .B(G128), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n247), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G125), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n243), .A2(new_n245), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n243), .A2(KEYINPUT1), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n254), .A2(new_n255), .A3(G128), .ZN(new_n256));
  INV_X1    g070(.A(G128), .ZN(new_n257));
  OAI211_X1 g071(.A(new_n243), .B(new_n245), .C1(KEYINPUT1), .C2(new_n257), .ZN(new_n258));
  AOI21_X1  g072(.A(G125), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n253), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(G953), .ZN(new_n261));
  AND2_X1   g075(.A1(new_n261), .A2(G224), .ZN(new_n262));
  XOR2_X1   g076(.A(new_n260), .B(new_n262), .Z(new_n263));
  NAND2_X1  g077(.A1(new_n232), .A2(new_n236), .ZN(new_n264));
  OAI21_X1  g078(.A(KEYINPUT75), .B1(new_n239), .B2(new_n212), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n264), .A2(new_n265), .A3(new_n187), .A4(new_n235), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n241), .A2(new_n263), .A3(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT79), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT7), .ZN(new_n269));
  OAI22_X1  g083(.A1(new_n253), .A2(new_n259), .B1(new_n269), .B2(new_n262), .ZN(new_n270));
  INV_X1    g084(.A(new_n259), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n262), .A2(new_n269), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n271), .B(new_n272), .C1(new_n252), .C2(new_n251), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n211), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n275), .A2(KEYINPUT76), .A3(new_n195), .A4(new_n192), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT76), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n277), .B1(new_n196), .B2(new_n211), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n196), .A2(new_n211), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n276), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n233), .B(KEYINPUT8), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n274), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  OR2_X1    g096(.A1(new_n282), .A2(KEYINPUT77), .ZN(new_n283));
  AOI22_X1  g097(.A1(new_n282), .A2(KEYINPUT77), .B1(new_n232), .B2(new_n233), .ZN(new_n284));
  AOI21_X1  g098(.A(G902), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n267), .A2(new_n268), .A3(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(G210), .B1(G237), .B2(G902), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(KEYINPUT78), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n286), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n267), .A2(new_n285), .A3(new_n287), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(KEYINPUT79), .ZN(new_n293));
  NAND4_X1  g107(.A1(new_n267), .A2(new_n268), .A3(new_n285), .A4(new_n289), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n291), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(G214), .B1(G237), .B2(G902), .ZN(new_n296));
  XNOR2_X1  g110(.A(KEYINPUT9), .B(G234), .ZN(new_n297));
  OAI21_X1  g111(.A(G221), .B1(new_n297), .B2(G902), .ZN(new_n298));
  XOR2_X1   g112(.A(new_n298), .B(KEYINPUT70), .Z(new_n299));
  INV_X1    g113(.A(G469), .ZN(new_n300));
  INV_X1    g114(.A(G902), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  XNOR2_X1  g116(.A(G110), .B(G140), .ZN(new_n303));
  AND2_X1   g117(.A1(new_n261), .A2(G227), .ZN(new_n304));
  XNOR2_X1  g118(.A(new_n303), .B(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT11), .ZN(new_n306));
  INV_X1    g120(.A(G134), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n306), .B1(new_n307), .B2(G137), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(G137), .ZN(new_n309));
  INV_X1    g123(.A(G137), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n310), .A2(KEYINPUT11), .A3(G134), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n308), .A2(new_n309), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G131), .ZN(new_n313));
  INV_X1    g127(.A(G131), .ZN(new_n314));
  NAND4_X1  g128(.A1(new_n308), .A2(new_n311), .A3(new_n314), .A4(new_n309), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n227), .A2(new_n251), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n225), .A2(new_n319), .ZN(new_n320));
  NAND4_X1  g134(.A1(new_n207), .A2(new_n258), .A3(new_n256), .A4(new_n210), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT10), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n321), .B(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n317), .B1(new_n320), .B2(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n318), .B1(new_n238), .B2(new_n224), .ZN(new_n326));
  NOR3_X1   g140(.A1(new_n326), .A2(new_n316), .A3(new_n323), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n305), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n320), .A2(new_n317), .A3(new_n324), .ZN(new_n329));
  AOI22_X1  g143(.A1(new_n207), .A2(new_n210), .B1(new_n256), .B2(new_n258), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT74), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n330), .B1(new_n331), .B2(new_n321), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n256), .A2(new_n258), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n211), .A2(new_n331), .A3(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n316), .B1(new_n332), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(KEYINPUT12), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT12), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n338), .B(new_n316), .C1(new_n332), .C2(new_n335), .ZN(new_n339));
  INV_X1    g153(.A(new_n305), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n329), .A2(new_n337), .A3(new_n339), .A4(new_n340), .ZN(new_n341));
  AOI21_X1  g155(.A(G902), .B1(new_n328), .B2(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n302), .B1(new_n342), .B2(new_n300), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n337), .A2(new_n339), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n305), .B1(new_n344), .B2(new_n327), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n316), .B1(new_n326), .B2(new_n323), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n329), .A2(new_n346), .A3(new_n340), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n345), .A2(G469), .A3(new_n347), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n299), .B1(new_n343), .B2(new_n348), .ZN(new_n349));
  XNOR2_X1  g163(.A(G113), .B(G122), .ZN(new_n350));
  XNOR2_X1  g164(.A(KEYINPUT80), .B(G104), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n350), .B(new_n351), .ZN(new_n352));
  NOR3_X1   g166(.A1(new_n252), .A2(KEYINPUT16), .A3(G140), .ZN(new_n353));
  XNOR2_X1  g167(.A(G125), .B(G140), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n353), .B1(new_n354), .B2(KEYINPUT16), .ZN(new_n355));
  AND2_X1   g169(.A1(new_n355), .A2(G146), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n355), .A2(G146), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(G237), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n359), .A2(new_n261), .A3(G214), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n360), .B(new_n244), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n361), .A2(KEYINPUT17), .A3(G131), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(G131), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n360), .B(G143), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(new_n314), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  OAI211_X1 g180(.A(new_n358), .B(new_n362), .C1(new_n366), .C2(KEYINPUT17), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT18), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n364), .B1(new_n368), .B2(new_n314), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n361), .A2(KEYINPUT18), .A3(G131), .ZN(new_n370));
  XNOR2_X1  g184(.A(new_n354), .B(new_n242), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n369), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n352), .B1(new_n367), .B2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT17), .ZN(new_n374));
  AND3_X1   g188(.A1(new_n363), .A2(new_n365), .A3(new_n374), .ZN(new_n375));
  OR2_X1    g189(.A1(new_n355), .A2(G146), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n355), .A2(G146), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n376), .A2(new_n362), .A3(new_n377), .ZN(new_n378));
  OAI211_X1 g192(.A(new_n372), .B(new_n352), .C1(new_n375), .C2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n301), .B1(new_n373), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(G475), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n354), .B(KEYINPUT19), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(new_n242), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n366), .A2(new_n377), .A3(new_n384), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n352), .B1(new_n385), .B2(new_n372), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n380), .A2(new_n386), .ZN(new_n387));
  NOR2_X1   g201(.A1(G475), .A2(G902), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  NOR3_X1   g203(.A1(new_n387), .A2(KEYINPUT20), .A3(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT20), .ZN(new_n391));
  AND2_X1   g205(.A1(new_n385), .A2(new_n372), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n379), .B1(new_n392), .B2(new_n352), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n391), .B1(new_n393), .B2(new_n388), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n382), .B1(new_n390), .B2(new_n394), .ZN(new_n395));
  XNOR2_X1  g209(.A(G128), .B(G143), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(new_n307), .ZN(new_n397));
  XNOR2_X1  g211(.A(G116), .B(G122), .ZN(new_n398));
  XNOR2_X1  g212(.A(new_n398), .B(new_n200), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT13), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n400), .B1(new_n257), .B2(G143), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n244), .A2(KEYINPUT13), .A3(G128), .ZN(new_n402));
  OAI211_X1 g216(.A(new_n401), .B(new_n402), .C1(G128), .C2(new_n244), .ZN(new_n403));
  AND3_X1   g217(.A1(new_n403), .A2(KEYINPUT81), .A3(G134), .ZN(new_n404));
  AOI21_X1  g218(.A(KEYINPUT81), .B1(new_n403), .B2(G134), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n397), .B(new_n399), .C1(new_n404), .C2(new_n405), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n396), .B(new_n307), .ZN(new_n407));
  INV_X1    g221(.A(G116), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n408), .A2(KEYINPUT14), .A3(G122), .ZN(new_n409));
  INV_X1    g223(.A(new_n398), .ZN(new_n410));
  OAI211_X1 g224(.A(G107), .B(new_n409), .C1(new_n410), .C2(KEYINPUT14), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n407), .B(new_n411), .C1(G107), .C2(new_n410), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n406), .A2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(G217), .ZN(new_n414));
  NOR3_X1   g228(.A1(new_n297), .A2(new_n414), .A3(G953), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n406), .A2(new_n412), .A3(new_n415), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT82), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n419), .A2(new_n420), .A3(new_n301), .ZN(new_n421));
  INV_X1    g235(.A(G478), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n422), .A2(KEYINPUT15), .ZN(new_n423));
  OR2_X1    g237(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n421), .A2(new_n423), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(G234), .A2(G237), .ZN(new_n427));
  AND3_X1   g241(.A1(new_n427), .A2(G952), .A3(new_n261), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  XOR2_X1   g243(.A(KEYINPUT21), .B(G898), .Z(new_n430));
  XNOR2_X1  g244(.A(new_n430), .B(KEYINPUT83), .ZN(new_n431));
  AND3_X1   g245(.A1(new_n427), .A2(G902), .A3(G953), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n429), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  NOR3_X1   g249(.A1(new_n395), .A2(new_n426), .A3(new_n435), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n295), .A2(new_n296), .A3(new_n349), .A4(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT28), .ZN(new_n438));
  AND3_X1   g252(.A1(new_n316), .A2(KEYINPUT64), .A3(new_n251), .ZN(new_n439));
  AOI21_X1  g253(.A(KEYINPUT64), .B1(new_n316), .B2(new_n251), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n307), .A2(G137), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n310), .A2(G134), .ZN(new_n443));
  OAI21_X1  g257(.A(G131), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND4_X1  g258(.A1(new_n256), .A2(new_n315), .A3(new_n258), .A4(new_n444), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n445), .B(KEYINPUT65), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n229), .B1(new_n441), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n316), .A2(new_n251), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(KEYINPUT66), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT66), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n316), .A2(new_n450), .A3(new_n251), .ZN(new_n451));
  INV_X1    g265(.A(new_n229), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n449), .A2(new_n451), .A3(new_n452), .A4(new_n445), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n438), .B1(new_n447), .B2(new_n453), .ZN(new_n454));
  AND2_X1   g268(.A1(new_n452), .A2(new_n445), .ZN(new_n455));
  AOI21_X1  g269(.A(KEYINPUT28), .B1(new_n455), .B2(new_n448), .ZN(new_n456));
  XOR2_X1   g270(.A(KEYINPUT67), .B(KEYINPUT27), .Z(new_n457));
  NAND3_X1  g271(.A1(new_n359), .A2(new_n261), .A3(G210), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n457), .B(new_n458), .ZN(new_n459));
  XNOR2_X1  g273(.A(KEYINPUT26), .B(G101), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n459), .B(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  NOR3_X1   g276(.A1(new_n454), .A2(new_n456), .A3(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT30), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n464), .B1(new_n441), .B2(new_n446), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n449), .A2(new_n451), .A3(KEYINPUT30), .A4(new_n445), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n465), .A2(new_n229), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n461), .B1(new_n467), .B2(new_n453), .ZN(new_n468));
  NOR3_X1   g282(.A1(new_n463), .A2(new_n468), .A3(KEYINPUT29), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n449), .A2(new_n451), .A3(new_n445), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(new_n229), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n438), .B1(new_n471), .B2(new_n453), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n472), .A2(new_n456), .ZN(new_n473));
  AND2_X1   g287(.A1(new_n461), .A2(KEYINPUT29), .ZN(new_n474));
  AOI21_X1  g288(.A(G902), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(G472), .B1(new_n469), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n467), .A2(new_n453), .A3(new_n461), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(KEYINPUT31), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n462), .B1(new_n454), .B2(new_n456), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT31), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n467), .A2(new_n481), .A3(new_n453), .A4(new_n461), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n479), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT32), .ZN(new_n484));
  NOR2_X1   g298(.A1(G472), .A2(G902), .ZN(new_n485));
  AND3_X1   g299(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n484), .B1(new_n483), .B2(new_n485), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n477), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  XNOR2_X1  g302(.A(KEYINPUT22), .B(G137), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n261), .A2(G221), .A3(G234), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n489), .B(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n190), .A2(G128), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n257), .A2(KEYINPUT23), .A3(G119), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n190), .A2(G128), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n492), .B(new_n493), .C1(new_n494), .C2(KEYINPUT23), .ZN(new_n495));
  XOR2_X1   g309(.A(KEYINPUT24), .B(G110), .Z(new_n496));
  XNOR2_X1  g310(.A(G119), .B(G128), .ZN(new_n497));
  AOI22_X1  g311(.A1(new_n495), .A2(G110), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n498), .B1(new_n356), .B2(new_n357), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT69), .ZN(new_n500));
  XOR2_X1   g314(.A(KEYINPUT68), .B(G110), .Z(new_n501));
  OAI22_X1  g315(.A1(new_n495), .A2(new_n501), .B1(new_n496), .B2(new_n497), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n354), .A2(new_n242), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n502), .A2(new_n377), .A3(new_n503), .ZN(new_n504));
  AND3_X1   g318(.A1(new_n499), .A2(new_n500), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n500), .B1(new_n499), .B2(new_n504), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n491), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n491), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n499), .A2(new_n504), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n508), .B1(new_n509), .B2(KEYINPUT69), .ZN(new_n510));
  AND2_X1   g324(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n511), .A2(KEYINPUT25), .A3(new_n301), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n507), .A2(new_n301), .A3(new_n510), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT25), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n414), .B1(G234), .B2(new_n301), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n517), .A2(G902), .ZN(new_n518));
  AOI22_X1  g332(.A1(new_n516), .A2(new_n517), .B1(new_n511), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n488), .A2(new_n519), .ZN(new_n520));
  OR2_X1    g334(.A1(new_n437), .A2(new_n520), .ZN(new_n521));
  XNOR2_X1  g335(.A(KEYINPUT84), .B(G101), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n521), .B(new_n522), .ZN(G3));
  NAND2_X1  g337(.A1(new_n483), .A2(new_n301), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(G472), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n483), .A2(new_n485), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n328), .A2(new_n341), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n528), .A2(new_n300), .A3(new_n301), .ZN(new_n529));
  INV_X1    g343(.A(new_n302), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n529), .A2(new_n530), .A3(new_n348), .ZN(new_n531));
  INV_X1    g345(.A(new_n299), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n519), .ZN(new_n534));
  NOR3_X1   g348(.A1(new_n527), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  XOR2_X1   g349(.A(new_n535), .B(KEYINPUT85), .Z(new_n536));
  INV_X1    g350(.A(new_n395), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT33), .ZN(new_n538));
  AOI21_X1  g352(.A(KEYINPUT86), .B1(new_n406), .B2(new_n412), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n419), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n539), .A2(new_n538), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n541), .A2(new_n418), .A3(new_n417), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n422), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n419), .A2(new_n422), .A3(new_n301), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n544), .B1(new_n422), .B2(new_n301), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  NOR3_X1   g361(.A1(new_n537), .A2(new_n547), .A3(new_n435), .ZN(new_n548));
  AND3_X1   g362(.A1(new_n267), .A2(new_n285), .A3(new_n287), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n287), .B1(new_n267), .B2(new_n285), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n548), .B(new_n296), .C1(new_n549), .C2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n536), .A2(new_n552), .ZN(new_n553));
  XOR2_X1   g367(.A(KEYINPUT34), .B(G104), .Z(new_n554));
  XNOR2_X1  g368(.A(new_n553), .B(new_n554), .ZN(G6));
  INV_X1    g369(.A(new_n296), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n267), .A2(new_n285), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(new_n288), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n556), .B1(new_n558), .B2(new_n292), .ZN(new_n559));
  AOI22_X1  g373(.A1(new_n424), .A2(new_n425), .B1(G475), .B2(new_n381), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT87), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n394), .A2(new_n561), .ZN(new_n562));
  OAI21_X1  g376(.A(KEYINPUT20), .B1(new_n387), .B2(new_n389), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n393), .A2(new_n391), .A3(new_n388), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n563), .A2(KEYINPUT87), .A3(new_n564), .ZN(new_n565));
  AND4_X1   g379(.A1(new_n434), .A2(new_n560), .A3(new_n562), .A4(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n559), .A2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n536), .A2(new_n568), .ZN(new_n569));
  XOR2_X1   g383(.A(KEYINPUT35), .B(G107), .Z(new_n570));
  XNOR2_X1  g384(.A(new_n569), .B(new_n570), .ZN(G9));
  NAND2_X1  g385(.A1(new_n516), .A2(new_n517), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT36), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n491), .A2(new_n573), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n574), .B(KEYINPUT88), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT89), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n575), .B(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n577), .B(new_n509), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(new_n518), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n572), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n525), .A2(new_n526), .A3(new_n580), .ZN(new_n581));
  OR2_X1    g395(.A1(new_n437), .A2(new_n581), .ZN(new_n582));
  XNOR2_X1  g396(.A(KEYINPUT37), .B(G110), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n583), .B(KEYINPUT90), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n582), .B(new_n584), .ZN(G12));
  AND4_X1   g399(.A1(new_n488), .A2(new_n559), .A3(new_n349), .A4(new_n580), .ZN(new_n586));
  AND2_X1   g400(.A1(new_n565), .A2(new_n562), .ZN(new_n587));
  XOR2_X1   g401(.A(new_n428), .B(KEYINPUT91), .Z(new_n588));
  OAI21_X1  g402(.A(new_n588), .B1(G900), .B2(new_n433), .ZN(new_n589));
  XOR2_X1   g403(.A(new_n589), .B(KEYINPUT92), .Z(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n587), .A2(new_n560), .A3(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n586), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n594), .B(G128), .ZN(G30));
  XOR2_X1   g409(.A(KEYINPUT96), .B(KEYINPUT39), .Z(new_n596));
  XNOR2_X1  g410(.A(new_n590), .B(new_n596), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n533), .A2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT40), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NOR3_X1   g414(.A1(new_n533), .A2(KEYINPUT40), .A3(new_n597), .ZN(new_n601));
  INV_X1    g415(.A(new_n426), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n537), .A2(new_n602), .ZN(new_n603));
  AOI22_X1  g417(.A1(new_n516), .A2(new_n517), .B1(new_n578), .B2(new_n518), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n603), .A2(new_n604), .A3(new_n296), .ZN(new_n605));
  OR3_X1    g419(.A1(new_n600), .A2(new_n601), .A3(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(KEYINPUT93), .B(KEYINPUT38), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n295), .B(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n462), .B1(new_n467), .B2(new_n453), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n471), .A2(new_n453), .A3(new_n462), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(new_n301), .ZN(new_n612));
  OAI21_X1  g426(.A(G472), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT94), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n615), .B1(new_n486), .B2(new_n487), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(KEYINPUT95), .ZN(new_n617));
  NOR3_X1   g431(.A1(new_n606), .A2(new_n609), .A3(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(new_n244), .ZN(G45));
  NAND4_X1  g433(.A1(new_n488), .A2(new_n559), .A3(new_n349), .A4(new_n580), .ZN(new_n620));
  AND3_X1   g434(.A1(new_n395), .A2(new_n546), .A3(new_n591), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(new_n242), .ZN(G48));
  INV_X1    g438(.A(G472), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n468), .A2(KEYINPUT29), .ZN(new_n626));
  INV_X1    g440(.A(new_n463), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n625), .B1(new_n628), .B2(new_n475), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n526), .A2(KEYINPUT32), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n629), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n632), .A2(new_n534), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n342), .A2(new_n300), .ZN(new_n634));
  AOI211_X1 g448(.A(G469), .B(G902), .C1(new_n328), .C2(new_n341), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n634), .A2(new_n635), .A3(new_n299), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n552), .A2(new_n633), .A3(KEYINPUT97), .A4(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT97), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n488), .A2(new_n519), .A3(new_n636), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n638), .B1(new_n639), .B2(new_n551), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(KEYINPUT41), .B(G113), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G15));
  NAND3_X1  g457(.A1(new_n633), .A2(new_n568), .A3(new_n636), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(G116), .ZN(G18));
  NAND3_X1  g459(.A1(new_n488), .A2(new_n436), .A3(new_n580), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n559), .A2(new_n636), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(new_n190), .ZN(G21));
  OAI21_X1  g463(.A(new_n462), .B1(new_n472), .B2(new_n456), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n479), .A2(new_n482), .A3(new_n650), .ZN(new_n651));
  AOI22_X1  g465(.A1(new_n524), .A2(G472), .B1(new_n485), .B2(new_n651), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n652), .A2(new_n636), .A3(new_n519), .A4(new_n434), .ZN(new_n653));
  OAI211_X1 g467(.A(new_n603), .B(new_n296), .C1(new_n549), .C2(new_n550), .ZN(new_n654));
  OR2_X1    g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(G122), .ZN(G24));
  NAND2_X1  g470(.A1(new_n651), .A2(new_n485), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n625), .B1(new_n483), .B2(new_n301), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n658), .A2(new_n659), .A3(new_n604), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n660), .A2(new_n559), .A3(new_n621), .A4(new_n636), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G125), .ZN(G27));
  OAI21_X1  g476(.A(KEYINPUT99), .B1(new_n632), .B2(new_n534), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n291), .A2(new_n293), .A3(new_n296), .A4(new_n294), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT98), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n665), .B1(new_n345), .B2(new_n347), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n347), .A2(new_n665), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  NOR3_X1   g482(.A1(new_n666), .A2(new_n668), .A3(new_n300), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n529), .A2(new_n530), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n532), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n664), .A2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT99), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n488), .A2(new_n673), .A3(new_n519), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n663), .A2(new_n672), .A3(new_n621), .A4(new_n674), .ZN(new_n675));
  AND2_X1   g489(.A1(new_n345), .A2(new_n347), .ZN(new_n676));
  OAI211_X1 g490(.A(G469), .B(new_n667), .C1(new_n676), .C2(new_n665), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n299), .B1(new_n677), .B2(new_n343), .ZN(new_n678));
  AOI22_X1  g492(.A1(KEYINPUT79), .A2(new_n292), .B1(new_n286), .B2(new_n290), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n678), .A2(new_n679), .A3(new_n296), .A4(new_n294), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n680), .A2(new_n520), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n622), .A2(KEYINPUT42), .ZN(new_n682));
  AOI22_X1  g496(.A1(new_n675), .A2(KEYINPUT42), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G131), .ZN(G33));
  NAND3_X1  g498(.A1(new_n672), .A2(new_n633), .A3(new_n593), .ZN(new_n685));
  XNOR2_X1  g499(.A(KEYINPUT100), .B(G134), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(G36));
  OAI21_X1  g501(.A(G469), .B1(new_n676), .B2(KEYINPUT45), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n666), .A2(new_n668), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n688), .B1(KEYINPUT45), .B2(new_n689), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n690), .A2(new_n302), .ZN(new_n691));
  AND2_X1   g505(.A1(new_n691), .A2(KEYINPUT46), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n529), .B1(new_n691), .B2(KEYINPUT46), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n532), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  OR2_X1    g508(.A1(new_n694), .A2(new_n597), .ZN(new_n695));
  OR3_X1    g509(.A1(new_n547), .A2(KEYINPUT43), .A3(new_n395), .ZN(new_n696));
  OAI21_X1  g510(.A(KEYINPUT43), .B1(new_n547), .B2(new_n395), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n527), .A2(new_n580), .A3(new_n696), .A4(new_n697), .ZN(new_n698));
  XOR2_X1   g512(.A(new_n698), .B(KEYINPUT44), .Z(new_n699));
  OR3_X1    g513(.A1(new_n695), .A2(new_n664), .A3(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(KEYINPUT101), .B(G137), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(G39));
  INV_X1    g516(.A(KEYINPUT47), .ZN(new_n703));
  OR2_X1    g517(.A1(new_n694), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n694), .A2(new_n703), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NOR4_X1   g520(.A1(new_n664), .A2(new_n488), .A3(new_n519), .A4(new_n622), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G140), .ZN(G42));
  INV_X1    g523(.A(new_n588), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n696), .A2(new_n710), .A3(new_n697), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(KEYINPUT109), .ZN(new_n712));
  NOR3_X1   g526(.A1(new_n534), .A2(new_n658), .A3(new_n659), .ZN(new_n713));
  AND2_X1   g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n636), .A2(new_n556), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(KEYINPUT110), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n714), .A2(new_n609), .A3(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT50), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(KEYINPUT111), .ZN(new_n719));
  INV_X1    g533(.A(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n717), .B(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(KEYINPUT112), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n634), .A2(new_n635), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(new_n532), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n664), .A2(new_n724), .ZN(new_n725));
  AND2_X1   g539(.A1(new_n712), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(new_n660), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n617), .A2(new_n519), .A3(new_n428), .A4(new_n725), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n537), .A2(new_n547), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n727), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(new_n723), .ZN(new_n731));
  OAI211_X1 g545(.A(new_n704), .B(new_n705), .C1(new_n532), .C2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n664), .ZN(new_n733));
  AND2_X1   g547(.A1(new_n714), .A2(new_n733), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n730), .B1(new_n732), .B2(new_n734), .ZN(new_n735));
  AOI21_X1  g549(.A(KEYINPUT51), .B1(new_n722), .B2(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n735), .A2(new_n721), .A3(KEYINPUT51), .ZN(new_n737));
  AND2_X1   g551(.A1(new_n663), .A2(new_n674), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n726), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(KEYINPUT48), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n537), .A2(new_n547), .ZN(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  OR2_X1    g556(.A1(new_n728), .A2(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(G952), .ZN(new_n744));
  INV_X1    g558(.A(new_n647), .ZN(new_n745));
  AOI211_X1 g559(.A(new_n744), .B(G953), .C1(new_n714), .C2(new_n745), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n737), .A2(new_n740), .A3(new_n743), .A4(new_n746), .ZN(new_n747));
  OR2_X1    g561(.A1(new_n736), .A2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT52), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT105), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n604), .A2(new_n591), .ZN(new_n751));
  INV_X1    g565(.A(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n616), .A2(new_n678), .A3(new_n752), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n750), .B1(new_n753), .B2(new_n654), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n671), .A2(new_n751), .ZN(new_n755));
  INV_X1    g569(.A(new_n654), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n755), .A2(new_n756), .A3(KEYINPUT105), .A4(new_n616), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n632), .A2(new_n604), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n759), .A2(new_n349), .A3(new_n559), .A4(new_n621), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n525), .A2(new_n580), .A3(new_n621), .A4(new_n657), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n296), .B1(new_n549), .B2(new_n550), .ZN(new_n762));
  NOR3_X1   g576(.A1(new_n761), .A2(new_n724), .A3(new_n762), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n763), .B1(new_n586), .B2(new_n593), .ZN(new_n764));
  AND4_X1   g578(.A1(new_n749), .A2(new_n758), .A3(new_n760), .A4(new_n764), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n661), .B1(new_n620), .B2(new_n592), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n766), .A2(new_n623), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n749), .B1(new_n767), .B2(new_n758), .ZN(new_n768));
  OAI21_X1  g582(.A(KEYINPUT107), .B1(new_n765), .B2(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(new_n758), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n594), .A2(new_n760), .A3(new_n661), .ZN(new_n771));
  OAI21_X1  g585(.A(KEYINPUT52), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT107), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n767), .A2(new_n749), .A3(new_n758), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n772), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n769), .A2(new_n775), .ZN(new_n776));
  AND4_X1   g590(.A1(new_n382), .A2(new_n587), .A3(new_n602), .A4(new_n591), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n488), .A2(new_n777), .A3(new_n349), .A4(new_n580), .ZN(new_n778));
  OAI22_X1  g592(.A1(new_n778), .A2(new_n664), .B1(new_n680), .B2(new_n761), .ZN(new_n779));
  NOR3_X1   g593(.A1(new_n680), .A2(new_n520), .A3(new_n592), .ZN(new_n780));
  OAI21_X1  g594(.A(KEYINPUT104), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  OR2_X1    g595(.A1(new_n778), .A2(new_n664), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT104), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n672), .A2(new_n621), .A3(new_n660), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n782), .A2(new_n685), .A3(new_n783), .A4(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n781), .A2(new_n785), .ZN(new_n786));
  OAI22_X1  g600(.A1(new_n639), .A2(new_n567), .B1(new_n653), .B2(new_n654), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n787), .A2(new_n648), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n641), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n786), .A2(new_n789), .A3(new_n683), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n295), .A2(new_n296), .A3(new_n548), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(KEYINPUT102), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT102), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n295), .A2(new_n793), .A3(new_n296), .A4(new_n548), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n792), .A2(new_n535), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(new_n521), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(KEYINPUT103), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT103), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n795), .A2(new_n521), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n537), .A2(new_n426), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n800), .A2(new_n435), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n535), .A2(new_n296), .A3(new_n295), .A4(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n582), .A2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n797), .A2(new_n799), .A3(new_n804), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n790), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g620(.A(KEYINPUT53), .B1(new_n776), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n675), .A2(KEYINPUT42), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n681), .A2(new_n682), .ZN(new_n809));
  AND4_X1   g623(.A1(new_n641), .A2(new_n808), .A3(new_n809), .A4(new_n788), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n803), .B1(new_n796), .B2(KEYINPUT103), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n810), .A2(new_n799), .A3(new_n811), .A4(new_n786), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT53), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n772), .A2(new_n774), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n812), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n807), .A2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT54), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n776), .A2(new_n806), .ZN(new_n819));
  OAI21_X1  g633(.A(KEYINPUT108), .B1(new_n819), .B2(new_n813), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n812), .B1(new_n769), .B2(new_n775), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT108), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n821), .A2(new_n822), .A3(KEYINPUT53), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n813), .B1(new_n812), .B2(new_n814), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT106), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  OAI211_X1 g640(.A(KEYINPUT106), .B(new_n813), .C1(new_n812), .C2(new_n814), .ZN(new_n827));
  AOI22_X1  g641(.A1(new_n820), .A2(new_n823), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n818), .B1(new_n828), .B2(new_n817), .ZN(new_n829));
  OAI22_X1  g643(.A1(new_n748), .A2(new_n829), .B1(G952), .B2(G953), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n731), .A2(KEYINPUT49), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n731), .A2(KEYINPUT49), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n537), .A2(new_n296), .A3(new_n532), .A4(new_n546), .ZN(new_n833));
  NOR4_X1   g647(.A1(new_n831), .A2(new_n832), .A3(new_n534), .A4(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n609), .A2(new_n834), .A3(new_n617), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n830), .A2(new_n835), .ZN(G75));
  NOR2_X1   g650(.A1(new_n816), .A2(new_n301), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(G210), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n241), .A2(new_n266), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n839), .B(new_n263), .ZN(new_n840));
  XNOR2_X1  g654(.A(KEYINPUT113), .B(KEYINPUT55), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n841), .B(KEYINPUT114), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n840), .B(new_n842), .ZN(new_n843));
  XOR2_X1   g657(.A(KEYINPUT116), .B(KEYINPUT56), .Z(new_n844));
  NOR2_X1   g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n838), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n744), .A2(G953), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(KEYINPUT117), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT115), .ZN(new_n850));
  AOI21_X1  g664(.A(KEYINPUT56), .B1(new_n838), .B2(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n837), .A2(KEYINPUT115), .A3(G210), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n849), .B1(new_n853), .B2(new_n843), .ZN(G51));
  INV_X1    g668(.A(new_n848), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n302), .B(KEYINPUT57), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n819), .A2(new_n813), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT118), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n806), .A2(KEYINPUT53), .A3(new_n772), .A4(new_n774), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n857), .A2(new_n858), .A3(new_n817), .A4(new_n859), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n860), .B1(new_n817), .B2(new_n816), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n858), .B1(new_n816), .B2(new_n817), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n856), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(new_n528), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n837), .A2(new_n690), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n855), .B1(new_n864), .B2(new_n865), .ZN(G54));
  AND2_X1   g680(.A1(KEYINPUT58), .A2(G475), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n393), .A2(new_n867), .ZN(new_n868));
  OAI211_X1 g682(.A(G902), .B(new_n868), .C1(new_n807), .C2(new_n815), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT119), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n859), .B1(new_n821), .B2(KEYINPUT53), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n872), .A2(KEYINPUT119), .A3(G902), .A4(new_n868), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  OAI211_X1 g688(.A(G902), .B(new_n867), .C1(new_n807), .C2(new_n815), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n875), .A2(KEYINPUT120), .A3(new_n387), .ZN(new_n876));
  AOI21_X1  g690(.A(KEYINPUT120), .B1(new_n875), .B2(new_n387), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n874), .B(new_n848), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n878), .A2(KEYINPUT121), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n855), .B1(new_n871), .B2(new_n873), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT121), .ZN(new_n881));
  OAI211_X1 g695(.A(new_n880), .B(new_n881), .C1(new_n877), .C2(new_n876), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n879), .A2(new_n882), .ZN(G60));
  AND2_X1   g697(.A1(new_n540), .A2(new_n542), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n422), .A2(new_n301), .ZN(new_n885));
  XOR2_X1   g699(.A(new_n885), .B(KEYINPUT59), .Z(new_n886));
  OAI211_X1 g700(.A(new_n884), .B(new_n886), .C1(new_n861), .C2(new_n862), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(new_n848), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n884), .B1(new_n829), .B2(new_n886), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n888), .A2(new_n889), .ZN(G63));
  INV_X1    g704(.A(KEYINPUT61), .ZN(new_n891));
  XNOR2_X1  g705(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n414), .A2(new_n301), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n892), .B(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n872), .A2(new_n578), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(KEYINPUT123), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n872), .A2(new_n894), .ZN(new_n897));
  INV_X1    g711(.A(new_n511), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n896), .A2(new_n848), .A3(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n895), .A2(KEYINPUT123), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n891), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT124), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n899), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n897), .A2(KEYINPUT124), .A3(new_n898), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n855), .A2(new_n891), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n904), .A2(new_n895), .A3(new_n905), .A4(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n902), .A2(new_n907), .ZN(G66));
  AOI21_X1  g722(.A(new_n261), .B1(new_n431), .B2(G224), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n811), .A2(new_n799), .A3(new_n789), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n909), .B1(new_n910), .B2(new_n261), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n839), .B1(G898), .B2(new_n261), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n911), .B(new_n912), .Z(G69));
  INV_X1    g727(.A(new_n465), .ZN(new_n914));
  INV_X1    g728(.A(new_n466), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(KEYINPUT125), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(new_n383), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n918), .B1(G900), .B2(G953), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n738), .A2(new_n756), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n685), .B1(new_n695), .B2(new_n920), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n921), .A2(new_n771), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n922), .A2(new_n683), .A3(new_n700), .A4(new_n708), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n919), .B1(new_n923), .B2(G953), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n742), .A2(new_n800), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n633), .A2(new_n733), .A3(new_n598), .A4(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n700), .A2(new_n708), .A3(new_n926), .ZN(new_n927));
  OAI21_X1  g741(.A(KEYINPUT62), .B1(new_n618), .B2(new_n771), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT127), .ZN(new_n929));
  NOR3_X1   g743(.A1(new_n618), .A2(KEYINPUT62), .A3(new_n771), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n927), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n931), .A2(G953), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n918), .B(KEYINPUT126), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n924), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n261), .B1(G227), .B2(G900), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n934), .B(new_n935), .ZN(G72));
  NAND2_X1  g750(.A1(G472), .A2(G902), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(KEYINPUT63), .Z(new_n938));
  OAI21_X1  g752(.A(new_n938), .B1(new_n923), .B2(new_n910), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n467), .A2(new_n453), .A3(new_n462), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n855), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(new_n938), .ZN(new_n943));
  INV_X1    g757(.A(new_n910), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n943), .B1(new_n931), .B2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n610), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n942), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(new_n828), .ZN(new_n948));
  NOR3_X1   g762(.A1(new_n941), .A2(new_n610), .A3(new_n943), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n947), .B1(new_n948), .B2(new_n949), .ZN(G57));
endmodule


