//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 0 1 0 1 1 0 0 1 1 1 1 0 0 0 0 0 0 0 0 0 0 0 0 1 0 1 1 1 0 1 1 1 1 0 1 0 1 1 0 1 0 0 0 0 1 1 1 0 1 1 0 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:35 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005;
  INV_X1    g000(.A(G140), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G125), .ZN(new_n188));
  INV_X1    g002(.A(G125), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G140), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n188), .A2(new_n190), .A3(KEYINPUT16), .ZN(new_n191));
  OR3_X1    g005(.A1(new_n189), .A2(KEYINPUT16), .A3(G140), .ZN(new_n192));
  AND3_X1   g006(.A1(new_n191), .A2(G146), .A3(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G146), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n188), .A2(new_n190), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n193), .B1(new_n194), .B2(new_n196), .ZN(new_n197));
  OR2_X1    g011(.A1(KEYINPUT68), .A2(G128), .ZN(new_n198));
  NAND2_X1  g012(.A1(KEYINPUT68), .A2(G128), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n198), .A2(G119), .A3(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT79), .ZN(new_n201));
  INV_X1    g015(.A(G128), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n201), .B1(new_n202), .B2(G119), .ZN(new_n203));
  INV_X1    g017(.A(G119), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n204), .A2(KEYINPUT79), .A3(G128), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n200), .A2(new_n203), .A3(new_n205), .ZN(new_n206));
  XNOR2_X1  g020(.A(KEYINPUT24), .B(G110), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  AOI21_X1  g022(.A(KEYINPUT23), .B1(new_n202), .B2(G119), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n209), .B1(new_n204), .B2(G128), .ZN(new_n210));
  INV_X1    g024(.A(G110), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n198), .A2(KEYINPUT23), .A3(G119), .A4(new_n199), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n210), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  AND3_X1   g027(.A1(new_n208), .A2(new_n213), .A3(KEYINPUT81), .ZN(new_n214));
  AOI21_X1  g028(.A(KEYINPUT81), .B1(new_n208), .B2(new_n213), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n197), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  AOI21_X1  g030(.A(G146), .B1(new_n191), .B2(new_n192), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n193), .A2(new_n217), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n206), .A2(new_n207), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n211), .B1(new_n210), .B2(new_n212), .ZN(new_n220));
  NOR4_X1   g034(.A1(new_n218), .A2(new_n219), .A3(new_n220), .A4(KEYINPUT80), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT80), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n219), .A2(new_n220), .ZN(new_n223));
  OR2_X1    g037(.A1(new_n193), .A2(new_n217), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n222), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n216), .B1(new_n221), .B2(new_n225), .ZN(new_n226));
  AND2_X1   g040(.A1(KEYINPUT73), .A2(G953), .ZN(new_n227));
  NOR2_X1   g041(.A1(KEYINPUT73), .A2(G953), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n229), .A2(G221), .A3(G234), .ZN(new_n230));
  XNOR2_X1  g044(.A(KEYINPUT22), .B(G137), .ZN(new_n231));
  XNOR2_X1  g045(.A(new_n230), .B(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n226), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(G902), .ZN(new_n235));
  OAI211_X1 g049(.A(new_n216), .B(new_n232), .C1(new_n221), .C2(new_n225), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n234), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  NOR2_X1   g051(.A1(KEYINPUT82), .A2(KEYINPUT25), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(new_n238), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n234), .A2(new_n235), .A3(new_n236), .A4(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(KEYINPUT82), .A2(KEYINPUT25), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n239), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(G234), .ZN(new_n244));
  OAI21_X1  g058(.A(G217), .B1(new_n244), .B2(G902), .ZN(new_n245));
  XNOR2_X1  g059(.A(new_n245), .B(KEYINPUT78), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n243), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n245), .A2(new_n235), .ZN(new_n249));
  XNOR2_X1  g063(.A(new_n249), .B(KEYINPUT84), .ZN(new_n250));
  INV_X1    g064(.A(new_n234), .ZN(new_n251));
  INV_X1    g065(.A(new_n236), .ZN(new_n252));
  OAI21_X1  g066(.A(KEYINPUT83), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  NOR3_X1   g068(.A1(new_n251), .A2(KEYINPUT83), .A3(new_n252), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n250), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n248), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT2), .ZN(new_n258));
  INV_X1    g072(.A(G113), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n258), .A2(new_n259), .A3(KEYINPUT70), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT70), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n261), .B1(KEYINPUT2), .B2(G113), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(KEYINPUT2), .A2(G113), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  OR2_X1    g079(.A1(KEYINPUT71), .A2(G116), .ZN(new_n266));
  NAND2_X1  g080(.A1(KEYINPUT71), .A2(G116), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n266), .A2(G119), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n204), .A2(G116), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n265), .A2(new_n270), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n263), .A2(new_n268), .A3(new_n264), .A4(new_n269), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT66), .ZN(new_n274));
  INV_X1    g088(.A(G137), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n274), .B1(new_n275), .B2(G134), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(G134), .ZN(new_n277));
  INV_X1    g091(.A(G134), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n278), .A2(KEYINPUT66), .A3(G137), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n276), .A2(new_n277), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(G131), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(KEYINPUT67), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT65), .ZN(new_n283));
  INV_X1    g097(.A(G143), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n283), .B1(new_n284), .B2(G146), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n194), .A2(KEYINPUT65), .A3(G143), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n202), .A2(KEYINPUT1), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n284), .A2(G146), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n285), .A2(new_n286), .A3(new_n287), .A4(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n194), .A2(G143), .ZN(new_n290));
  AOI22_X1  g104(.A1(new_n198), .A2(new_n199), .B1(new_n290), .B2(KEYINPUT1), .ZN(new_n291));
  AND2_X1   g105(.A1(new_n290), .A2(new_n288), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n289), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(KEYINPUT11), .B1(new_n278), .B2(G137), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT11), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n295), .A2(new_n275), .A3(G134), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G131), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n275), .A2(G134), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n297), .A2(new_n298), .A3(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT67), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n280), .A2(new_n302), .A3(G131), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n282), .A2(new_n293), .A3(new_n301), .A4(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(KEYINPUT72), .ZN(new_n305));
  AND2_X1   g119(.A1(new_n303), .A2(new_n301), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT72), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n306), .A2(new_n307), .A3(new_n293), .A4(new_n282), .ZN(new_n308));
  AND3_X1   g122(.A1(new_n285), .A2(new_n286), .A3(new_n288), .ZN(new_n309));
  NAND2_X1  g123(.A1(KEYINPUT0), .A2(G128), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  XNOR2_X1  g126(.A(new_n310), .B(KEYINPUT64), .ZN(new_n313));
  NOR2_X1   g127(.A1(KEYINPUT0), .A2(G128), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n314), .B1(new_n290), .B2(new_n288), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  AOI211_X1 g130(.A(G131), .B(new_n299), .C1(new_n294), .C2(new_n296), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n298), .B1(new_n297), .B2(new_n300), .ZN(new_n318));
  OAI211_X1 g132(.A(new_n312), .B(new_n316), .C1(new_n317), .C2(new_n318), .ZN(new_n319));
  NAND4_X1  g133(.A1(new_n305), .A2(new_n308), .A3(KEYINPUT30), .A4(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT69), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n304), .A2(new_n319), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT30), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n321), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  AOI211_X1 g138(.A(KEYINPUT69), .B(KEYINPUT30), .C1(new_n304), .C2(new_n319), .ZN(new_n325));
  OAI211_X1 g139(.A(new_n273), .B(new_n320), .C1(new_n324), .C2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(new_n273), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n305), .A2(new_n308), .A3(new_n327), .A4(new_n319), .ZN(new_n328));
  INV_X1    g142(.A(G237), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n229), .A2(G210), .A3(new_n329), .ZN(new_n330));
  XNOR2_X1  g144(.A(new_n330), .B(KEYINPUT27), .ZN(new_n331));
  XNOR2_X1  g145(.A(KEYINPUT26), .B(G101), .ZN(new_n332));
  XNOR2_X1  g146(.A(new_n331), .B(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n326), .A2(new_n328), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(KEYINPUT31), .ZN(new_n335));
  INV_X1    g149(.A(new_n333), .ZN(new_n336));
  AND2_X1   g150(.A1(new_n304), .A2(new_n319), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT74), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n273), .B1(new_n322), .B2(KEYINPUT74), .ZN(new_n340));
  AOI21_X1  g154(.A(KEYINPUT28), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT28), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n322), .A2(new_n273), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n342), .B1(new_n328), .B2(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n336), .B1(new_n341), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT31), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n326), .A2(new_n346), .A3(new_n328), .A4(new_n333), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n335), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  NOR2_X1   g162(.A1(G472), .A2(G902), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(KEYINPUT75), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT75), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n348), .A2(new_n352), .A3(new_n349), .ZN(new_n353));
  XNOR2_X1  g167(.A(KEYINPUT76), .B(KEYINPUT32), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n351), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  AND2_X1   g169(.A1(new_n348), .A2(new_n349), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n333), .B1(new_n341), .B2(new_n344), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n326), .A2(new_n328), .A3(new_n336), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT29), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  AND2_X1   g175(.A1(new_n308), .A2(new_n319), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n362), .A2(KEYINPUT77), .A3(new_n327), .A4(new_n305), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n308), .A2(new_n319), .ZN(new_n364));
  INV_X1    g178(.A(new_n305), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n273), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT77), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n328), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n363), .A2(new_n366), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(KEYINPUT28), .ZN(new_n370));
  INV_X1    g184(.A(new_n341), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n370), .A2(KEYINPUT29), .A3(new_n371), .A4(new_n333), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n361), .A2(new_n372), .A3(new_n235), .ZN(new_n373));
  AOI22_X1  g187(.A1(new_n356), .A2(KEYINPUT32), .B1(new_n373), .B2(G472), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n257), .B1(new_n355), .B2(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(G210), .B1(G237), .B2(G902), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n376), .B(KEYINPUT94), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(KEYINPUT93), .ZN(new_n378));
  XNOR2_X1  g192(.A(G110), .B(G122), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(G104), .ZN(new_n381));
  OAI21_X1  g195(.A(KEYINPUT3), .B1(new_n381), .B2(G107), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT3), .ZN(new_n383));
  INV_X1    g197(.A(G107), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n383), .A2(new_n384), .A3(G104), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n381), .A2(G107), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n382), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(KEYINPUT86), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT4), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT86), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n382), .A2(new_n385), .A3(new_n390), .A4(new_n386), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n388), .A2(new_n389), .A3(G101), .A4(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n273), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n388), .A2(G101), .A3(new_n391), .ZN(new_n394));
  INV_X1    g208(.A(G101), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n382), .A2(new_n385), .A3(new_n395), .A4(new_n386), .ZN(new_n396));
  AND2_X1   g210(.A1(new_n396), .A2(KEYINPUT4), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n394), .A2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT87), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n394), .A2(KEYINPUT87), .A3(new_n397), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n393), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  AND3_X1   g216(.A1(new_n268), .A2(KEYINPUT5), .A3(new_n269), .ZN(new_n403));
  OAI21_X1  g217(.A(G113), .B1(new_n269), .B2(KEYINPUT5), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(new_n272), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n381), .A2(G107), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n384), .A2(G104), .ZN(new_n408));
  OAI21_X1  g222(.A(G101), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n396), .A2(new_n409), .ZN(new_n410));
  NOR3_X1   g224(.A1(new_n405), .A2(new_n406), .A3(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n380), .B1(new_n402), .B2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n411), .ZN(new_n413));
  AND3_X1   g227(.A1(new_n394), .A2(KEYINPUT87), .A3(new_n397), .ZN(new_n414));
  AOI21_X1  g228(.A(KEYINPUT87), .B1(new_n394), .B2(new_n397), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  OAI211_X1 g230(.A(new_n379), .B(new_n413), .C1(new_n416), .C2(new_n393), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n412), .A2(new_n417), .A3(KEYINPUT6), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT6), .ZN(new_n419));
  OAI211_X1 g233(.A(new_n419), .B(new_n380), .C1(new_n402), .C2(new_n411), .ZN(new_n420));
  AOI22_X1  g234(.A1(new_n309), .A2(new_n311), .B1(new_n313), .B2(new_n315), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n421), .A2(new_n189), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n293), .A2(G125), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(G953), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(G224), .ZN(new_n426));
  XNOR2_X1  g240(.A(new_n424), .B(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n418), .A2(new_n420), .A3(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT91), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n418), .A2(KEYINPUT91), .A3(new_n420), .A4(new_n427), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n424), .B1(KEYINPUT7), .B2(new_n426), .ZN(new_n433));
  XOR2_X1   g247(.A(new_n379), .B(KEYINPUT8), .Z(new_n434));
  INV_X1    g248(.A(new_n410), .ZN(new_n435));
  XOR2_X1   g249(.A(new_n404), .B(KEYINPUT92), .Z(new_n436));
  OAI211_X1 g250(.A(new_n272), .B(new_n435), .C1(new_n436), .C2(new_n403), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n410), .B1(new_n405), .B2(new_n406), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n434), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT7), .ZN(new_n440));
  INV_X1    g254(.A(new_n426), .ZN(new_n441));
  NOR4_X1   g255(.A1(new_n422), .A2(new_n423), .A3(new_n440), .A4(new_n441), .ZN(new_n442));
  NOR3_X1   g256(.A1(new_n433), .A2(new_n439), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(new_n417), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n235), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n378), .B1(new_n432), .B2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n378), .ZN(new_n448));
  AOI211_X1 g262(.A(new_n448), .B(new_n445), .C1(new_n430), .C2(new_n431), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  OAI21_X1  g264(.A(G214), .B1(G237), .B2(G902), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  NOR2_X1   g267(.A1(KEYINPUT89), .A2(KEYINPUT12), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n290), .A2(new_n288), .ZN(new_n455));
  AND2_X1   g269(.A1(KEYINPUT68), .A2(G128), .ZN(new_n456));
  NOR2_X1   g270(.A1(KEYINPUT68), .A2(G128), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT1), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n459), .B1(G143), .B2(new_n194), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n455), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  AND3_X1   g275(.A1(new_n410), .A2(new_n289), .A3(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n285), .A2(new_n286), .A3(new_n288), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n284), .A2(G146), .ZN(new_n464));
  OAI21_X1  g278(.A(G128), .B1(new_n464), .B2(new_n459), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(KEYINPUT88), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT88), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n463), .A2(new_n465), .A3(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n467), .A2(new_n289), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n462), .B1(new_n470), .B2(new_n435), .ZN(new_n471));
  INV_X1    g285(.A(new_n318), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(new_n301), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n454), .B1(new_n471), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n454), .ZN(new_n476));
  AND4_X1   g290(.A1(new_n285), .A2(new_n286), .A3(new_n287), .A4(new_n288), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n477), .B1(new_n466), .B2(KEYINPUT88), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n410), .B1(new_n478), .B2(new_n469), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n473), .B(new_n476), .C1(new_n479), .C2(new_n462), .ZN(new_n480));
  NAND2_X1  g294(.A1(KEYINPUT89), .A2(KEYINPUT12), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n475), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n229), .A2(G227), .ZN(new_n483));
  XOR2_X1   g297(.A(G110), .B(G140), .Z(new_n484));
  XNOR2_X1  g298(.A(new_n483), .B(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n435), .A2(new_n293), .A3(KEYINPUT10), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n470), .A2(new_n435), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT10), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n392), .A2(new_n421), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n493), .B1(new_n414), .B2(new_n415), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n491), .A2(new_n494), .A3(new_n474), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n482), .A2(new_n486), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n492), .B1(new_n400), .B2(new_n401), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n487), .B1(new_n479), .B2(KEYINPUT10), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n473), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n486), .B1(new_n499), .B2(new_n495), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n496), .B1(new_n500), .B2(KEYINPUT90), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT90), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n482), .A2(new_n502), .A3(new_n486), .A4(new_n495), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(G469), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n504), .A2(new_n505), .A3(new_n235), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n499), .A2(new_n495), .A3(new_n486), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n486), .B1(new_n482), .B2(new_n495), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(G469), .B1(new_n510), .B2(G902), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n506), .A2(new_n511), .ZN(new_n512));
  XNOR2_X1  g326(.A(KEYINPUT9), .B(G234), .ZN(new_n513));
  OAI21_X1  g327(.A(G221), .B1(new_n513), .B2(G902), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n514), .B(KEYINPUT85), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n512), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g331(.A1(G475), .A2(G902), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n518), .B(KEYINPUT99), .ZN(new_n519));
  XNOR2_X1  g333(.A(G113), .B(G122), .ZN(new_n520));
  XNOR2_X1  g334(.A(KEYINPUT98), .B(G104), .ZN(new_n521));
  XOR2_X1   g335(.A(new_n520), .B(new_n521), .Z(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  OR2_X1    g337(.A1(KEYINPUT73), .A2(G953), .ZN(new_n524));
  NAND2_X1  g338(.A1(KEYINPUT73), .A2(G953), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n524), .A2(G214), .A3(new_n329), .A4(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(new_n284), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n229), .A2(G143), .A3(G214), .A4(new_n329), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(G131), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT96), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n529), .A2(KEYINPUT96), .A3(G131), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n527), .A2(new_n528), .A3(new_n298), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT97), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n532), .A2(KEYINPUT97), .A3(new_n533), .A4(new_n534), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n195), .A2(KEYINPUT19), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n195), .B(KEYINPUT95), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n539), .B1(new_n540), .B2(KEYINPUT19), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n193), .B1(new_n541), .B2(new_n194), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n537), .A2(new_n538), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n540), .A2(G146), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n544), .B1(G146), .B2(new_n195), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n529), .A2(KEYINPUT18), .A3(G131), .ZN(new_n546));
  NAND2_X1  g360(.A1(KEYINPUT18), .A2(G131), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n527), .A2(new_n528), .A3(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n545), .A2(new_n546), .A3(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n523), .B1(new_n543), .B2(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(KEYINPUT96), .B1(new_n529), .B2(G131), .ZN(new_n551));
  AOI211_X1 g365(.A(new_n531), .B(new_n298), .C1(new_n527), .C2(new_n528), .ZN(new_n552));
  OAI21_X1  g366(.A(KEYINPUT17), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n218), .B(new_n553), .C1(new_n535), .C2(KEYINPUT17), .ZN(new_n554));
  AND3_X1   g368(.A1(new_n554), .A2(new_n523), .A3(new_n549), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n519), .B1(new_n550), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(KEYINPUT20), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT20), .ZN(new_n558));
  OAI211_X1 g372(.A(new_n558), .B(new_n519), .C1(new_n550), .C2(new_n555), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n523), .B1(new_n554), .B2(new_n549), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n235), .B1(new_n555), .B2(new_n560), .ZN(new_n561));
  XNOR2_X1  g375(.A(KEYINPUT100), .B(G475), .ZN(new_n562));
  AOI22_X1  g376(.A1(new_n557), .A2(new_n559), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  AND2_X1   g377(.A1(new_n425), .A2(G952), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n564), .B1(new_n244), .B2(new_n329), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  AOI211_X1 g380(.A(new_n235), .B(new_n229), .C1(G234), .C2(G237), .ZN(new_n567));
  XNOR2_X1  g381(.A(KEYINPUT21), .B(G898), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n266), .A2(G122), .A3(new_n267), .ZN(new_n571));
  INV_X1    g385(.A(G116), .ZN(new_n572));
  OR2_X1    g386(.A1(new_n572), .A2(G122), .ZN(new_n573));
  AND3_X1   g387(.A1(new_n571), .A2(new_n384), .A3(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n198), .A2(G143), .A3(new_n199), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n575), .B1(new_n202), .B2(G143), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(G134), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n575), .B(new_n278), .C1(new_n202), .C2(G143), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n574), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT14), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n571), .A2(new_n580), .A3(new_n573), .ZN(new_n581));
  OAI211_X1 g395(.A(new_n581), .B(G107), .C1(new_n580), .C2(new_n571), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT13), .ZN(new_n584));
  OAI221_X1 g398(.A(new_n575), .B1(new_n584), .B2(new_n278), .C1(new_n202), .C2(G143), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n384), .B1(new_n571), .B2(new_n573), .ZN(new_n586));
  AOI21_X1  g400(.A(KEYINPUT13), .B1(new_n458), .B2(G143), .ZN(new_n587));
  OAI221_X1 g401(.A(new_n585), .B1(new_n574), .B2(new_n586), .C1(new_n577), .C2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n583), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(G217), .ZN(new_n590));
  NOR3_X1   g404(.A1(new_n513), .A2(new_n590), .A3(G953), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n583), .A2(new_n588), .A3(new_n591), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n593), .A2(KEYINPUT101), .A3(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT101), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n589), .A2(new_n596), .A3(new_n592), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n595), .A2(new_n235), .A3(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(G478), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n599), .A2(KEYINPUT15), .ZN(new_n600));
  XOR2_X1   g414(.A(new_n598), .B(new_n600), .Z(new_n601));
  NAND3_X1  g415(.A1(new_n563), .A2(new_n570), .A3(new_n601), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n517), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n375), .A2(new_n453), .A3(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(G101), .ZN(G3));
  INV_X1    g419(.A(new_n377), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n606), .B1(new_n432), .B2(new_n446), .ZN(new_n607));
  AOI211_X1 g421(.A(new_n377), .B(new_n445), .C1(new_n430), .C2(new_n431), .ZN(new_n608));
  OR2_X1    g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n598), .A2(new_n599), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(KEYINPUT102), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT102), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n598), .A2(new_n612), .A3(new_n599), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT33), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n595), .A2(new_n614), .A3(new_n597), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n593), .A2(KEYINPUT33), .A3(new_n594), .ZN(new_n616));
  AND2_X1   g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n599), .A2(G902), .ZN(new_n618));
  AOI22_X1  g432(.A1(new_n611), .A2(new_n613), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NOR3_X1   g433(.A1(new_n563), .A2(new_n569), .A3(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT103), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n609), .A2(new_n620), .A3(new_n621), .A4(new_n451), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n451), .B1(new_n607), .B2(new_n608), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n557), .A2(new_n559), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n561), .A2(new_n562), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n619), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n626), .A2(new_n627), .A3(new_n570), .ZN(new_n628));
  OAI21_X1  g442(.A(KEYINPUT103), .B1(new_n623), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n622), .A2(new_n629), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n515), .B1(new_n506), .B2(new_n511), .ZN(new_n631));
  INV_X1    g445(.A(new_n242), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n632), .B1(new_n237), .B2(new_n238), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n246), .B1(new_n633), .B2(new_n241), .ZN(new_n634));
  INV_X1    g448(.A(new_n255), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(new_n253), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n634), .B1(new_n250), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n631), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n348), .A2(new_n235), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(G472), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n351), .A2(new_n640), .A3(new_n353), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n638), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n630), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT34), .B(G104), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G6));
  INV_X1    g459(.A(new_n623), .ZN(new_n646));
  INV_X1    g460(.A(new_n601), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n563), .A2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n646), .A2(new_n570), .A3(new_n649), .ZN(new_n650));
  NOR3_X1   g464(.A1(new_n650), .A2(new_n641), .A3(new_n638), .ZN(new_n651));
  XNOR2_X1  g465(.A(KEYINPUT35), .B(G107), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G9));
  INV_X1    g467(.A(KEYINPUT105), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n233), .A2(KEYINPUT36), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n226), .A2(new_n656), .ZN(new_n657));
  OAI211_X1 g471(.A(new_n216), .B(new_n655), .C1(new_n221), .C2(new_n225), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n657), .A2(new_n250), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(KEYINPUT104), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n248), .A2(new_n654), .A3(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT104), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n659), .B(new_n662), .ZN(new_n663));
  OAI21_X1  g477(.A(KEYINPUT105), .B1(new_n634), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n641), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n666), .A2(new_n453), .A3(new_n603), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT37), .B(G110), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G12));
  AOI21_X1  g483(.A(new_n665), .B1(new_n355), .B2(new_n374), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n623), .A2(new_n517), .ZN(new_n671));
  INV_X1    g485(.A(G900), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n566), .B1(new_n567), .B2(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n648), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n670), .A2(new_n671), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G128), .ZN(G30));
  XOR2_X1   g490(.A(new_n450), .B(KEYINPUT38), .Z(new_n677));
  NOR2_X1   g491(.A1(new_n601), .A2(new_n452), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n626), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n248), .A2(new_n660), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  XOR2_X1   g495(.A(new_n673), .B(KEYINPUT39), .Z(new_n682));
  NAND2_X1  g496(.A1(new_n631), .A2(new_n682), .ZN(new_n683));
  OR2_X1    g497(.A1(new_n683), .A2(KEYINPUT40), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n348), .A2(KEYINPUT32), .A3(new_n349), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n235), .B1(new_n369), .B2(new_n333), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n336), .B1(new_n326), .B2(new_n328), .ZN(new_n687));
  OAI21_X1  g501(.A(G472), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  AND2_X1   g502(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  AOI22_X1  g503(.A1(new_n683), .A2(KEYINPUT40), .B1(new_n355), .B2(new_n689), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n677), .A2(new_n681), .A3(new_n684), .A4(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G143), .ZN(G45));
  NOR3_X1   g506(.A1(new_n563), .A2(new_n619), .A3(new_n673), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n670), .A2(new_n671), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G146), .ZN(G48));
  AND2_X1   g509(.A1(new_n622), .A2(new_n629), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n355), .A2(new_n374), .ZN(new_n697));
  AND4_X1   g511(.A1(new_n502), .A2(new_n482), .A3(new_n486), .A4(new_n495), .ZN(new_n698));
  NOR3_X1   g512(.A1(new_n497), .A2(new_n498), .A3(new_n473), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n474), .B1(new_n491), .B2(new_n494), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n485), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(new_n502), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n698), .B1(new_n702), .B2(new_n496), .ZN(new_n703));
  OAI21_X1  g517(.A(G469), .B1(new_n703), .B2(G902), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n704), .A2(new_n516), .A3(new_n506), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(KEYINPUT106), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT106), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n704), .A2(new_n707), .A3(new_n516), .A4(new_n506), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n697), .A2(new_n637), .A3(new_n706), .A4(new_n708), .ZN(new_n709));
  OAI21_X1  g523(.A(KEYINPUT107), .B1(new_n696), .B2(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(new_n709), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT107), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n711), .A2(new_n712), .A3(new_n630), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(KEYINPUT41), .B(G113), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n714), .B(new_n715), .ZN(G15));
  NOR2_X1   g530(.A1(new_n709), .A2(new_n650), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(new_n572), .ZN(G18));
  INV_X1    g532(.A(new_n602), .ZN(new_n719));
  INV_X1    g533(.A(new_n665), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n697), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n646), .A2(new_n708), .A3(new_n706), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(new_n204), .ZN(G21));
  NAND2_X1  g538(.A1(new_n335), .A2(new_n347), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n333), .B1(new_n370), .B2(new_n371), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n349), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  AND3_X1   g541(.A1(new_n637), .A2(new_n640), .A3(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n728), .A2(new_n706), .A3(new_n708), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n609), .A2(new_n570), .A3(new_n626), .A4(new_n678), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  XOR2_X1   g545(.A(new_n731), .B(G122), .Z(G24));
  INV_X1    g546(.A(new_n673), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n626), .A2(new_n627), .A3(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n640), .A2(new_n680), .A3(new_n727), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n736), .A2(new_n646), .A3(new_n708), .A4(new_n706), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G125), .ZN(G27));
  AOI211_X1 g552(.A(G469), .B(G902), .C1(new_n501), .C2(new_n503), .ZN(new_n739));
  AND2_X1   g553(.A1(new_n482), .A2(new_n495), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n507), .B1(new_n740), .B2(new_n486), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n505), .B1(new_n741), .B2(new_n235), .ZN(new_n742));
  OAI21_X1  g556(.A(KEYINPUT108), .B1(new_n739), .B2(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT108), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n506), .A2(new_n744), .A3(new_n511), .ZN(new_n745));
  AND3_X1   g559(.A1(new_n743), .A2(new_n516), .A3(new_n745), .ZN(new_n746));
  NOR3_X1   g560(.A1(new_n447), .A2(new_n449), .A3(new_n452), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n375), .A2(new_n746), .A3(new_n693), .A4(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT42), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT109), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n746), .A2(new_n747), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n373), .A2(G472), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT32), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n350), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n753), .A2(new_n755), .A3(new_n685), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n693), .A2(new_n756), .A3(KEYINPUT42), .A4(new_n637), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n751), .B1(new_n752), .B2(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n743), .A2(new_n516), .A3(new_n745), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n432), .A2(new_n446), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(new_n448), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n432), .A2(new_n378), .A3(new_n446), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n761), .A2(new_n451), .A3(new_n762), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n759), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n756), .A2(new_n637), .ZN(new_n765));
  INV_X1    g579(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n734), .A2(new_n749), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n764), .A2(new_n766), .A3(KEYINPUT109), .A4(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n750), .A2(new_n758), .A3(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G131), .ZN(G33));
  NAND3_X1  g584(.A1(new_n764), .A2(new_n375), .A3(new_n674), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G134), .ZN(G36));
  XNOR2_X1  g586(.A(KEYINPUT111), .B(KEYINPUT43), .ZN(new_n773));
  NOR3_X1   g587(.A1(new_n626), .A2(new_n619), .A3(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT111), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(KEYINPUT43), .ZN(new_n776));
  INV_X1    g590(.A(new_n776), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n777), .B1(new_n627), .B2(new_n563), .ZN(new_n778));
  OAI211_X1 g592(.A(new_n641), .B(new_n680), .C1(new_n774), .C2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT44), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n763), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  OR2_X1    g595(.A1(new_n774), .A2(new_n778), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n782), .A2(KEYINPUT44), .A3(new_n641), .A4(new_n680), .ZN(new_n783));
  INV_X1    g597(.A(new_n682), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT110), .ZN(new_n785));
  OAI211_X1 g599(.A(KEYINPUT45), .B(new_n507), .C1(new_n740), .C2(new_n486), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT45), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n787), .B1(new_n508), .B2(new_n509), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n786), .A2(new_n788), .A3(G469), .ZN(new_n789));
  NAND2_X1  g603(.A1(G469), .A2(G902), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT46), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n785), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n789), .A2(KEYINPUT110), .A3(KEYINPUT46), .A4(new_n790), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n739), .B1(new_n791), .B2(new_n792), .ZN(new_n796));
  AOI211_X1 g610(.A(new_n515), .B(new_n784), .C1(new_n795), .C2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n781), .A2(new_n783), .A3(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G137), .ZN(G39));
  AOI21_X1  g613(.A(new_n515), .B1(new_n795), .B2(new_n796), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT112), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(KEYINPUT47), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  NOR4_X1   g617(.A1(new_n697), .A2(new_n763), .A3(new_n734), .A4(new_n637), .ZN(new_n804));
  XNOR2_X1  g618(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n803), .B(new_n804), .C1(new_n800), .C2(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(G140), .ZN(G42));
  NAND2_X1  g621(.A1(new_n355), .A2(new_n689), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n704), .A2(new_n506), .ZN(new_n809));
  XOR2_X1   g623(.A(new_n809), .B(KEYINPUT113), .Z(new_n810));
  INV_X1    g624(.A(new_n810), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n808), .B1(new_n811), .B2(KEYINPUT49), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n637), .A2(new_n451), .A3(new_n516), .ZN(new_n813));
  NOR4_X1   g627(.A1(new_n677), .A2(new_n626), .A3(new_n619), .A4(new_n813), .ZN(new_n814));
  OAI211_X1 g628(.A(new_n812), .B(new_n814), .C1(KEYINPUT49), .C2(new_n811), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT54), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n563), .A2(new_n601), .A3(new_n733), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n763), .A2(new_n517), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(new_n670), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n764), .A2(new_n736), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n771), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n626), .A2(new_n627), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n569), .B1(new_n822), .B2(new_n648), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n642), .A2(new_n453), .A3(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n824), .A2(new_n604), .A3(new_n667), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n821), .A2(new_n825), .ZN(new_n826));
  OAI22_X1  g640(.A1(new_n709), .A2(new_n650), .B1(new_n729), .B2(new_n730), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n827), .A2(new_n723), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n714), .A2(new_n826), .A3(new_n769), .A4(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT53), .ZN(new_n830));
  OAI211_X1 g644(.A(new_n670), .B(new_n671), .C1(new_n674), .C2(new_n693), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n607), .A2(new_n608), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n832), .A2(new_n679), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n743), .A2(new_n745), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n680), .A2(new_n515), .A3(new_n673), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n833), .A2(new_n834), .A3(new_n808), .A4(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n831), .A2(new_n737), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(KEYINPUT52), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT52), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n831), .A2(new_n839), .A3(new_n737), .A4(new_n836), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n829), .A2(new_n830), .A3(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT115), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n842), .B(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n841), .B1(new_n829), .B2(KEYINPUT114), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n845), .B1(KEYINPUT114), .B2(new_n829), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(new_n830), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n816), .B1(new_n844), .B2(new_n847), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n696), .A2(KEYINPUT107), .A3(new_n709), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n712), .B1(new_n711), .B2(new_n630), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n828), .B(new_n769), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(KEYINPUT116), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT116), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n714), .A2(new_n853), .A3(new_n769), .A4(new_n828), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n824), .A2(new_n604), .A3(new_n667), .ZN(new_n855));
  AOI22_X1  g669(.A1(new_n818), .A2(new_n670), .B1(new_n764), .B2(new_n736), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n855), .A2(KEYINPUT53), .A3(new_n771), .A4(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n841), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n852), .A2(new_n854), .A3(new_n858), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n830), .B1(new_n829), .B2(new_n841), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n859), .A2(new_n860), .A3(new_n816), .ZN(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n677), .A2(new_n451), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n706), .A2(new_n708), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n782), .A2(new_n566), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n863), .A2(new_n864), .A3(new_n728), .A4(new_n865), .ZN(new_n866));
  XOR2_X1   g680(.A(new_n866), .B(KEYINPUT50), .Z(new_n867));
  OAI21_X1  g681(.A(new_n803), .B1(new_n800), .B2(new_n805), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n868), .B1(new_n516), .B2(new_n811), .ZN(new_n869));
  AND2_X1   g683(.A1(new_n865), .A2(new_n728), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n869), .A2(new_n747), .A3(new_n870), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n864), .A2(new_n566), .A3(new_n747), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n872), .A2(new_n355), .A3(new_n637), .A4(new_n689), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n873), .A2(new_n626), .A3(new_n627), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n872), .A2(new_n782), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n875), .A2(new_n735), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n867), .A2(new_n871), .A3(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT51), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n867), .A2(KEYINPUT51), .A3(new_n871), .A4(new_n877), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n875), .A2(new_n765), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(KEYINPUT48), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n870), .A2(new_n646), .A3(new_n864), .ZN(new_n884));
  OAI211_X1 g698(.A(new_n884), .B(new_n564), .C1(new_n822), .C2(new_n873), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n880), .A2(new_n881), .A3(new_n886), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n848), .A2(new_n862), .A3(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(G952), .A2(G953), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n815), .B1(new_n888), .B2(new_n889), .ZN(G75));
  NOR2_X1   g704(.A1(new_n229), .A2(G952), .ZN(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n235), .B1(new_n859), .B2(new_n860), .ZN(new_n893));
  AOI21_X1  g707(.A(KEYINPUT56), .B1(new_n893), .B2(new_n377), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n418), .A2(new_n420), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(new_n427), .ZN(new_n896));
  XOR2_X1   g710(.A(KEYINPUT117), .B(KEYINPUT55), .Z(new_n897));
  XNOR2_X1  g711(.A(new_n896), .B(new_n897), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n892), .B1(new_n894), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n894), .A2(new_n898), .ZN(new_n900));
  OR2_X1    g714(.A1(new_n900), .A2(KEYINPUT118), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(KEYINPUT118), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n899), .B1(new_n901), .B2(new_n902), .ZN(G51));
  AOI211_X1 g717(.A(new_n235), .B(new_n789), .C1(new_n859), .C2(new_n860), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n859), .A2(new_n860), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(KEYINPUT54), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(new_n861), .ZN(new_n907));
  XOR2_X1   g721(.A(new_n790), .B(KEYINPUT57), .Z(new_n908));
  AOI21_X1  g722(.A(new_n703), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n904), .B1(new_n909), .B2(KEYINPUT119), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT119), .ZN(new_n911));
  INV_X1    g725(.A(new_n908), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n912), .B1(new_n906), .B2(new_n861), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n911), .B1(new_n913), .B2(new_n703), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n891), .B1(new_n910), .B2(new_n914), .ZN(G54));
  AND3_X1   g729(.A1(new_n893), .A2(KEYINPUT58), .A3(G475), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n550), .A2(new_n555), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  OAI21_X1  g732(.A(KEYINPUT120), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n891), .B1(new_n916), .B2(new_n918), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NOR3_X1   g735(.A1(new_n916), .A2(KEYINPUT120), .A3(new_n918), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n921), .A2(new_n922), .ZN(G60));
  NAND2_X1  g737(.A1(G478), .A2(G902), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT59), .Z(new_n925));
  INV_X1    g739(.A(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n907), .A2(new_n617), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(new_n892), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n926), .B1(new_n848), .B2(new_n862), .ZN(new_n929));
  INV_X1    g743(.A(new_n617), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n928), .B1(new_n929), .B2(new_n930), .ZN(G63));
  NAND2_X1  g745(.A1(G217), .A2(G902), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT60), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n933), .B1(new_n859), .B2(new_n860), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n934), .A2(new_n658), .A3(new_n657), .ZN(new_n935));
  OAI211_X1 g749(.A(new_n935), .B(new_n892), .C1(new_n636), .C2(new_n934), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT61), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n936), .B(new_n937), .ZN(G66));
  INV_X1    g752(.A(new_n568), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n425), .B1(new_n939), .B2(G224), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n714), .A2(new_n828), .A3(new_n855), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n940), .B1(new_n941), .B2(new_n229), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n895), .B1(G898), .B2(new_n229), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n942), .B(new_n943), .Z(G69));
  AND2_X1   g758(.A1(new_n831), .A2(new_n737), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(new_n691), .ZN(new_n946));
  OR2_X1    g760(.A1(new_n946), .A2(KEYINPUT62), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT121), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n947), .B(new_n948), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n822), .A2(new_n648), .ZN(new_n950));
  NOR3_X1   g764(.A1(new_n950), .A2(new_n683), .A3(new_n763), .ZN(new_n951));
  AND2_X1   g765(.A1(new_n951), .A2(new_n375), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT122), .ZN(new_n953));
  AND3_X1   g767(.A1(new_n953), .A2(new_n798), .A3(new_n806), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n946), .A2(KEYINPUT62), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n229), .B1(new_n949), .B2(new_n956), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n320), .B1(new_n324), .B2(new_n325), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(new_n541), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT124), .ZN(new_n961));
  AND3_X1   g775(.A1(new_n769), .A2(new_n806), .A3(new_n798), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n831), .A2(new_n771), .A3(new_n737), .ZN(new_n963));
  NOR3_X1   g777(.A1(new_n765), .A2(new_n832), .A3(new_n679), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n963), .B1(new_n797), .B2(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n961), .B1(new_n962), .B2(new_n965), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n769), .A2(new_n806), .A3(new_n798), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n797), .A2(new_n964), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n945), .A2(new_n968), .A3(new_n771), .ZN(new_n969));
  NOR3_X1   g783(.A1(new_n967), .A2(new_n969), .A3(KEYINPUT124), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n229), .B1(new_n966), .B2(new_n970), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n229), .A2(G900), .ZN(new_n972));
  INV_X1    g786(.A(new_n972), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n971), .A2(KEYINPUT125), .A3(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT125), .ZN(new_n975));
  INV_X1    g789(.A(new_n229), .ZN(new_n976));
  AND2_X1   g790(.A1(new_n769), .A2(new_n798), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n977), .A2(new_n961), .A3(new_n806), .A4(new_n965), .ZN(new_n978));
  OAI21_X1  g792(.A(KEYINPUT124), .B1(new_n967), .B2(new_n969), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n976), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n975), .B1(new_n980), .B2(new_n972), .ZN(new_n981));
  INV_X1    g795(.A(new_n959), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n974), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n960), .A2(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(KEYINPUT123), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n229), .B1(G227), .B2(G900), .ZN(new_n987));
  INV_X1    g801(.A(new_n987), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n984), .A2(new_n986), .A3(new_n988), .ZN(new_n989));
  OAI211_X1 g803(.A(new_n960), .B(new_n983), .C1(new_n985), .C2(new_n987), .ZN(new_n990));
  AND2_X1   g804(.A1(new_n989), .A2(new_n990), .ZN(G72));
  NAND2_X1  g805(.A1(G472), .A2(G902), .ZN(new_n992));
  XOR2_X1   g806(.A(new_n992), .B(KEYINPUT63), .Z(new_n993));
  XNOR2_X1  g807(.A(new_n947), .B(KEYINPUT121), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n994), .A2(new_n955), .A3(new_n954), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n993), .B1(new_n995), .B2(new_n941), .ZN(new_n996));
  AND2_X1   g810(.A1(new_n996), .A2(new_n687), .ZN(new_n997));
  INV_X1    g811(.A(new_n687), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n998), .A2(new_n358), .A3(new_n993), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n999), .B(KEYINPUT127), .Z(new_n1000));
  AOI21_X1  g814(.A(new_n1000), .B1(new_n844), .B2(new_n847), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n978), .A2(new_n979), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n993), .B1(new_n1002), .B2(new_n941), .ZN(new_n1003));
  XOR2_X1   g817(.A(new_n358), .B(KEYINPUT126), .Z(new_n1004));
  AND2_X1   g818(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NOR4_X1   g819(.A1(new_n997), .A2(new_n891), .A3(new_n1001), .A4(new_n1005), .ZN(G57));
endmodule


