//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 1 0 0 0 0 0 0 0 1 1 1 0 0 0 0 0 1 1 1 1 0 1 0 1 1 0 1 0 0 1 0 0 0 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 1 0 0 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:24 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1250, new_n1251, new_n1252, new_n1253, new_n1255,
    new_n1256, new_n1257, new_n1258, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1319, new_n1320, new_n1321, new_n1322;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  AND2_X1   g0007(.A1(KEYINPUT64), .A2(G68), .ZN(new_n208));
  NOR2_X1   g0008(.A1(KEYINPUT64), .A2(G68), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  AND2_X1   g0010(.A1(new_n210), .A2(G238), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G87), .A2(G250), .ZN(new_n215));
  NAND4_X1  g0015(.A1(new_n212), .A2(new_n213), .A3(new_n214), .A4(new_n215), .ZN(new_n216));
  OAI21_X1  g0016(.A(new_n207), .B1(new_n211), .B2(new_n216), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT1), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n207), .A2(G13), .ZN(new_n219));
  OAI211_X1 g0019(.A(new_n219), .B(G250), .C1(G257), .C2(G264), .ZN(new_n220));
  INV_X1    g0020(.A(KEYINPUT0), .ZN(new_n221));
  NOR2_X1   g0021(.A1(G58), .A2(G68), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n223), .A2(G50), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(G20), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  AOI22_X1  g0028(.A1(new_n220), .A2(new_n221), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n229), .B1(new_n221), .B2(new_n220), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n218), .A2(new_n230), .ZN(G361));
  XOR2_X1   g0031(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n232));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G226), .B(G232), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G250), .B(G257), .Z(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n236), .B(new_n239), .Z(G358));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G58), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(KEYINPUT66), .B(KEYINPUT67), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G87), .B(G116), .Z(new_n246));
  XNOR2_X1  g0046(.A(G97), .B(G107), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(KEYINPUT3), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT3), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G33), .ZN(new_n253));
  INV_X1    g0053(.A(G1698), .ZN(new_n254));
  NAND4_X1  g0054(.A1(new_n251), .A2(new_n253), .A3(G226), .A4(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(KEYINPUT76), .ZN(new_n256));
  XNOR2_X1  g0056(.A(KEYINPUT3), .B(G33), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT76), .ZN(new_n258));
  NAND4_X1  g0058(.A1(new_n257), .A2(new_n258), .A3(G226), .A4(new_n254), .ZN(new_n259));
  NAND2_X1  g0059(.A1(G33), .A2(G97), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n257), .A2(G232), .A3(G1698), .ZN(new_n261));
  NAND4_X1  g0061(.A1(new_n256), .A2(new_n259), .A3(new_n260), .A4(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n226), .B1(G33), .B2(G41), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G1), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n265), .B1(G41), .B2(G45), .ZN(new_n266));
  INV_X1    g0066(.A(G274), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(G33), .A2(G41), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n269), .A2(G1), .A3(G13), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT68), .ZN(new_n271));
  AND3_X1   g0071(.A1(new_n270), .A2(new_n271), .A3(new_n266), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n271), .B1(new_n270), .B2(new_n266), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n268), .B1(new_n274), .B2(G238), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n264), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(KEYINPUT13), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT13), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n264), .A2(new_n275), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G200), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n250), .A2(G20), .ZN(new_n282));
  NOR2_X1   g0082(.A1(G20), .A2(G33), .ZN(new_n283));
  AOI22_X1  g0083(.A1(new_n282), .A2(G77), .B1(new_n283), .B2(G50), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n284), .B1(new_n227), .B2(new_n210), .ZN(new_n285));
  NAND3_X1  g0085(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(new_n226), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  XOR2_X1   g0088(.A(KEYINPUT77), .B(KEYINPUT78), .Z(new_n289));
  XNOR2_X1  g0089(.A(new_n289), .B(KEYINPUT11), .ZN(new_n290));
  OR2_X1    g0090(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n265), .A2(G20), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n265), .A2(G13), .A3(G20), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  OAI21_X1  g0094(.A(KEYINPUT72), .B1(new_n294), .B2(new_n287), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  NOR3_X1   g0096(.A1(new_n294), .A2(new_n287), .A3(KEYINPUT72), .ZN(new_n297));
  OAI211_X1 g0097(.A(G68), .B(new_n292), .C1(new_n296), .C2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n288), .A2(new_n290), .ZN(new_n299));
  XNOR2_X1  g0099(.A(KEYINPUT64), .B(G68), .ZN(new_n300));
  AND3_X1   g0100(.A1(new_n300), .A2(new_n294), .A3(KEYINPUT12), .ZN(new_n301));
  AOI21_X1  g0101(.A(KEYINPUT12), .B1(new_n294), .B2(new_n203), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n291), .A2(new_n298), .A3(new_n299), .A4(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n277), .A2(G190), .A3(new_n279), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n281), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n279), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n278), .B1(new_n264), .B2(new_n275), .ZN(new_n310));
  OAI21_X1  g0110(.A(G169), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(KEYINPUT14), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT14), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n280), .A2(new_n313), .A3(G169), .ZN(new_n314));
  INV_X1    g0114(.A(G179), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n312), .B(new_n314), .C1(new_n280), .C2(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n308), .B1(new_n316), .B2(new_n304), .ZN(new_n317));
  NOR2_X1   g0117(.A1(KEYINPUT75), .A2(KEYINPUT10), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n252), .A2(G33), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n250), .A2(KEYINPUT3), .ZN(new_n320));
  OAI21_X1  g0120(.A(G77), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n251), .A2(new_n253), .A3(G222), .A4(new_n254), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n251), .A2(new_n253), .A3(G223), .A4(G1698), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n321), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(new_n263), .ZN(new_n325));
  INV_X1    g0125(.A(new_n268), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n270), .A2(new_n266), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(KEYINPUT68), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n270), .A2(new_n271), .A3(new_n266), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n328), .A2(G226), .A3(new_n329), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n325), .A2(new_n326), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(G200), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(KEYINPUT74), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n325), .A2(G190), .A3(new_n330), .A4(new_n326), .ZN(new_n334));
  NAND2_X1  g0134(.A1(KEYINPUT75), .A2(KEYINPUT10), .ZN(new_n335));
  AND2_X1   g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT74), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n331), .A2(new_n337), .A3(G200), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n333), .A2(new_n336), .A3(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT69), .ZN(new_n340));
  NOR3_X1   g0140(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n340), .B1(new_n341), .B2(new_n227), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n204), .A2(KEYINPUT69), .A3(G20), .ZN(new_n343));
  OR2_X1    g0143(.A1(KEYINPUT8), .A2(G58), .ZN(new_n344));
  NAND2_X1  g0144(.A1(KEYINPUT8), .A2(G58), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n282), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n283), .A2(G150), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n342), .A2(new_n343), .A3(new_n346), .A4(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(new_n287), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT9), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(KEYINPUT73), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT70), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n352), .B1(new_n294), .B2(new_n287), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n293), .A2(KEYINPUT70), .A3(new_n226), .A4(new_n286), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n353), .A2(G50), .A3(new_n292), .A4(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n294), .A2(new_n201), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n349), .A2(new_n351), .A3(new_n355), .A4(new_n356), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n350), .A2(KEYINPUT73), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n348), .A2(new_n287), .B1(new_n201), .B2(new_n294), .ZN(new_n360));
  INV_X1    g0160(.A(new_n358), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n360), .A2(new_n351), .A3(new_n355), .A4(new_n361), .ZN(new_n362));
  AND2_X1   g0162(.A1(new_n359), .A2(new_n362), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n318), .B1(new_n339), .B2(new_n363), .ZN(new_n364));
  AND3_X1   g0164(.A1(new_n338), .A2(new_n335), .A3(new_n334), .ZN(new_n365));
  INV_X1    g0165(.A(new_n318), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n359), .A2(new_n362), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n365), .A2(new_n366), .A3(new_n367), .A4(new_n333), .ZN(new_n368));
  INV_X1    g0168(.A(G169), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n331), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n360), .A2(new_n355), .ZN(new_n371));
  OAI211_X1 g0171(.A(new_n370), .B(new_n371), .C1(G179), .C2(new_n331), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n364), .A2(new_n368), .A3(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n344), .A2(new_n283), .A3(new_n345), .ZN(new_n374));
  INV_X1    g0174(.A(G77), .ZN(new_n375));
  XNOR2_X1  g0175(.A(KEYINPUT15), .B(G87), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n227), .A2(G33), .ZN(new_n377));
  OAI221_X1 g0177(.A(new_n374), .B1(new_n227), .B2(new_n375), .C1(new_n376), .C2(new_n377), .ZN(new_n378));
  AOI22_X1  g0178(.A1(new_n378), .A2(new_n287), .B1(new_n375), .B2(new_n294), .ZN(new_n379));
  OAI211_X1 g0179(.A(G77), .B(new_n292), .C1(new_n296), .C2(new_n297), .ZN(new_n380));
  AND2_X1   g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g0181(.A(G107), .B1(new_n319), .B2(new_n320), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n251), .A2(new_n253), .A3(G232), .A4(new_n254), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n251), .A2(new_n253), .A3(G238), .A4(G1698), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n382), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(KEYINPUT71), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT71), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n382), .A2(new_n383), .A3(new_n384), .A4(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n386), .A2(new_n263), .A3(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n268), .B1(new_n274), .B2(G244), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n389), .A2(G190), .A3(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n328), .A2(G244), .A3(new_n329), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n326), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n270), .B1(new_n385), .B2(KEYINPUT71), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n393), .B1(new_n388), .B2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(G200), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n381), .B(new_n391), .C1(new_n395), .C2(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n389), .A2(new_n315), .A3(new_n390), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n379), .A2(new_n380), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n398), .B(new_n399), .C1(new_n395), .C2(G169), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n397), .A2(new_n400), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n373), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n317), .A2(new_n402), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n251), .A2(new_n253), .A3(G226), .A4(G1698), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n251), .A2(new_n253), .A3(G223), .A4(new_n254), .ZN(new_n405));
  NAND2_X1  g0205(.A1(G33), .A2(G87), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(new_n263), .ZN(new_n408));
  INV_X1    g0208(.A(new_n327), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n268), .B1(new_n409), .B2(G232), .ZN(new_n410));
  INV_X1    g0210(.A(G190), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n408), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(KEYINPUT80), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT80), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n408), .A2(new_n410), .A3(new_n414), .A4(new_n411), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n408), .A2(new_n410), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(new_n396), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n413), .A2(new_n415), .A3(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT16), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n283), .A2(G159), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n222), .B1(new_n210), .B2(G58), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n420), .B1(new_n421), .B2(new_n227), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT7), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n423), .B1(new_n257), .B2(G20), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n251), .A2(new_n253), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n425), .A2(KEYINPUT7), .A3(new_n227), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n300), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n419), .B1(new_n422), .B2(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(KEYINPUT7), .B1(new_n425), .B2(new_n227), .ZN(new_n429));
  AOI211_X1 g0229(.A(new_n423), .B(G20), .C1(new_n251), .C2(new_n253), .ZN(new_n430));
  OAI21_X1  g0230(.A(G68), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n223), .B1(new_n300), .B2(new_n202), .ZN(new_n432));
  AOI22_X1  g0232(.A1(new_n432), .A2(G20), .B1(G159), .B2(new_n283), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n431), .A2(new_n433), .A3(KEYINPUT16), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n428), .A2(new_n434), .A3(new_n287), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n344), .A2(new_n345), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n353), .A2(new_n292), .A3(new_n437), .A4(new_n354), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n436), .A2(new_n294), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n418), .A2(new_n435), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(KEYINPUT17), .ZN(new_n443));
  INV_X1    g0243(.A(new_n287), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n203), .B1(new_n424), .B2(new_n426), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n422), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n444), .B1(new_n446), .B2(KEYINPUT16), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n440), .B1(new_n447), .B2(new_n428), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT17), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n448), .A2(new_n449), .A3(new_n418), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n443), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n435), .A2(new_n441), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n416), .A2(G169), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n408), .A2(new_n410), .A3(G179), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(KEYINPUT18), .B1(new_n452), .B2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT79), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n451), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT18), .ZN(new_n460));
  AOI221_X4 g0260(.A(new_n460), .B1(new_n453), .B2(new_n454), .C1(new_n435), .C2(new_n441), .ZN(new_n461));
  NOR3_X1   g0261(.A1(new_n461), .A2(new_n456), .A3(new_n457), .ZN(new_n462));
  OAI21_X1  g0262(.A(KEYINPUT81), .B1(new_n459), .B2(new_n462), .ZN(new_n463));
  OR3_X1    g0263(.A1(new_n459), .A2(new_n462), .A3(KEYINPUT81), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n403), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n265), .A2(G45), .A3(G274), .ZN(new_n466));
  OR2_X1    g0266(.A1(KEYINPUT5), .A2(G41), .ZN(new_n467));
  NAND2_X1  g0267(.A1(KEYINPUT5), .A2(G41), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(G45), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n470), .A2(G1), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n467), .A2(new_n468), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n263), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n469), .B1(new_n473), .B2(G257), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n251), .A2(new_n253), .A3(G244), .A4(new_n254), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT4), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n257), .A2(KEYINPUT4), .A3(G244), .A4(new_n254), .ZN(new_n478));
  NAND2_X1  g0278(.A1(G33), .A2(G283), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n257), .A2(G250), .A3(G1698), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n477), .A2(new_n478), .A3(new_n479), .A4(new_n480), .ZN(new_n481));
  AND3_X1   g0281(.A1(new_n481), .A2(KEYINPUT83), .A3(new_n263), .ZN(new_n482));
  AOI21_X1  g0282(.A(KEYINPUT83), .B1(new_n481), .B2(new_n263), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n315), .B(new_n474), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT6), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n247), .A2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(G107), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n487), .A2(KEYINPUT6), .A3(G97), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(G20), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n283), .A2(G77), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n487), .B1(new_n424), .B2(new_n426), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n287), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n293), .A2(G97), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n265), .A2(G33), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n293), .A2(new_n496), .A3(new_n226), .A4(new_n286), .ZN(new_n497));
  XNOR2_X1  g0297(.A(new_n497), .B(KEYINPUT82), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n495), .B1(new_n498), .B2(G97), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n494), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n481), .A2(new_n263), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(new_n474), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n369), .ZN(new_n503));
  AND3_X1   g0303(.A1(new_n484), .A2(new_n500), .A3(new_n503), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n474), .B1(new_n482), .B2(new_n483), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(KEYINPUT84), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT84), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n507), .B(new_n474), .C1(new_n482), .C2(new_n483), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n506), .A2(G200), .A3(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(new_n502), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n500), .B1(G190), .B2(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n504), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n293), .A2(G107), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT25), .ZN(new_n514));
  XNOR2_X1  g0314(.A(new_n513), .B(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n515), .B1(new_n498), .B2(G107), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT23), .ZN(new_n517));
  NOR3_X1   g0317(.A1(new_n517), .A2(new_n227), .A3(G107), .ZN(new_n518));
  AOI21_X1  g0318(.A(KEYINPUT23), .B1(new_n487), .B2(G20), .ZN(new_n519));
  NAND2_X1  g0319(.A1(G33), .A2(G116), .ZN(new_n520));
  OAI22_X1  g0320(.A1(new_n518), .A2(new_n519), .B1(G20), .B2(new_n520), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n251), .A2(new_n253), .A3(new_n227), .A4(G87), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(KEYINPUT22), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT22), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n257), .A2(new_n524), .A3(new_n227), .A4(G87), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n521), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n287), .B1(new_n526), .B2(KEYINPUT24), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT24), .ZN(new_n528));
  AOI211_X1 g0328(.A(new_n528), .B(new_n521), .C1(new_n523), .C2(new_n525), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n516), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n251), .A2(new_n253), .A3(G250), .A4(new_n254), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n251), .A2(new_n253), .A3(G257), .A4(G1698), .ZN(new_n532));
  NAND2_X1  g0332(.A1(G33), .A2(G294), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n263), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n473), .A2(G264), .ZN(new_n536));
  INV_X1    g0336(.A(new_n469), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(KEYINPUT86), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n263), .A2(new_n534), .B1(new_n473), .B2(G264), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT86), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n540), .A2(new_n541), .A3(new_n537), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n539), .A2(new_n542), .A3(new_n411), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n538), .A2(new_n396), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n530), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n369), .B1(new_n539), .B2(new_n542), .ZN(new_n546));
  INV_X1    g0346(.A(new_n546), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n535), .A2(new_n536), .A3(G179), .A4(new_n537), .ZN(new_n548));
  XNOR2_X1  g0348(.A(new_n548), .B(KEYINPUT87), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n545), .B1(new_n550), .B2(new_n530), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT85), .ZN(new_n552));
  OAI21_X1  g0352(.A(G250), .B1(new_n470), .B2(G1), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n466), .B1(new_n263), .B2(new_n553), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n251), .A2(new_n253), .A3(G238), .A4(new_n254), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n251), .A2(new_n253), .A3(G244), .A4(G1698), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n555), .A2(new_n556), .A3(new_n520), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n554), .B1(new_n557), .B2(new_n263), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n558), .A2(new_n369), .ZN(new_n559));
  AOI211_X1 g0359(.A(new_n315), .B(new_n554), .C1(new_n557), .C2(new_n263), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n552), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n558), .A2(G179), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n562), .B(KEYINPUT85), .C1(new_n369), .C2(new_n558), .ZN(new_n563));
  INV_X1    g0363(.A(new_n376), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n498), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n257), .A2(new_n227), .A3(G68), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT19), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n227), .B1(new_n260), .B2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(G87), .ZN(new_n569));
  INV_X1    g0369(.A(G97), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n569), .A2(new_n570), .A3(new_n487), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n567), .B1(new_n377), .B2(new_n570), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n566), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n574), .A2(new_n287), .B1(new_n294), .B2(new_n376), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n565), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n561), .A2(new_n563), .A3(new_n576), .ZN(new_n577));
  OR2_X1    g0377(.A1(new_n558), .A2(new_n396), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n498), .A2(G87), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n558), .A2(G190), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n578), .A2(new_n579), .A3(new_n575), .A4(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n577), .A2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT21), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n469), .B1(new_n473), .B2(G270), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n251), .A2(new_n253), .A3(G257), .A4(new_n254), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n251), .A2(new_n253), .A3(G264), .A4(G1698), .ZN(new_n586));
  INV_X1    g0386(.A(G303), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n585), .B(new_n586), .C1(new_n587), .C2(new_n257), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n263), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n584), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(G169), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n496), .A2(G116), .ZN(new_n592));
  INV_X1    g0392(.A(new_n297), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n592), .B1(new_n593), .B2(new_n295), .ZN(new_n594));
  INV_X1    g0394(.A(G116), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n294), .A2(new_n595), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n286), .A2(new_n226), .B1(G20), .B2(new_n595), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n479), .B(new_n227), .C1(G33), .C2(new_n570), .ZN(new_n598));
  AND3_X1   g0398(.A1(new_n597), .A2(KEYINPUT20), .A3(new_n598), .ZN(new_n599));
  AOI21_X1  g0399(.A(KEYINPUT20), .B1(new_n597), .B2(new_n598), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n596), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n594), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n583), .B1(new_n591), .B2(new_n602), .ZN(new_n603));
  OAI211_X1 g0403(.A(G116), .B(new_n496), .C1(new_n296), .C2(new_n297), .ZN(new_n604));
  OR2_X1    g0404(.A1(new_n599), .A2(new_n600), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n604), .A2(new_n605), .A3(new_n596), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n606), .A2(KEYINPUT21), .A3(G169), .A4(new_n590), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n590), .A2(G200), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n584), .A2(new_n589), .A3(G190), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n608), .A2(new_n602), .A3(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n584), .A2(new_n589), .A3(G179), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n606), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n603), .A2(new_n607), .A3(new_n610), .A4(new_n613), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n582), .A2(new_n614), .ZN(new_n615));
  AND4_X1   g0415(.A1(new_n465), .A2(new_n512), .A3(new_n551), .A4(new_n615), .ZN(G372));
  NAND2_X1  g0416(.A1(new_n452), .A2(new_n455), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n460), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n452), .A2(KEYINPUT18), .A3(new_n455), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n369), .B1(new_n277), .B2(new_n279), .ZN(new_n622));
  OAI22_X1  g0422(.A1(new_n622), .A2(new_n313), .B1(new_n280), .B2(new_n315), .ZN(new_n623));
  INV_X1    g0423(.A(new_n314), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n304), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT90), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n400), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n389), .A2(new_n390), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n369), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n629), .A2(KEYINPUT90), .A3(new_n398), .A4(new_n399), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n625), .A2(new_n627), .A3(new_n630), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n451), .A2(new_n307), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n621), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n364), .A2(new_n368), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n372), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n465), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n576), .B1(new_n559), .B2(new_n560), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n484), .A2(new_n503), .A3(new_n500), .ZN(new_n639));
  OAI21_X1  g0439(.A(KEYINPUT26), .B1(new_n582), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n484), .A2(new_n503), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT89), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n581), .A2(new_n638), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n484), .A2(KEYINPUT89), .A3(new_n503), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n643), .A2(new_n645), .A3(new_n500), .A4(new_n646), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n638), .B(new_n640), .C1(new_n647), .C2(KEYINPUT26), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT87), .ZN(new_n649));
  XNOR2_X1  g0449(.A(new_n548), .B(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n530), .B1(new_n650), .B2(new_n546), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n603), .A2(new_n607), .A3(new_n613), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n474), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT83), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n501), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n481), .A2(KEYINPUT83), .A3(new_n263), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n655), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(G200), .B1(new_n659), .B2(new_n507), .ZN(new_n660));
  INV_X1    g0460(.A(new_n508), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n511), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n545), .A2(new_n644), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n662), .A2(new_n639), .A3(new_n663), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n654), .B1(new_n664), .B2(KEYINPUT88), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT88), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n512), .A2(new_n666), .A3(new_n663), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n648), .B1(new_n665), .B2(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n636), .B1(new_n637), .B2(new_n668), .ZN(G369));
  AND2_X1   g0469(.A1(new_n227), .A2(G13), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(new_n265), .ZN(new_n671));
  OR2_X1    g0471(.A1(new_n671), .A2(KEYINPUT27), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(KEYINPUT27), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n672), .A2(G213), .A3(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(G343), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n677), .A2(new_n602), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n653), .A2(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n679), .B1(new_n614), .B2(new_n678), .ZN(new_n680));
  AND2_X1   g0480(.A1(new_n680), .A2(G330), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n653), .A2(new_n677), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n543), .A2(new_n544), .ZN(new_n684));
  INV_X1    g0484(.A(new_n530), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n530), .A2(new_n676), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(KEYINPUT91), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT91), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n530), .A2(new_n689), .A3(new_n676), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n651), .A2(new_n686), .A3(new_n688), .A4(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n692), .B1(new_n652), .B2(new_n676), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n682), .B1(new_n683), .B2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  OAI22_X1  g0495(.A1(new_n691), .A2(new_n683), .B1(new_n651), .B2(new_n676), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n695), .A2(new_n697), .ZN(G399));
  INV_X1    g0498(.A(new_n219), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n699), .A2(G41), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n571), .A2(G116), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n701), .A2(G1), .A3(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n703), .B1(new_n224), .B2(new_n701), .ZN(new_n704));
  XNOR2_X1  g0504(.A(new_n704), .B(KEYINPUT28), .ZN(new_n705));
  NOR3_X1   g0505(.A1(new_n582), .A2(KEYINPUT26), .A3(new_n639), .ZN(new_n706));
  INV_X1    g0506(.A(new_n638), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n647), .A2(KEYINPUT26), .ZN(new_n709));
  OAI211_X1 g0509(.A(new_n708), .B(new_n709), .C1(new_n664), .C2(new_n654), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n710), .A2(KEYINPUT29), .A3(new_n677), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n664), .A2(KEYINPUT88), .ZN(new_n712));
  INV_X1    g0512(.A(new_n654), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n712), .A2(new_n667), .A3(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n648), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n676), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n711), .B1(new_n716), .B2(KEYINPUT29), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n540), .A2(new_n558), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n510), .A2(KEYINPUT30), .A3(new_n612), .A4(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT30), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n501), .A2(new_n540), .A3(new_n558), .A4(new_n474), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n720), .B1(new_n721), .B2(new_n611), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n558), .A2(G179), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n723), .A2(new_n538), .A3(new_n590), .ZN(new_n724));
  OAI211_X1 g0524(.A(new_n719), .B(new_n722), .C1(new_n659), .C2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT31), .ZN(new_n726));
  AND3_X1   g0526(.A1(new_n725), .A2(new_n726), .A3(new_n676), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n512), .A2(new_n551), .A3(new_n615), .A4(new_n677), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n726), .B1(new_n725), .B2(new_n676), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n727), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(G330), .ZN(new_n731));
  AND2_X1   g0531(.A1(new_n717), .A2(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n705), .B1(new_n732), .B2(G1), .ZN(G364));
  AOI21_X1  g0533(.A(new_n265), .B1(new_n670), .B2(G45), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  OR3_X1    g0535(.A1(new_n735), .A2(new_n700), .A3(KEYINPUT92), .ZN(new_n736));
  OAI21_X1  g0536(.A(KEYINPUT92), .B1(new_n735), .B2(new_n700), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n396), .A2(G179), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n740), .A2(G20), .A3(new_n411), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(new_n487), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n315), .A2(new_n396), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n743), .A2(G20), .A3(new_n411), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n742), .B1(G68), .B2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n227), .A2(new_n315), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n747), .A2(G190), .A3(new_n396), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n746), .B1(new_n202), .B2(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(G190), .A2(G200), .ZN(new_n750));
  AND2_X1   g0550(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n257), .B1(new_n752), .B2(new_n375), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n227), .A2(new_n411), .ZN(new_n754));
  AND2_X1   g0554(.A1(new_n743), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n754), .A2(new_n740), .ZN(new_n757));
  OAI22_X1  g0557(.A1(new_n756), .A2(new_n201), .B1(new_n757), .B2(new_n569), .ZN(new_n758));
  NOR3_X1   g0558(.A1(new_n749), .A2(new_n753), .A3(new_n758), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n750), .A2(G20), .A3(new_n315), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(G159), .ZN(new_n762));
  XNOR2_X1  g0562(.A(new_n762), .B(KEYINPUT32), .ZN(new_n763));
  NOR3_X1   g0563(.A1(new_n411), .A2(G179), .A3(G200), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n227), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n763), .B1(G97), .B2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n748), .ZN(new_n768));
  INV_X1    g0568(.A(new_n741), .ZN(new_n769));
  AOI22_X1  g0569(.A1(G322), .A2(new_n768), .B1(new_n769), .B2(G283), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n257), .B1(new_n755), .B2(G326), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n772), .B1(G294), .B2(new_n766), .ZN(new_n773));
  AOI22_X1  g0573(.A1(new_n751), .A2(G311), .B1(new_n761), .B2(G329), .ZN(new_n774));
  XOR2_X1   g0574(.A(KEYINPUT33), .B(G317), .Z(new_n775));
  OAI21_X1  g0575(.A(new_n774), .B1(new_n744), .B2(new_n775), .ZN(new_n776));
  AND2_X1   g0576(.A1(new_n757), .A2(KEYINPUT94), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n757), .A2(KEYINPUT94), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n776), .B1(G303), .B2(new_n780), .ZN(new_n781));
  AOI22_X1  g0581(.A1(new_n759), .A2(new_n767), .B1(new_n773), .B2(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n226), .B1(G20), .B2(new_n369), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n739), .B1(new_n782), .B2(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(G13), .A2(G33), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(G20), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(new_n783), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n425), .A2(new_n219), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n790), .B1(new_n470), .B2(new_n225), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(KEYINPUT93), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n792), .B1(new_n245), .B2(new_n470), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n699), .A2(new_n425), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n794), .A2(G355), .B1(new_n595), .B2(new_n699), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n785), .B1(new_n789), .B2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n788), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n797), .B1(new_n680), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n682), .A2(new_n738), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n680), .A2(G330), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n799), .B1(new_n800), .B2(new_n801), .ZN(G396));
  NAND2_X1  g0602(.A1(new_n399), .A2(new_n676), .ZN(new_n803));
  AND3_X1   g0603(.A1(new_n397), .A2(new_n400), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n627), .A2(new_n630), .ZN(new_n805));
  INV_X1    g0605(.A(new_n803), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n804), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n716), .B(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n739), .B1(new_n809), .B2(new_n731), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n810), .B1(new_n731), .B2(new_n809), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n783), .A2(new_n786), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n739), .B1(G77), .B2(new_n813), .ZN(new_n814));
  XOR2_X1   g0614(.A(new_n814), .B(KEYINPUT95), .Z(new_n815));
  NOR2_X1   g0615(.A1(new_n779), .A2(new_n487), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n768), .A2(G294), .B1(new_n751), .B2(G116), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n257), .B1(new_n761), .B2(G311), .ZN(new_n818));
  OAI211_X1 g0618(.A(new_n817), .B(new_n818), .C1(new_n570), .C2(new_n765), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n741), .A2(new_n569), .ZN(new_n820));
  INV_X1    g0620(.A(G283), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n756), .A2(new_n587), .B1(new_n821), .B2(new_n744), .ZN(new_n822));
  NOR4_X1   g0622(.A1(new_n816), .A2(new_n819), .A3(new_n820), .A4(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  OR2_X1    g0624(.A1(new_n824), .A2(KEYINPUT96), .ZN(new_n825));
  AOI22_X1  g0625(.A1(G137), .A2(new_n755), .B1(new_n751), .B2(G159), .ZN(new_n826));
  INV_X1    g0626(.A(G143), .ZN(new_n827));
  INV_X1    g0627(.A(G150), .ZN(new_n828));
  OAI221_X1 g0628(.A(new_n826), .B1(new_n827), .B2(new_n748), .C1(new_n828), .C2(new_n744), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n829), .B(KEYINPUT34), .ZN(new_n830));
  INV_X1    g0630(.A(G132), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n257), .B1(new_n760), .B2(new_n831), .C1(new_n741), .C2(new_n203), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n832), .B1(G58), .B2(new_n766), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n830), .B(new_n833), .C1(new_n201), .C2(new_n779), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n824), .A2(KEYINPUT96), .ZN(new_n835));
  AND3_X1   g0635(.A1(new_n825), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n815), .B1(new_n836), .B2(new_n784), .C1(new_n808), .C2(new_n787), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n811), .A2(new_n837), .ZN(G384));
  XNOR2_X1  g0638(.A(new_n489), .B(KEYINPUT97), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT35), .ZN(new_n840));
  OR2_X1    g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n839), .A2(new_n840), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n841), .A2(new_n842), .A3(G116), .A4(new_n228), .ZN(new_n843));
  XOR2_X1   g0643(.A(new_n843), .B(KEYINPUT36), .Z(new_n844));
  OAI211_X1 g0644(.A(new_n225), .B(G77), .C1(new_n202), .C2(new_n300), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n201), .A2(G68), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n265), .B(G13), .C1(new_n845), .C2(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n637), .A2(new_n731), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n449), .B1(new_n448), .B2(new_n418), .ZN(new_n850));
  AND4_X1   g0650(.A1(new_n449), .A2(new_n418), .A3(new_n435), .A4(new_n441), .ZN(new_n851));
  OAI22_X1  g0651(.A1(new_n850), .A2(new_n851), .B1(new_n461), .B2(new_n456), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n448), .A2(new_n674), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AND3_X1   g0654(.A1(new_n428), .A2(new_n287), .A3(new_n434), .ZN(new_n855));
  INV_X1    g0655(.A(new_n674), .ZN(new_n856));
  OAI22_X1  g0656(.A1(new_n855), .A2(new_n440), .B1(new_n455), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n442), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(KEYINPUT37), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT37), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n857), .A2(new_n860), .A3(new_n442), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(KEYINPUT38), .B1(new_n854), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n419), .B1(new_n422), .B2(new_n445), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n864), .A2(new_n434), .A3(new_n287), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n441), .ZN(new_n866));
  AOI21_X1  g0666(.A(KEYINPUT98), .B1(new_n866), .B2(new_n856), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT98), .ZN(new_n868));
  AOI211_X1 g0668(.A(new_n868), .B(new_n674), .C1(new_n865), .C2(new_n441), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  AOI22_X1  g0670(.A1(new_n443), .A2(new_n450), .B1(new_n456), .B2(new_n457), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n618), .A2(KEYINPUT79), .A3(new_n619), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  AND3_X1   g0673(.A1(new_n857), .A2(new_n860), .A3(new_n442), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n448), .A2(new_n418), .B1(new_n866), .B2(new_n455), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n440), .B1(new_n447), .B2(new_n864), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n868), .B1(new_n876), .B2(new_n674), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n866), .A2(KEYINPUT98), .A3(new_n856), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n875), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n874), .B1(new_n879), .B2(KEYINPUT37), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n873), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n863), .B1(new_n881), .B2(KEYINPUT38), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n304), .A2(new_n676), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n625), .A2(new_n307), .A3(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n316), .A2(new_n304), .A3(new_n676), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n730), .A2(new_n886), .A3(new_n808), .ZN(new_n887));
  OAI21_X1  g0687(.A(KEYINPUT40), .B1(new_n882), .B2(new_n887), .ZN(new_n888));
  OAI22_X1  g0688(.A1(new_n459), .A2(new_n462), .B1(new_n867), .B2(new_n869), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n866), .A2(new_n455), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n442), .ZN(new_n891));
  NOR3_X1   g0691(.A1(new_n891), .A2(new_n867), .A3(new_n869), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n861), .B1(new_n892), .B2(new_n860), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n889), .A2(KEYINPUT38), .A3(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT38), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n895), .B1(new_n873), .B2(new_n880), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT40), .ZN(new_n898));
  AOI211_X1 g0698(.A(new_n727), .B(new_n807), .C1(new_n728), .C2(new_n729), .ZN(new_n899));
  NAND4_X1  g0699(.A1(new_n897), .A2(new_n898), .A3(new_n886), .A4(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n888), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n849), .B1(new_n901), .B2(G330), .ZN(new_n902));
  AND2_X1   g0702(.A1(new_n465), .A2(new_n730), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n902), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  AOI211_X1 g0704(.A(new_n676), .B(new_n807), .C1(new_n714), .C2(new_n715), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n400), .A2(new_n676), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n897), .B(new_n886), .C1(new_n905), .C2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n621), .A2(new_n674), .ZN(new_n908));
  INV_X1    g0708(.A(new_n625), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n677), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  NOR3_X1   g0711(.A1(new_n873), .A2(new_n880), .A3(new_n895), .ZN(new_n912));
  NOR3_X1   g0712(.A1(new_n912), .A2(KEYINPUT39), .A3(new_n863), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT39), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n914), .B1(new_n894), .B2(new_n896), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n911), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  AND3_X1   g0716(.A1(new_n907), .A2(new_n908), .A3(new_n916), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n904), .B(new_n917), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n465), .B(new_n711), .C1(new_n716), .C2(KEYINPUT29), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT99), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT29), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n668), .B2(new_n676), .ZN(new_n923));
  NAND4_X1  g0723(.A1(new_n923), .A2(KEYINPUT99), .A3(new_n465), .A4(new_n711), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n635), .B1(new_n921), .B2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  OAI22_X1  g0726(.A1(new_n918), .A2(new_n926), .B1(new_n265), .B2(new_n670), .ZN(new_n927));
  AND2_X1   g0727(.A1(new_n918), .A2(new_n926), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n848), .B1(new_n927), .B2(new_n928), .ZN(G367));
  NAND2_X1  g0729(.A1(new_n579), .A2(new_n575), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n676), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n645), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n638), .B2(new_n931), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(KEYINPUT43), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n500), .A2(new_n676), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n512), .A2(new_n935), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n643), .A2(new_n500), .A3(new_n646), .A4(new_n676), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n652), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n676), .B1(new_n939), .B2(new_n639), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n691), .A2(new_n683), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(new_n512), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(KEYINPUT42), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT42), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n941), .A2(new_n944), .A3(new_n512), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n934), .B1(new_n940), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(KEYINPUT100), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT100), .ZN(new_n949));
  OAI211_X1 g0749(.A(new_n949), .B(new_n934), .C1(new_n940), .C2(new_n946), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n951), .B1(KEYINPUT43), .B2(new_n933), .ZN(new_n952));
  AND2_X1   g0752(.A1(new_n936), .A2(new_n937), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n695), .A2(new_n953), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n933), .A2(KEYINPUT43), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n948), .A2(new_n955), .A3(new_n950), .ZN(new_n956));
  AND3_X1   g0756(.A1(new_n952), .A2(new_n954), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n954), .B1(new_n952), .B2(new_n956), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  XOR2_X1   g0759(.A(KEYINPUT101), .B(KEYINPUT41), .Z(new_n960));
  XOR2_X1   g0760(.A(new_n700), .B(new_n960), .Z(new_n961));
  INV_X1    g0761(.A(KEYINPUT44), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT102), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n963), .B1(new_n953), .B2(new_n696), .ZN(new_n964));
  NAND4_X1  g0764(.A1(new_n696), .A2(new_n963), .A3(new_n936), .A4(new_n937), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n962), .B1(new_n964), .B2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT45), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n953), .B2(new_n696), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n697), .A2(new_n938), .A3(KEYINPUT45), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(KEYINPUT102), .B1(new_n697), .B2(new_n938), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n972), .A2(KEYINPUT44), .A3(new_n965), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n967), .A2(new_n971), .A3(new_n695), .A4(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT103), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n971), .A2(new_n973), .ZN(new_n977));
  AOI21_X1  g0777(.A(KEYINPUT44), .B1(new_n972), .B2(new_n965), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n694), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n976), .A2(new_n979), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n975), .B(new_n694), .C1(new_n977), .C2(new_n978), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT104), .ZN(new_n982));
  INV_X1    g0782(.A(new_n941), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n682), .A2(new_n693), .A3(new_n683), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n695), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n982), .B1(new_n732), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n717), .A2(new_n731), .ZN(new_n988));
  NOR3_X1   g0788(.A1(new_n988), .A2(KEYINPUT104), .A3(new_n985), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n980), .B(new_n981), .C1(new_n987), .C2(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n961), .B1(new_n990), .B2(new_n732), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n959), .B1(new_n991), .B2(new_n735), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n239), .A2(new_n790), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n789), .B1(new_n219), .B2(new_n376), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n739), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(G159), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n752), .A2(new_n201), .B1(new_n996), .B2(new_n744), .ZN(new_n997));
  INV_X1    g0797(.A(new_n757), .ZN(new_n998));
  AOI211_X1 g0798(.A(new_n425), .B(new_n997), .C1(G58), .C2(new_n998), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n768), .A2(G150), .B1(G137), .B2(new_n761), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(G77), .A2(new_n769), .B1(new_n755), .B2(G143), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n766), .A2(G68), .ZN(new_n1002));
  NAND4_X1  g0802(.A1(new_n999), .A2(new_n1000), .A3(new_n1001), .A4(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(G311), .ZN(new_n1004));
  OAI22_X1  g0804(.A1(new_n756), .A2(new_n1004), .B1(new_n587), .B2(new_n748), .ZN(new_n1005));
  AOI211_X1 g0805(.A(new_n257), .B(new_n1005), .C1(G317), .C2(new_n761), .ZN(new_n1006));
  INV_X1    g0806(.A(G294), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n744), .A2(new_n1007), .B1(new_n741), .B2(new_n570), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1008), .B1(G283), .B2(new_n751), .ZN(new_n1009));
  OAI211_X1 g0809(.A(new_n1006), .B(new_n1009), .C1(new_n487), .C2(new_n765), .ZN(new_n1010));
  NOR3_X1   g0810(.A1(new_n757), .A2(KEYINPUT46), .A3(new_n595), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n780), .A2(G116), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1011), .B1(new_n1012), .B2(KEYINPUT46), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1003), .B1(new_n1010), .B2(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n1015));
  OR2_X1    g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n784), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n995), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(new_n798), .B2(new_n933), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n992), .A2(new_n1019), .ZN(G387));
  NAND2_X1  g0820(.A1(new_n693), .A2(new_n788), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n794), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n1022), .A2(new_n702), .B1(G107), .B2(new_n219), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n236), .A2(G45), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n470), .B1(new_n203), .B2(new_n375), .C1(new_n702), .C2(KEYINPUT106), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(KEYINPUT106), .B2(new_n702), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n436), .A2(G50), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT50), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n790), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1023), .B1(new_n1024), .B2(new_n1029), .ZN(new_n1030));
  AND2_X1   g0830(.A1(new_n1030), .A2(KEYINPUT107), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n789), .B1(new_n1030), .B2(KEYINPUT107), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n739), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n748), .A2(new_n201), .B1(new_n828), .B2(new_n760), .ZN(new_n1034));
  AOI211_X1 g0834(.A(new_n425), .B(new_n1034), .C1(G97), .C2(new_n769), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n745), .A2(new_n437), .B1(new_n755), .B2(G159), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(G77), .A2(new_n998), .B1(new_n751), .B2(G68), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n766), .A2(new_n564), .ZN(new_n1038));
  NAND4_X1  g0838(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .A4(new_n1038), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(G322), .A2(new_n755), .B1(new_n751), .B2(G303), .ZN(new_n1040));
  INV_X1    g0840(.A(G317), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n1040), .B1(new_n1004), .B2(new_n744), .C1(new_n1041), .C2(new_n748), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT48), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n1043), .B1(new_n821), .B2(new_n765), .C1(new_n1007), .C2(new_n757), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT108), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT49), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n425), .B1(new_n741), .B2(new_n595), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(G326), .B2(new_n761), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1039), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1033), .B1(new_n1052), .B2(new_n783), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n1021), .A2(new_n1053), .B1(new_n986), .B2(new_n735), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n732), .A2(new_n986), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1055), .A2(new_n700), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n732), .A2(new_n986), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1054), .B1(new_n1056), .B2(new_n1057), .ZN(G393));
  NAND2_X1  g0858(.A1(new_n979), .A2(new_n974), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n701), .B1(new_n1059), .B2(new_n1055), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n990), .A2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n979), .A2(new_n735), .A3(new_n974), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n248), .A2(new_n790), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n789), .B1(new_n570), .B2(new_n219), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n739), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n756), .A2(new_n828), .B1(new_n996), .B2(new_n748), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT51), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n766), .A2(G77), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n752), .A2(new_n436), .B1(new_n201), .B2(new_n744), .ZN(new_n1069));
  NOR3_X1   g0869(.A1(new_n1069), .A2(new_n425), .A3(new_n820), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n757), .A2(new_n300), .B1(new_n760), .B2(new_n827), .ZN(new_n1071));
  XOR2_X1   g0871(.A(new_n1071), .B(KEYINPUT109), .Z(new_n1072));
  NAND4_X1  g0872(.A1(new_n1067), .A2(new_n1068), .A3(new_n1070), .A4(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT110), .ZN(new_n1074));
  OR2_X1    g0874(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n756), .A2(new_n1041), .B1(new_n1004), .B2(new_n748), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT52), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n745), .A2(G303), .B1(new_n998), .B2(G283), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n751), .A2(G294), .B1(new_n761), .B2(G322), .ZN(new_n1079));
  AOI211_X1 g0879(.A(new_n257), .B(new_n742), .C1(G116), .C2(new_n766), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n1077), .A2(new_n1078), .A3(new_n1079), .A4(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1075), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1065), .B1(new_n1083), .B2(new_n783), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1084), .B1(new_n938), .B2(new_n798), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1061), .A2(new_n1062), .A3(new_n1085), .ZN(G390));
  NAND3_X1  g0886(.A1(new_n899), .A2(G330), .A3(new_n886), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n897), .A2(KEYINPUT39), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n854), .A2(new_n862), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(new_n895), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n894), .A2(new_n1091), .A3(new_n914), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1089), .A2(new_n1092), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n886), .B1(new_n905), .B2(new_n906), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1093), .B1(new_n1094), .B2(new_n910), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n886), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n710), .A2(new_n677), .A3(new_n808), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n906), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1096), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n910), .B1(new_n912), .B2(new_n863), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1088), .B1(new_n1095), .B2(new_n1101), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n913), .A2(new_n915), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n714), .A2(new_n715), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1104), .A2(new_n677), .A3(new_n808), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1096), .B1(new_n1105), .B2(new_n1098), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1103), .B1(new_n1106), .B2(new_n911), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1101), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1107), .A2(new_n1087), .A3(new_n1108), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1102), .A2(new_n735), .A3(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(KEYINPUT111), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT111), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n1102), .A2(new_n1112), .A3(new_n1109), .A4(new_n735), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n899), .A2(G330), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(new_n1096), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n1116), .A2(new_n1087), .A3(new_n1098), .A4(new_n1097), .ZN(new_n1117));
  AND2_X1   g0917(.A1(new_n1116), .A2(new_n1087), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n906), .B1(new_n716), .B2(new_n808), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1117), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n849), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1120), .A2(new_n925), .A3(new_n1121), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n910), .B1(new_n1119), .B2(new_n1096), .ZN(new_n1123));
  AOI211_X1 g0923(.A(new_n1088), .B(new_n1101), .C1(new_n1123), .C2(new_n1103), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1087), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1122), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  AOI211_X1 g0926(.A(new_n635), .B(new_n849), .C1(new_n921), .C2(new_n924), .ZN(new_n1127));
  NAND4_X1  g0927(.A1(new_n1102), .A2(new_n1127), .A3(new_n1109), .A4(new_n1120), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1126), .A2(new_n1128), .A3(new_n700), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n738), .B1(new_n436), .B2(new_n812), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n757), .A2(new_n828), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1131), .B(KEYINPUT53), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(KEYINPUT54), .B(G143), .ZN(new_n1133));
  INV_X1    g0933(.A(G137), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n752), .A2(new_n1133), .B1(new_n1134), .B2(new_n744), .ZN(new_n1135));
  XOR2_X1   g0935(.A(new_n1135), .B(KEYINPUT112), .Z(new_n1136));
  INV_X1    g0936(.A(G125), .ZN(new_n1137));
  OAI221_X1 g0937(.A(new_n257), .B1(new_n760), .B2(new_n1137), .C1(new_n741), .C2(new_n201), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(G159), .B2(new_n766), .ZN(new_n1139));
  INV_X1    g0939(.A(G128), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n756), .A2(new_n1140), .B1(new_n831), .B2(new_n748), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(new_n1141), .B(KEYINPUT113), .ZN(new_n1142));
  AND4_X1   g0942(.A1(new_n1132), .A2(new_n1136), .A3(new_n1139), .A4(new_n1142), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n425), .B1(new_n779), .B2(new_n569), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n1144), .B(KEYINPUT114), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n745), .A2(G107), .B1(new_n751), .B2(G97), .ZN(new_n1146));
  OAI221_X1 g0946(.A(new_n1146), .B1(new_n595), .B2(new_n748), .C1(new_n1007), .C2(new_n760), .ZN(new_n1147));
  OAI221_X1 g0947(.A(new_n1068), .B1(new_n203), .B2(new_n741), .C1(new_n821), .C2(new_n756), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1143), .B1(new_n1145), .B2(new_n1149), .ZN(new_n1150));
  OAI221_X1 g0950(.A(new_n1130), .B1(new_n784), .B2(new_n1150), .C1(new_n1093), .C2(new_n787), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1114), .A2(new_n1129), .A3(new_n1151), .ZN(G378));
  XNOR2_X1  g0952(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(KEYINPUT118), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n373), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n371), .A2(new_n856), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n364), .A2(new_n368), .A3(KEYINPUT118), .A4(new_n372), .ZN(new_n1158));
  AND3_X1   g0958(.A1(new_n1156), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1157), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1154), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1157), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1156), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1164), .A2(new_n1153), .A3(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1161), .A2(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1168), .A2(new_n787), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n756), .A2(new_n595), .B1(new_n752), .B2(new_n376), .ZN(new_n1170));
  OAI221_X1 g0970(.A(new_n1002), .B1(new_n487), .B2(new_n748), .C1(new_n821), .C2(new_n760), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n1170), .B(new_n1171), .C1(G97), .C2(new_n745), .ZN(new_n1172));
  OR2_X1    g0972(.A1(new_n257), .A2(G41), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(G77), .B2(new_n998), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(new_n1174), .B(KEYINPUT116), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n741), .A2(new_n202), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n1176), .B(KEYINPUT115), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1172), .A2(new_n1175), .A3(new_n1177), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(KEYINPUT117), .B(KEYINPUT58), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  OR2_X1    g0980(.A1(new_n1178), .A2(new_n1180), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n1140), .A2(new_n748), .B1(new_n744), .B2(new_n831), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n751), .A2(G137), .ZN(new_n1183));
  OAI221_X1 g0983(.A(new_n1183), .B1(new_n757), .B2(new_n1133), .C1(new_n756), .C2(new_n1137), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n1182), .B(new_n1184), .C1(G150), .C2(new_n766), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT59), .ZN(new_n1186));
  OR2_X1    g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n769), .A2(G159), .ZN(new_n1189));
  AOI211_X1 g0989(.A(G33), .B(G41), .C1(new_n761), .C2(G124), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1187), .A2(new_n1188), .A3(new_n1189), .A4(new_n1190), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n1173), .B(new_n201), .C1(G33), .C2(G41), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1178), .A2(new_n1180), .ZN(new_n1193));
  AND4_X1   g0993(.A1(new_n1181), .A2(new_n1191), .A3(new_n1192), .A4(new_n1193), .ZN(new_n1194));
  OAI221_X1 g0994(.A(new_n739), .B1(G50), .B2(new_n813), .C1(new_n1194), .C2(new_n784), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1169), .A2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT119), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1168), .B1(new_n901), .B2(G330), .ZN(new_n1198));
  INV_X1    g0998(.A(G330), .ZN(new_n1199));
  AOI211_X1 g0999(.A(new_n1199), .B(new_n1167), .C1(new_n888), .C2(new_n900), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1197), .B1(new_n1198), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1201), .A2(new_n917), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n907), .A2(new_n908), .A3(new_n916), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1197), .B(new_n1203), .C1(new_n1198), .C2(new_n1200), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1202), .A2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1196), .B1(new_n1205), .B2(new_n735), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1127), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1207), .B1(new_n1208), .B2(new_n1120), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1203), .B1(new_n1198), .B2(new_n1200), .ZN(new_n1210));
  OAI211_X1 g1010(.A(new_n899), .B(new_n886), .C1(new_n912), .C2(new_n863), .ZN(new_n1211));
  AND3_X1   g1011(.A1(new_n730), .A2(new_n886), .A3(new_n808), .ZN(new_n1212));
  AOI21_X1  g1012(.A(KEYINPUT40), .B1(new_n894), .B2(new_n896), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n1211), .A2(KEYINPUT40), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1167), .B1(new_n1214), .B2(new_n1199), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n901), .A2(G330), .A3(new_n1168), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n917), .A2(new_n1215), .A3(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1210), .A2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(KEYINPUT57), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n700), .B1(new_n1209), .B2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1128), .A2(new_n1127), .ZN(new_n1221));
  AOI21_X1  g1021(.A(KEYINPUT57), .B1(new_n1205), .B2(new_n1221), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1206), .B1(new_n1220), .B2(new_n1222), .ZN(G375));
  OAI21_X1  g1023(.A(new_n425), .B1(new_n741), .B2(new_n375), .ZN(new_n1224));
  XOR2_X1   g1024(.A(new_n1224), .B(KEYINPUT122), .Z(new_n1225));
  AOI22_X1  g1025(.A1(new_n745), .A2(G116), .B1(new_n751), .B2(G107), .ZN(new_n1226));
  OAI221_X1 g1026(.A(new_n1225), .B1(KEYINPUT121), .B2(new_n1226), .C1(new_n570), .C2(new_n779), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n564), .A2(new_n766), .B1(new_n768), .B2(G283), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1229), .A2(KEYINPUT123), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(KEYINPUT123), .ZN(new_n1231));
  OAI22_X1  g1031(.A1(new_n756), .A2(new_n1007), .B1(new_n587), .B2(new_n760), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(new_n1226), .B2(KEYINPUT121), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1231), .A2(new_n1233), .ZN(new_n1234));
  NOR3_X1   g1034(.A1(new_n1227), .A2(new_n1230), .A3(new_n1234), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1177), .B1(new_n996), .B2(new_n779), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n752), .A2(new_n828), .B1(new_n1134), .B2(new_n748), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n756), .A2(new_n831), .B1(new_n1140), .B2(new_n760), .ZN(new_n1238));
  OAI221_X1 g1038(.A(new_n257), .B1(new_n744), .B2(new_n1133), .C1(new_n201), .C2(new_n765), .ZN(new_n1239));
  NOR4_X1   g1039(.A1(new_n1236), .A2(new_n1237), .A3(new_n1238), .A4(new_n1239), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n783), .B1(new_n1235), .B2(new_n1240), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1241), .B(new_n739), .C1(G68), .C2(new_n813), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(new_n1096), .B2(new_n786), .ZN(new_n1243));
  XNOR2_X1  g1043(.A(new_n734), .B(KEYINPUT120), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1243), .B1(new_n1120), .B2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n961), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1122), .A2(new_n1246), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1127), .A2(new_n1120), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1245), .B1(new_n1247), .B2(new_n1248), .ZN(G381));
  AND3_X1   g1049(.A1(new_n1114), .A2(new_n1129), .A3(new_n1151), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n1250), .B(new_n1206), .C1(new_n1222), .C2(new_n1220), .ZN(new_n1251));
  OR2_X1    g1051(.A1(G393), .A2(G396), .ZN(new_n1252));
  OR4_X1    g1052(.A1(G384), .A2(G390), .A3(new_n1252), .A4(G381), .ZN(new_n1253));
  OR3_X1    g1053(.A1(new_n1251), .A2(new_n1253), .A3(G387), .ZN(G407));
  NAND2_X1  g1054(.A1(new_n675), .A2(G213), .ZN(new_n1255));
  OR2_X1    g1055(.A1(new_n1251), .A2(new_n1255), .ZN(new_n1256));
  OR2_X1    g1056(.A1(new_n1256), .A2(KEYINPUT124), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1256), .A2(KEYINPUT124), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1257), .A2(G213), .A3(G407), .A4(new_n1258), .ZN(G409));
  INV_X1    g1059(.A(KEYINPUT126), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(G375), .A2(G378), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1255), .ZN(new_n1262));
  NOR3_X1   g1062(.A1(new_n1198), .A2(new_n1200), .A3(new_n1203), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(new_n1093), .A2(new_n911), .B1(new_n621), .B2(new_n674), .ZN(new_n1264));
  AOI22_X1  g1064(.A1(new_n1215), .A2(new_n1216), .B1(new_n907), .B2(new_n1264), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1244), .B1(new_n1263), .B2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1196), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n1202), .A2(new_n1204), .B1(new_n1128), .B2(new_n1127), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1268), .B1(new_n1269), .B2(new_n1246), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1262), .B1(new_n1250), .B2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1248), .A2(KEYINPUT60), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT60), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1273), .B1(new_n1127), .B2(new_n1120), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n701), .B1(new_n1127), .B2(new_n1120), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1272), .A2(new_n1274), .A3(new_n1275), .ZN(new_n1276));
  AND3_X1   g1076(.A1(new_n1276), .A2(G384), .A3(new_n1245), .ZN(new_n1277));
  AOI21_X1  g1077(.A(G384), .B1(new_n1276), .B2(new_n1245), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1261), .A2(new_n1271), .A3(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT63), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1261), .A2(new_n1271), .A3(new_n1279), .A4(KEYINPUT63), .ZN(new_n1283));
  XOR2_X1   g1083(.A(G393), .B(G396), .Z(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  AND3_X1   g1085(.A1(new_n992), .A2(new_n1019), .A3(G390), .ZN(new_n1286));
  AOI21_X1  g1086(.A(G390), .B1(new_n992), .B2(new_n1019), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1285), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(G390), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(G387), .A2(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n992), .A2(new_n1019), .A3(G390), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1290), .A2(new_n1284), .A3(new_n1291), .ZN(new_n1292));
  AND2_X1   g1092(.A1(new_n1288), .A2(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1282), .A2(new_n1283), .A3(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1261), .A2(new_n1271), .ZN(new_n1295));
  OR2_X1    g1095(.A1(new_n1255), .A2(KEYINPUT125), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1262), .A2(G2897), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1279), .A2(new_n1296), .A3(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1276), .A2(new_n1245), .ZN(new_n1299));
  INV_X1    g1099(.A(G384), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1276), .A2(G384), .A3(new_n1245), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1301), .A2(new_n1302), .A3(new_n1296), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1297), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1295), .A2(new_n1298), .A3(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT61), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1260), .B1(new_n1294), .B2(new_n1308), .ZN(new_n1309));
  AND3_X1   g1109(.A1(new_n1283), .A2(new_n1292), .A3(new_n1288), .ZN(new_n1310));
  AOI22_X1  g1110(.A1(new_n1261), .A2(new_n1271), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1311));
  AOI21_X1  g1111(.A(KEYINPUT61), .B1(new_n1311), .B2(new_n1298), .ZN(new_n1312));
  NAND4_X1  g1112(.A1(new_n1310), .A2(new_n1312), .A3(KEYINPUT126), .A4(new_n1282), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1309), .A2(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1288), .A2(new_n1292), .ZN(new_n1315));
  XNOR2_X1  g1115(.A(new_n1280), .B(KEYINPUT62), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1315), .B1(new_n1316), .B2(new_n1308), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1314), .A2(new_n1317), .ZN(G405));
  NAND2_X1  g1118(.A1(new_n1261), .A2(new_n1251), .ZN(new_n1319));
  XOR2_X1   g1119(.A(new_n1319), .B(new_n1279), .Z(new_n1320));
  NAND3_X1  g1120(.A1(new_n1320), .A2(KEYINPUT127), .A3(new_n1315), .ZN(new_n1321));
  XNOR2_X1  g1121(.A(new_n1315), .B(KEYINPUT127), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1321), .B1(new_n1320), .B2(new_n1322), .ZN(G402));
endmodule


