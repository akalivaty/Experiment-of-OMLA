//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 0 1 1 1 1 1 0 1 0 0 0 0 0 1 1 0 0 0 0 0 0 1 0 1 1 0 1 0 0 0 0 0 0 0 0 0 0 0 0 1 0 1 1 0 1 1 0 1 0 0 0 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:21 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1246, new_n1247, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0006(.A1(G68), .A2(G238), .B1(G97), .B2(G257), .ZN(new_n207));
  NAND2_X1  g0007(.A1(G50), .A2(G226), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G116), .A2(G270), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G58), .A2(G232), .ZN(new_n210));
  NAND4_X1  g0010(.A1(new_n207), .A2(new_n208), .A3(new_n209), .A4(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(G77), .ZN(new_n212));
  INV_X1    g0012(.A(G244), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  AND2_X1   g0014(.A1(G87), .A2(G250), .ZN(new_n215));
  NOR3_X1   g0015(.A1(new_n211), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G107), .A2(G264), .ZN(new_n217));
  INV_X1    g0017(.A(G1), .ZN(new_n218));
  INV_X1    g0018(.A(G20), .ZN(new_n219));
  OAI21_X1  g0019(.A(KEYINPUT64), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  OR3_X1    g0020(.A1(new_n218), .A2(new_n219), .A3(KEYINPUT64), .ZN(new_n221));
  AOI22_X1  g0021(.A1(new_n216), .A2(new_n217), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT1), .Z(new_n223));
  NAND2_X1  g0023(.A1(new_n221), .A2(new_n220), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n224), .A2(G13), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n225), .B(G250), .C1(G257), .C2(G264), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT0), .Z(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n228), .A2(new_n219), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n202), .A2(new_n203), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(G50), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  AOI211_X1 g0032(.A(new_n223), .B(new_n227), .C1(new_n229), .C2(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G250), .B(G257), .Z(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XNOR2_X1  g0041(.A(G68), .B(G77), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT65), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G87), .B(G97), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(KEYINPUT66), .B(G107), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n245), .B(new_n249), .ZN(G351));
  INV_X1    g0050(.A(KEYINPUT18), .ZN(new_n251));
  XNOR2_X1  g0051(.A(KEYINPUT8), .B(G58), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n218), .A2(G13), .A3(G20), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g0056(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(new_n228), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n258), .B1(new_n218), .B2(G20), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n256), .B1(new_n260), .B2(new_n253), .ZN(new_n261));
  INV_X1    g0061(.A(new_n258), .ZN(new_n262));
  AND2_X1   g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  NOR2_X1   g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  AOI21_X1  g0065(.A(KEYINPUT7), .B1(new_n265), .B2(new_n219), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT7), .ZN(new_n267));
  NOR4_X1   g0067(.A1(new_n263), .A2(new_n264), .A3(new_n267), .A4(G20), .ZN(new_n268));
  OAI21_X1  g0068(.A(G68), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  NOR2_X1   g0069(.A1(G20), .A2(G33), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G159), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(G58), .A2(G68), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n219), .B1(new_n230), .B2(new_n274), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n269), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT16), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n262), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT73), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n276), .A2(new_n280), .ZN(new_n281));
  OAI21_X1  g0081(.A(KEYINPUT73), .B1(new_n273), .B2(new_n275), .ZN(new_n282));
  NAND4_X1  g0082(.A1(new_n269), .A2(new_n281), .A3(KEYINPUT16), .A4(new_n282), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n261), .B1(new_n279), .B2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G33), .ZN(new_n285));
  INV_X1    g0085(.A(G41), .ZN(new_n286));
  OAI211_X1 g0086(.A(G1), .B(G13), .C1(new_n285), .C2(new_n286), .ZN(new_n287));
  OR2_X1    g0087(.A1(G223), .A2(G1698), .ZN(new_n288));
  INV_X1    g0088(.A(G226), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G1698), .ZN(new_n290));
  OAI211_X1 g0090(.A(new_n288), .B(new_n290), .C1(new_n263), .C2(new_n264), .ZN(new_n291));
  INV_X1    g0091(.A(G87), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n285), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n287), .B1(new_n291), .B2(new_n294), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n218), .B1(G41), .B2(G45), .ZN(new_n296));
  INV_X1    g0096(.A(G274), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G179), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n287), .A2(G232), .A3(new_n296), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n299), .A2(KEYINPUT74), .A3(new_n300), .A4(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT74), .ZN(new_n303));
  INV_X1    g0103(.A(new_n298), .ZN(new_n304));
  NOR2_X1   g0104(.A1(G223), .A2(G1698), .ZN(new_n305));
  OR2_X1    g0105(.A1(KEYINPUT3), .A2(G33), .ZN(new_n306));
  NAND2_X1  g0106(.A1(KEYINPUT3), .A2(G33), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n305), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n293), .B1(new_n308), .B2(new_n290), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n301), .B(new_n304), .C1(new_n309), .C2(new_n287), .ZN(new_n310));
  INV_X1    g0110(.A(G169), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n303), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n310), .A2(G179), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n302), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n251), .B1(new_n284), .B2(new_n314), .ZN(new_n315));
  XNOR2_X1  g0115(.A(KEYINPUT3), .B(G33), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n267), .B1(new_n316), .B2(G20), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n265), .A2(KEYINPUT7), .A3(new_n219), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n203), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n276), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n278), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n283), .A2(new_n321), .A3(new_n258), .ZN(new_n322));
  INV_X1    g0122(.A(new_n261), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(G169), .B1(new_n299), .B2(new_n301), .ZN(new_n325));
  OAI22_X1  g0125(.A1(new_n325), .A2(new_n303), .B1(G179), .B2(new_n310), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n324), .A2(new_n326), .A3(KEYINPUT18), .A4(new_n302), .ZN(new_n327));
  AND2_X1   g0127(.A1(new_n315), .A2(new_n327), .ZN(new_n328));
  AND3_X1   g0128(.A1(new_n287), .A2(G232), .A3(new_n296), .ZN(new_n329));
  INV_X1    g0129(.A(G190), .ZN(new_n330));
  NOR4_X1   g0130(.A1(new_n295), .A2(new_n329), .A3(new_n330), .A4(new_n298), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n331), .B1(G200), .B2(new_n310), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n332), .A2(new_n322), .A3(new_n323), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT75), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n334), .A2(KEYINPUT17), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  XNOR2_X1  g0136(.A(KEYINPUT75), .B(KEYINPUT17), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n284), .A2(new_n332), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n328), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT13), .ZN(new_n341));
  INV_X1    g0141(.A(G1698), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n289), .A2(new_n342), .ZN(new_n343));
  OAI221_X1 g0143(.A(new_n343), .B1(G232), .B2(new_n342), .C1(new_n263), .C2(new_n264), .ZN(new_n344));
  NAND2_X1  g0144(.A1(G33), .A2(G97), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n287), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n298), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n287), .A2(new_n296), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(KEYINPUT71), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT71), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n287), .A2(new_n351), .A3(new_n296), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n350), .A2(G238), .A3(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n341), .B1(new_n348), .B2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n348), .A2(new_n341), .A3(new_n353), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n355), .A2(KEYINPUT72), .A3(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT72), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n354), .A2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(G190), .B1(new_n358), .B2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n356), .ZN(new_n363));
  OAI21_X1  g0163(.A(G200), .B1(new_n363), .B2(new_n354), .ZN(new_n364));
  OAI22_X1  g0164(.A1(new_n271), .A2(new_n201), .B1(new_n219), .B2(G68), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n219), .A2(G33), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n366), .A2(new_n212), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n258), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  XOR2_X1   g0168(.A(new_n368), .B(KEYINPUT11), .Z(new_n369));
  NOR2_X1   g0169(.A1(new_n260), .A2(new_n203), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n254), .A2(G68), .ZN(new_n371));
  XNOR2_X1  g0171(.A(new_n371), .B(KEYINPUT12), .ZN(new_n372));
  NOR3_X1   g0172(.A1(new_n369), .A2(new_n370), .A3(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n362), .A2(new_n364), .A3(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n373), .ZN(new_n375));
  OAI21_X1  g0175(.A(G169), .B1(new_n363), .B2(new_n354), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(KEYINPUT14), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT14), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n378), .B(G169), .C1(new_n363), .C2(new_n354), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n300), .B1(new_n357), .B2(new_n360), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n375), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n253), .A2(new_n270), .B1(G20), .B2(G77), .ZN(new_n383));
  XOR2_X1   g0183(.A(KEYINPUT15), .B(G87), .Z(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n383), .B1(new_n366), .B2(new_n385), .ZN(new_n386));
  AOI22_X1  g0186(.A1(new_n386), .A2(new_n258), .B1(new_n212), .B2(new_n255), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n387), .B1(new_n212), .B2(new_n260), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n316), .A2(G232), .A3(new_n342), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n316), .A2(G238), .A3(G1698), .ZN(new_n390));
  INV_X1    g0190(.A(G107), .ZN(new_n391));
  OAI211_X1 g0191(.A(new_n389), .B(new_n390), .C1(new_n391), .C2(new_n316), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n347), .ZN(new_n393));
  INV_X1    g0193(.A(new_n349), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(G244), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n393), .A2(new_n304), .A3(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT68), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n393), .A2(KEYINPUT68), .A3(new_n304), .A4(new_n395), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n388), .B1(new_n400), .B2(G190), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n398), .A2(G200), .A3(new_n399), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n340), .A2(new_n374), .A3(new_n382), .A4(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n204), .A2(G20), .ZN(new_n405));
  INV_X1    g0205(.A(G150), .ZN(new_n406));
  OAI221_X1 g0206(.A(new_n405), .B1(new_n406), .B2(new_n271), .C1(new_n252), .C2(new_n366), .ZN(new_n407));
  AOI22_X1  g0207(.A1(new_n407), .A2(new_n258), .B1(new_n201), .B2(new_n255), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n259), .A2(G50), .ZN(new_n409));
  AOI21_X1  g0209(.A(KEYINPUT9), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  OAI211_X1 g0210(.A(G222), .B(new_n342), .C1(new_n263), .C2(new_n264), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT67), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n316), .A2(KEYINPUT67), .A3(G222), .A4(new_n342), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n265), .A2(G77), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n316), .A2(G223), .A3(G1698), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n413), .A2(new_n414), .A3(new_n415), .A4(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(new_n347), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n394), .A2(G226), .ZN(new_n419));
  AND3_X1   g0219(.A1(new_n418), .A2(new_n304), .A3(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n410), .B1(new_n420), .B2(G190), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n407), .A2(new_n258), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n255), .A2(new_n201), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n422), .A2(new_n409), .A3(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT9), .ZN(new_n425));
  OAI21_X1  g0225(.A(KEYINPUT69), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT69), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n408), .A2(new_n427), .A3(KEYINPUT9), .A4(new_n409), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n418), .A2(new_n304), .A3(new_n419), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n430), .A2(KEYINPUT70), .A3(G200), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(KEYINPUT70), .B1(new_n430), .B2(G200), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n421), .B(new_n429), .C1(new_n432), .C2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(KEYINPUT10), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT70), .ZN(new_n436));
  INV_X1    g0236(.A(G200), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n436), .B1(new_n420), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n431), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT10), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n439), .A2(new_n440), .A3(new_n429), .A4(new_n421), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n435), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n420), .A2(new_n300), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n443), .B(new_n424), .C1(G169), .C2(new_n420), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n400), .A2(new_n300), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n398), .A2(new_n311), .A3(new_n399), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n445), .A2(new_n388), .A3(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n442), .A2(new_n444), .A3(new_n447), .ZN(new_n448));
  OAI211_X1 g0248(.A(G257), .B(new_n342), .C1(new_n263), .C2(new_n264), .ZN(new_n449));
  OAI211_X1 g0249(.A(G264), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n306), .A2(G303), .A3(new_n307), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(new_n347), .ZN(new_n453));
  INV_X1    g0253(.A(G45), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n454), .A2(G1), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(G274), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n286), .A2(KEYINPUT5), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT5), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(G41), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n456), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n455), .A2(new_n457), .A3(new_n459), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n463), .A2(G270), .A3(new_n287), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(KEYINPUT79), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT79), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n463), .A2(new_n466), .A3(G270), .A4(new_n287), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n453), .A2(new_n462), .A3(new_n465), .A4(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n468), .A2(KEYINPUT21), .A3(G169), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n461), .B1(new_n452), .B2(new_n347), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n470), .A2(G179), .A3(new_n465), .A4(new_n467), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(G116), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n255), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n218), .A2(G33), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n262), .A2(G116), .A3(new_n254), .A4(new_n475), .ZN(new_n476));
  AOI22_X1  g0276(.A1(new_n257), .A2(new_n228), .B1(G20), .B2(new_n473), .ZN(new_n477));
  NAND2_X1  g0277(.A1(G33), .A2(G283), .ZN(new_n478));
  INV_X1    g0278(.A(G97), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n478), .B(new_n219), .C1(G33), .C2(new_n479), .ZN(new_n480));
  AND3_X1   g0280(.A1(new_n477), .A2(KEYINPUT20), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(KEYINPUT20), .B1(new_n477), .B2(new_n480), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n474), .B(new_n476), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n472), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n468), .A2(G169), .A3(new_n483), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT21), .ZN(new_n486));
  AND3_X1   g0286(.A1(new_n485), .A2(KEYINPUT80), .A3(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(KEYINPUT80), .B1(new_n485), .B2(new_n486), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n484), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n468), .A2(G200), .ZN(new_n490));
  INV_X1    g0290(.A(new_n483), .ZN(new_n491));
  AOI21_X1  g0291(.A(KEYINPUT81), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT81), .ZN(new_n493));
  AOI211_X1 g0293(.A(new_n493), .B(new_n483), .C1(new_n468), .C2(G200), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n468), .A2(new_n330), .ZN(new_n495));
  NOR3_X1   g0295(.A1(new_n492), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n489), .A2(new_n496), .ZN(new_n497));
  AND3_X1   g0297(.A1(new_n262), .A2(new_n254), .A3(new_n475), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(G107), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT85), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n500), .B(KEYINPUT25), .C1(new_n254), .C2(G107), .ZN(new_n501));
  OR2_X1    g0301(.A1(new_n500), .A2(KEYINPUT25), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n500), .A2(KEYINPUT25), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n255), .A2(new_n502), .A3(new_n391), .A4(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n499), .A2(new_n501), .A3(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT84), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT82), .ZN(new_n508));
  NAND2_X1  g0308(.A1(G33), .A2(G116), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n508), .B1(new_n509), .B2(G20), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n219), .A2(KEYINPUT82), .A3(G33), .A4(G116), .ZN(new_n511));
  AND2_X1   g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  OR2_X1    g0313(.A1(KEYINPUT83), .A2(KEYINPUT23), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n391), .A2(G20), .ZN(new_n515));
  NAND2_X1  g0315(.A1(KEYINPUT83), .A2(KEYINPUT23), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n517), .B1(new_n515), .B2(new_n516), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT22), .ZN(new_n519));
  AOI21_X1  g0319(.A(G20), .B1(new_n306), .B2(new_n307), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n519), .B1(new_n520), .B2(G87), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n219), .B(G87), .C1(new_n263), .C2(new_n264), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n522), .A2(KEYINPUT22), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n513), .B(new_n518), .C1(new_n521), .C2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(KEYINPUT24), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n522), .A2(KEYINPUT22), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n316), .A2(new_n519), .A3(new_n219), .A4(G87), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n512), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT24), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n528), .A2(new_n529), .A3(new_n518), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n525), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n507), .B1(new_n531), .B2(new_n258), .ZN(new_n532));
  AOI211_X1 g0332(.A(KEYINPUT84), .B(new_n262), .C1(new_n525), .C2(new_n530), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n506), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OAI211_X1 g0334(.A(G257), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(KEYINPUT86), .ZN(new_n536));
  XOR2_X1   g0336(.A(KEYINPUT87), .B(G294), .Z(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(G33), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT86), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n316), .A2(new_n539), .A3(G257), .A4(G1698), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n316), .A2(G250), .A3(new_n342), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n536), .A2(new_n538), .A3(new_n540), .A4(new_n541), .ZN(new_n542));
  AND2_X1   g0342(.A1(new_n463), .A2(new_n287), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n542), .A2(new_n347), .B1(G264), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n462), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n546), .A2(G169), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n546), .A2(new_n300), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n534), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n463), .A2(G257), .A3(new_n287), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT76), .ZN(new_n552));
  XNOR2_X1  g0352(.A(new_n551), .B(new_n552), .ZN(new_n553));
  OAI211_X1 g0353(.A(G244), .B(new_n342), .C1(new_n263), .C2(new_n264), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT4), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n316), .A2(KEYINPUT4), .A3(G244), .A4(new_n342), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n316), .A2(G250), .A3(G1698), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n556), .A2(new_n557), .A3(new_n558), .A4(new_n478), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n347), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n553), .A2(new_n560), .A3(new_n462), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n311), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n391), .A2(KEYINPUT6), .A3(G97), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT6), .ZN(new_n565));
  XNOR2_X1  g0365(.A(G97), .B(G107), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  OAI22_X1  g0367(.A1(new_n567), .A2(new_n219), .B1(new_n212), .B2(new_n271), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n391), .B1(new_n317), .B2(new_n318), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n258), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n262), .A2(new_n254), .A3(new_n475), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n571), .A2(new_n479), .ZN(new_n572));
  INV_X1    g0372(.A(new_n572), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n570), .B(new_n573), .C1(G97), .C2(new_n254), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n461), .B1(new_n559), .B2(new_n347), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n575), .A2(new_n300), .A3(new_n553), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n562), .A2(new_n574), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n561), .A2(G200), .ZN(new_n578));
  OAI21_X1  g0378(.A(G107), .B1(new_n266), .B2(new_n268), .ZN(new_n579));
  AND2_X1   g0379(.A1(G97), .A2(G107), .ZN(new_n580));
  NOR2_X1   g0380(.A1(G97), .A2(G107), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n565), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n563), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n583), .A2(G20), .B1(G77), .B2(new_n270), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n262), .B1(new_n579), .B2(new_n584), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n254), .A2(G97), .ZN(new_n586));
  NOR3_X1   g0386(.A1(new_n585), .A2(new_n572), .A3(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n575), .A2(G190), .A3(new_n553), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n578), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n498), .A2(new_n384), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n384), .A2(new_n254), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT19), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n219), .B1(new_n345), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n581), .A2(new_n292), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n219), .A2(G33), .A3(G97), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n594), .A2(new_n595), .B1(new_n593), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n316), .A2(new_n219), .A3(G68), .ZN(new_n598));
  AND2_X1   g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n590), .B(new_n592), .C1(new_n599), .C2(new_n262), .ZN(new_n600));
  OR2_X1    g0400(.A1(G238), .A2(G1698), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n213), .A2(G1698), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n601), .B(new_n602), .C1(new_n263), .C2(new_n264), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n509), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n347), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n218), .A2(G45), .ZN(new_n606));
  AND2_X1   g0406(.A1(G33), .A2(G41), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n606), .B(G250), .C1(new_n607), .C2(new_n228), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n608), .A2(KEYINPUT77), .A3(new_n456), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(KEYINPUT77), .B1(new_n608), .B2(new_n456), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n605), .B(new_n300), .C1(new_n610), .C2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n608), .A2(new_n456), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT77), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n615), .A2(new_n609), .B1(new_n347), .B2(new_n604), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n600), .B(new_n612), .C1(G169), .C2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT78), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n616), .A2(new_n618), .A3(G190), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n605), .B(G190), .C1(new_n610), .C2(new_n611), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(KEYINPUT78), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n605), .B1(new_n610), .B2(new_n611), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(G200), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n262), .B1(new_n597), .B2(new_n598), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n571), .A2(new_n292), .ZN(new_n625));
  NOR3_X1   g0425(.A1(new_n624), .A2(new_n625), .A3(new_n591), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n619), .A2(new_n621), .A3(new_n623), .A4(new_n626), .ZN(new_n627));
  AND4_X1   g0427(.A1(new_n577), .A2(new_n589), .A3(new_n617), .A4(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n526), .A2(new_n527), .ZN(new_n629));
  AND4_X1   g0429(.A1(new_n529), .A2(new_n629), .A3(new_n513), .A4(new_n518), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n529), .B1(new_n528), .B2(new_n518), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n258), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(KEYINPUT84), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n531), .A2(new_n507), .A3(new_n258), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n546), .A2(G190), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n437), .B1(new_n544), .B2(new_n462), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n635), .A2(new_n636), .A3(new_n506), .A4(new_n638), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n497), .A2(new_n550), .A3(new_n628), .A4(new_n639), .ZN(new_n640));
  NOR3_X1   g0440(.A1(new_n404), .A2(new_n448), .A3(new_n640), .ZN(G372));
  NOR2_X1   g0441(.A1(new_n404), .A2(new_n448), .ZN(new_n642));
  AND3_X1   g0442(.A1(new_n562), .A2(new_n574), .A3(new_n576), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT26), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n623), .A2(new_n626), .A3(new_n620), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n617), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n643), .A2(new_n644), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n627), .A2(new_n617), .ZN(new_n648));
  OAI21_X1  g0448(.A(KEYINPUT26), .B1(new_n648), .B2(new_n577), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n547), .B1(new_n635), .B2(new_n506), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n489), .B1(new_n651), .B2(new_n549), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n646), .A2(new_n577), .A3(new_n589), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(new_n639), .ZN(new_n654));
  OAI211_X1 g0454(.A(new_n617), .B(new_n650), .C1(new_n652), .C2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n642), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g0456(.A(new_n656), .B(KEYINPUT88), .Z(new_n657));
  INV_X1    g0457(.A(new_n444), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n315), .A2(new_n327), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n382), .A2(new_n447), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(new_n374), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n659), .B1(new_n661), .B2(new_n339), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n658), .B1(new_n662), .B2(new_n442), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n657), .A2(new_n663), .ZN(G369));
  INV_X1    g0464(.A(G13), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n665), .A2(G20), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  OR3_X1    g0467(.A1(new_n667), .A2(KEYINPUT27), .A3(G1), .ZN(new_n668));
  OAI21_X1  g0468(.A(KEYINPUT27), .B1(new_n667), .B2(G1), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n668), .A2(G213), .A3(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(G343), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n534), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(new_n639), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(new_n550), .ZN(new_n675));
  INV_X1    g0475(.A(new_n672), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n651), .A2(new_n549), .A3(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n489), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n678), .A2(new_n672), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n675), .A2(new_n677), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(new_n677), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(KEYINPUT89), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT89), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n680), .A2(new_n683), .A3(new_n677), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(G330), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n497), .B1(new_n491), .B2(new_n676), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n489), .A2(new_n483), .A3(new_n672), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n686), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n675), .A2(new_n677), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n685), .A2(new_n693), .ZN(G399));
  NAND2_X1  g0494(.A1(new_n225), .A2(new_n286), .ZN(new_n695));
  XNOR2_X1  g0495(.A(new_n695), .B(KEYINPUT90), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n595), .A2(G116), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(G1), .A3(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n699), .B1(new_n231), .B2(new_n697), .ZN(new_n700));
  XNOR2_X1  g0500(.A(new_n700), .B(KEYINPUT28), .ZN(new_n701));
  NOR3_X1   g0501(.A1(new_n648), .A2(new_n577), .A3(KEYINPUT26), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n644), .B1(new_n643), .B2(new_n646), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  OAI211_X1 g0504(.A(new_n617), .B(new_n704), .C1(new_n652), .C2(new_n654), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n705), .A2(KEYINPUT29), .A3(new_n676), .ZN(new_n706));
  INV_X1    g0506(.A(new_n617), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n646), .A2(new_n577), .A3(new_n589), .ZN(new_n708));
  AOI211_X1 g0508(.A(new_n505), .B(new_n637), .C1(new_n633), .C2(new_n634), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n708), .B1(new_n709), .B2(new_n636), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n550), .A2(new_n678), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n707), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n672), .B1(new_n712), .B2(new_n650), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n706), .B1(new_n713), .B2(KEYINPUT29), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n577), .A2(new_n589), .A3(new_n617), .A4(new_n627), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n715), .B1(new_n709), .B2(new_n636), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n716), .A2(new_n550), .A3(new_n497), .A4(new_n676), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT30), .ZN(new_n718));
  INV_X1    g0518(.A(new_n468), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n719), .A2(G179), .A3(new_n575), .A4(new_n553), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n544), .A2(new_n616), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n718), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n561), .A2(new_n471), .ZN(new_n723));
  INV_X1    g0523(.A(new_n721), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n723), .A2(new_n724), .A3(KEYINPUT30), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n616), .B1(new_n575), .B2(new_n553), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n726), .A2(new_n545), .A3(new_n300), .A4(new_n468), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n722), .A2(new_n725), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(new_n672), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(KEYINPUT31), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT31), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n728), .A2(new_n731), .A3(new_n672), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n686), .B1(new_n717), .B2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n714), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n701), .B1(new_n737), .B2(G1), .ZN(G364));
  OR2_X1    g0538(.A1(new_n311), .A2(KEYINPUT92), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n311), .A2(KEYINPUT92), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n739), .A2(G20), .A3(new_n740), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n741), .A2(G1), .A3(G13), .ZN(new_n742));
  XNOR2_X1  g0542(.A(new_n742), .B(KEYINPUT93), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n219), .A2(G190), .ZN(new_n744));
  NOR2_X1   g0544(.A1(G179), .A2(G200), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  XNOR2_X1  g0547(.A(KEYINPUT94), .B(G159), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  XOR2_X1   g0549(.A(new_n749), .B(KEYINPUT95), .Z(new_n750));
  AND2_X1   g0550(.A1(new_n750), .A2(KEYINPUT32), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(KEYINPUT32), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n300), .A2(new_n437), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(new_n744), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(new_n203), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n219), .B1(new_n745), .B2(G190), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(new_n479), .ZN(new_n757));
  NOR4_X1   g0557(.A1(new_n751), .A2(new_n752), .A3(new_n755), .A4(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n437), .A2(G179), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(new_n744), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(G107), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n219), .A2(new_n330), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(new_n759), .ZN(new_n764));
  OAI211_X1 g0564(.A(new_n762), .B(new_n316), .C1(new_n292), .C2(new_n764), .ZN(new_n765));
  XNOR2_X1  g0565(.A(new_n765), .B(KEYINPUT96), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n744), .A2(G179), .A3(new_n437), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n766), .B1(G77), .B2(new_n768), .ZN(new_n769));
  AND2_X1   g0569(.A1(new_n763), .A2(new_n753), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G50), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n763), .A2(G179), .A3(new_n437), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G58), .ZN(new_n774));
  NAND4_X1  g0574(.A1(new_n758), .A2(new_n769), .A3(new_n771), .A4(new_n774), .ZN(new_n775));
  AOI22_X1  g0575(.A1(new_n773), .A2(G322), .B1(new_n747), .B2(G329), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n770), .A2(G326), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n776), .A2(new_n265), .A3(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n778), .B1(G283), .B2(new_n761), .ZN(new_n779));
  INV_X1    g0579(.A(new_n764), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(G303), .ZN(new_n781));
  INV_X1    g0581(.A(new_n756), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(new_n537), .ZN(new_n783));
  INV_X1    g0583(.A(new_n754), .ZN(new_n784));
  XNOR2_X1  g0584(.A(KEYINPUT33), .B(G317), .ZN(new_n785));
  AOI22_X1  g0585(.A1(G311), .A2(new_n768), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NAND4_X1  g0586(.A1(new_n779), .A2(new_n781), .A3(new_n783), .A4(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n743), .B1(new_n775), .B2(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n218), .B1(new_n666), .B2(G45), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n697), .A2(new_n789), .ZN(new_n790));
  XOR2_X1   g0590(.A(new_n790), .B(KEYINPUT91), .Z(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n743), .ZN(new_n793));
  NOR3_X1   g0593(.A1(G13), .A2(G20), .A3(G33), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n232), .A2(new_n454), .ZN(new_n796));
  INV_X1    g0596(.A(new_n225), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(new_n316), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n796), .B(new_n798), .C1(new_n245), .C2(new_n454), .ZN(new_n799));
  INV_X1    g0599(.A(G355), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n225), .A2(new_n316), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n799), .B1(G116), .B2(new_n225), .C1(new_n800), .C2(new_n801), .ZN(new_n802));
  AOI211_X1 g0602(.A(new_n788), .B(new_n792), .C1(new_n795), .C2(new_n802), .ZN(new_n803));
  XOR2_X1   g0603(.A(new_n794), .B(KEYINPUT97), .Z(new_n804));
  NAND3_X1  g0604(.A1(new_n687), .A2(new_n688), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n687), .A2(new_n686), .A3(new_n688), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n690), .A2(new_n792), .A3(new_n807), .ZN(new_n808));
  AND2_X1   g0608(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(G396));
  NAND4_X1  g0610(.A1(new_n445), .A2(new_n388), .A3(new_n446), .A4(new_n676), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n401), .A2(new_n402), .B1(new_n388), .B2(new_n672), .ZN(new_n812));
  AND3_X1   g0612(.A1(new_n445), .A2(new_n388), .A3(new_n446), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n811), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n713), .B(new_n814), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n815), .B(new_n735), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(new_n792), .ZN(new_n817));
  NOR2_X1   g0617(.A1(G13), .A2(G33), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n792), .B1(new_n818), .B2(new_n814), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n793), .A2(new_n818), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(new_n212), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n764), .A2(new_n391), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n757), .B(new_n822), .C1(G116), .C2(new_n768), .ZN(new_n823));
  INV_X1    g0623(.A(G311), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n746), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n760), .A2(new_n292), .ZN(new_n826));
  AOI211_X1 g0626(.A(new_n825), .B(new_n826), .C1(G303), .C2(new_n770), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n784), .A2(G283), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n316), .B1(new_n773), .B2(G294), .ZN(new_n829));
  NAND4_X1  g0629(.A1(new_n823), .A2(new_n827), .A3(new_n828), .A4(new_n829), .ZN(new_n830));
  AOI22_X1  g0630(.A1(G68), .A2(new_n761), .B1(new_n747), .B2(G132), .ZN(new_n831));
  OAI211_X1 g0631(.A(new_n831), .B(new_n316), .C1(new_n201), .C2(new_n764), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n832), .B1(G58), .B2(new_n782), .ZN(new_n833));
  XNOR2_X1  g0633(.A(new_n833), .B(KEYINPUT98), .ZN(new_n834));
  AOI22_X1  g0634(.A1(G143), .A2(new_n773), .B1(new_n768), .B2(new_n748), .ZN(new_n835));
  INV_X1    g0635(.A(G137), .ZN(new_n836));
  INV_X1    g0636(.A(new_n770), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n835), .B1(new_n836), .B2(new_n837), .C1(new_n406), .C2(new_n754), .ZN(new_n838));
  XOR2_X1   g0638(.A(new_n838), .B(KEYINPUT34), .Z(new_n839));
  OAI21_X1  g0639(.A(new_n830), .B1(new_n834), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(new_n793), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n819), .A2(new_n821), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n817), .A2(new_n842), .ZN(G384));
  NAND2_X1  g0643(.A1(new_n375), .A2(new_n672), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n374), .A2(new_n382), .A3(new_n844), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n375), .B(new_n672), .C1(new_n380), .C2(new_n381), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n814), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n655), .A2(new_n676), .A3(new_n849), .ZN(new_n850));
  XOR2_X1   g0650(.A(new_n811), .B(KEYINPUT101), .Z(new_n851));
  AOI21_X1  g0651(.A(new_n848), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n670), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n269), .A2(new_n281), .A3(new_n282), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT102), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n854), .A2(new_n855), .A3(new_n278), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n855), .A2(new_n278), .ZN(new_n857));
  NAND4_X1  g0657(.A1(new_n269), .A2(new_n281), .A3(new_n282), .A4(new_n857), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n856), .A2(new_n258), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(new_n323), .ZN(new_n860));
  OAI211_X1 g0660(.A(new_n853), .B(new_n860), .C1(new_n328), .C2(new_n339), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT103), .ZN(new_n862));
  NAND4_X1  g0662(.A1(new_n324), .A2(new_n326), .A3(new_n862), .A4(new_n302), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT37), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n324), .A2(new_n853), .ZN(new_n865));
  NAND4_X1  g0665(.A1(new_n863), .A2(new_n864), .A3(new_n333), .A4(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(KEYINPUT103), .B1(new_n284), .B2(new_n314), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n314), .A2(new_n670), .ZN(new_n869));
  AOI22_X1  g0669(.A1(new_n860), .A2(new_n869), .B1(new_n284), .B2(new_n332), .ZN(new_n870));
  OAI22_X1  g0670(.A1(new_n866), .A2(new_n868), .B1(new_n870), .B2(new_n864), .ZN(new_n871));
  AND3_X1   g0671(.A1(new_n861), .A2(KEYINPUT38), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(KEYINPUT38), .B1(new_n861), .B2(new_n871), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n852), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n861), .A2(new_n871), .A3(KEYINPUT38), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT104), .ZN(new_n876));
  INV_X1    g0676(.A(new_n335), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n877), .B1(new_n284), .B2(new_n332), .ZN(new_n878));
  AND4_X1   g0678(.A1(new_n322), .A2(new_n332), .A3(new_n323), .A4(new_n337), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n876), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n336), .A2(new_n338), .A3(KEYINPUT104), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n880), .A2(new_n659), .A3(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n865), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n865), .A2(new_n333), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n885), .A2(new_n864), .A3(new_n867), .A4(new_n863), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n284), .A2(new_n314), .ZN(new_n887));
  OAI21_X1  g0687(.A(KEYINPUT37), .B1(new_n884), .B2(new_n887), .ZN(new_n888));
  AOI22_X1  g0688(.A1(new_n882), .A2(new_n883), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n875), .B1(new_n889), .B2(KEYINPUT38), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT39), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  OR2_X1    g0692(.A1(new_n382), .A2(new_n672), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n873), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n895), .A2(KEYINPUT39), .A3(new_n875), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n892), .A2(new_n894), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n328), .A2(new_n670), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n874), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n642), .B(new_n706), .C1(new_n713), .C2(KEYINPUT29), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n663), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n899), .B(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT106), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n731), .B1(new_n728), .B2(new_n672), .ZN(new_n905));
  AND3_X1   g0705(.A1(new_n728), .A2(new_n731), .A3(new_n672), .ZN(new_n906));
  OAI22_X1  g0706(.A1(new_n640), .A2(new_n672), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n642), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n908), .B(KEYINPUT105), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT40), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT38), .ZN(new_n911));
  AND2_X1   g0711(.A1(new_n882), .A2(new_n883), .ZN(new_n912));
  AND2_X1   g0712(.A1(new_n886), .A2(new_n888), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n911), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n910), .B1(new_n914), .B2(new_n875), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n814), .B1(new_n845), .B2(new_n846), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(new_n907), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n907), .B(new_n916), .C1(new_n872), .C2(new_n873), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n915), .A2(new_n918), .B1(new_n919), .B2(new_n910), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n909), .B(new_n920), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n921), .A2(new_n686), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n904), .A2(new_n922), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n902), .B(KEYINPUT106), .ZN(new_n924));
  OAI221_X1 g0724(.A(new_n923), .B1(new_n218), .B2(new_n666), .C1(new_n924), .C2(new_n922), .ZN(new_n925));
  OAI211_X1 g0725(.A(G116), .B(new_n229), .C1(new_n583), .C2(KEYINPUT35), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n926), .B(KEYINPUT99), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT35), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n927), .B1(new_n928), .B2(new_n567), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n929), .B(KEYINPUT36), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n274), .A2(G77), .ZN(new_n931));
  OAI22_X1  g0731(.A1(new_n231), .A2(new_n931), .B1(G50), .B2(new_n203), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n932), .A2(G1), .A3(new_n665), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n930), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n934), .B(KEYINPUT100), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n925), .A2(new_n935), .ZN(G367));
  INV_X1    g0736(.A(new_n798), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n795), .B1(new_n240), .B2(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n938), .B1(new_n797), .B2(new_n384), .ZN(new_n939));
  INV_X1    g0739(.A(new_n804), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n646), .B1(new_n626), .B2(new_n676), .ZN(new_n941));
  OR3_X1    g0741(.A1(new_n617), .A2(new_n626), .A3(new_n676), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n791), .B1(new_n940), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n768), .A2(G50), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n784), .A2(new_n748), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n770), .A2(G143), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n782), .A2(G68), .ZN(new_n948));
  NAND4_X1  g0748(.A1(new_n945), .A2(new_n946), .A3(new_n947), .A4(new_n948), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n772), .A2(new_n406), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n316), .B1(new_n746), .B2(new_n836), .ZN(new_n951));
  OAI22_X1  g0751(.A1(new_n764), .A2(new_n202), .B1(new_n760), .B2(new_n212), .ZN(new_n952));
  NOR4_X1   g0752(.A1(new_n949), .A2(new_n950), .A3(new_n951), .A4(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n780), .A2(G116), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT46), .ZN(new_n955));
  AOI22_X1  g0755(.A1(new_n954), .A2(new_n955), .B1(G311), .B2(new_n770), .ZN(new_n956));
  AOI22_X1  g0756(.A1(G303), .A2(new_n773), .B1(new_n768), .B2(G283), .ZN(new_n957));
  OAI211_X1 g0757(.A(new_n956), .B(new_n957), .C1(new_n955), .C2(new_n954), .ZN(new_n958));
  INV_X1    g0758(.A(new_n537), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n959), .A2(new_n754), .B1(new_n479), .B2(new_n760), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n265), .B1(new_n756), .B2(new_n391), .ZN(new_n961));
  NOR3_X1   g0761(.A1(new_n958), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n747), .A2(G317), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n953), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n964), .B(KEYINPUT47), .Z(new_n965));
  AOI211_X1 g0765(.A(new_n939), .B(new_n944), .C1(new_n793), .C2(new_n965), .ZN(new_n966));
  OAI211_X1 g0766(.A(new_n577), .B(new_n589), .C1(new_n587), .C2(new_n676), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n643), .A2(new_n672), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n685), .A2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT45), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n685), .A2(KEYINPUT45), .A3(new_n969), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT44), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n685), .B2(new_n969), .ZN(new_n976));
  INV_X1    g0776(.A(new_n969), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n682), .A2(KEYINPUT44), .A3(new_n684), .A4(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n974), .A2(new_n979), .A3(new_n693), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n689), .A2(new_n679), .ZN(new_n981));
  INV_X1    g0781(.A(new_n691), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n981), .B(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n736), .B1(new_n980), .B2(new_n983), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n696), .B(KEYINPUT41), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n789), .B1(new_n984), .B2(new_n986), .ZN(new_n987));
  OR2_X1    g0787(.A1(new_n680), .A2(new_n967), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n988), .A2(KEYINPUT42), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n577), .B1(new_n550), .B2(new_n967), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(new_n676), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n988), .A2(KEYINPUT42), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n989), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n943), .A2(KEYINPUT43), .ZN(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n943), .A2(KEYINPUT43), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n993), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n995), .B1(new_n993), .B2(new_n996), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n998), .A2(new_n999), .B1(new_n693), .B2(new_n977), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n999), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n693), .A2(new_n977), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n1001), .A2(new_n1002), .A3(new_n997), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1000), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n966), .B1(new_n987), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(G387));
  OAI21_X1  g0807(.A(KEYINPUT108), .B1(new_n737), .B2(new_n983), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n737), .A2(new_n983), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n981), .B(new_n691), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT108), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1010), .A2(new_n736), .A3(new_n1011), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1008), .A2(new_n696), .A3(new_n1009), .A4(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n789), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n983), .A2(new_n1014), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n784), .A2(G311), .B1(new_n770), .B2(G322), .ZN(new_n1016));
  INV_X1    g0816(.A(G303), .ZN(new_n1017));
  INV_X1    g0817(.A(G317), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n1016), .B1(new_n1017), .B2(new_n767), .C1(new_n1018), .C2(new_n772), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT48), .ZN(new_n1020));
  INV_X1    g0820(.A(G283), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n1020), .B1(new_n1021), .B2(new_n756), .C1(new_n959), .C2(new_n764), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT49), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(G116), .A2(new_n761), .B1(new_n747), .B2(G326), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1023), .A2(new_n265), .A3(new_n1024), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n837), .A2(new_n272), .B1(new_n201), .B2(new_n772), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(G97), .B2(new_n761), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n764), .A2(new_n212), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n767), .A2(new_n203), .B1(new_n746), .B2(new_n406), .ZN(new_n1029));
  AOI211_X1 g0829(.A(new_n1028), .B(new_n1029), .C1(new_n384), .C2(new_n782), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n784), .A2(new_n253), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1027), .A2(new_n1030), .A3(new_n316), .A4(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n743), .B1(new_n1025), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n253), .A2(new_n201), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT107), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT50), .ZN(new_n1036));
  AOI21_X1  g0836(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1036), .A2(new_n698), .A3(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n798), .B1(new_n237), .B2(new_n454), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(new_n698), .B2(new_n801), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1041), .B1(G107), .B2(new_n225), .ZN(new_n1042));
  AOI211_X1 g0842(.A(new_n792), .B(new_n1033), .C1(new_n795), .C2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(new_n982), .B2(new_n940), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1013), .A2(new_n1015), .A3(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(KEYINPUT109), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT109), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n1013), .A2(new_n1047), .A3(new_n1015), .A4(new_n1044), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1046), .A2(new_n1048), .ZN(G393));
  AOI22_X1  g0849(.A1(new_n972), .A2(new_n973), .B1(new_n976), .B2(new_n978), .ZN(new_n1050));
  OR2_X1    g0850(.A1(new_n1050), .A2(new_n693), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1051), .A2(KEYINPUT110), .A3(new_n980), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT110), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n980), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n1050), .A2(new_n693), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1053), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1052), .A2(new_n1056), .A3(new_n1014), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1009), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1009), .B1(new_n1050), .B2(new_n693), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1059), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1058), .A2(new_n696), .A3(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n792), .B1(new_n977), .B2(new_n794), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n265), .B(new_n826), .C1(G50), .C2(new_n784), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n782), .A2(G77), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n747), .A2(G143), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n253), .A2(new_n768), .B1(new_n780), .B2(G68), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n1063), .A2(new_n1064), .A3(new_n1065), .A4(new_n1066), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n773), .A2(G159), .B1(new_n770), .B2(G150), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(KEYINPUT111), .B(KEYINPUT51), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1068), .B(new_n1069), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n1067), .A2(new_n1070), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT112), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n837), .A2(new_n1018), .B1(new_n824), .B2(new_n772), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT52), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n764), .A2(new_n1021), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n754), .A2(new_n1017), .B1(new_n756), .B2(new_n473), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n1075), .B(new_n1076), .C1(G322), .C2(new_n747), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n316), .B1(new_n768), .B2(G294), .ZN(new_n1078));
  AND4_X1   g0878(.A1(new_n762), .A2(new_n1074), .A3(new_n1077), .A4(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n793), .B1(new_n1072), .B2(new_n1079), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n795), .B1(new_n479), .B2(new_n225), .C1(new_n249), .C2(new_n937), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1062), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1057), .A2(new_n1061), .A3(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT113), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n1057), .A2(new_n1061), .A3(KEYINPUT113), .A4(new_n1082), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1085), .A2(new_n1086), .ZN(G390));
  NAND2_X1  g0887(.A1(new_n892), .A2(new_n896), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n818), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n756), .A2(new_n272), .ZN(new_n1090));
  INV_X1    g0890(.A(G125), .ZN(new_n1091));
  OAI221_X1 g0891(.A(new_n316), .B1(new_n746), .B2(new_n1091), .C1(new_n201), .C2(new_n760), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT114), .ZN(new_n1093));
  XOR2_X1   g0893(.A(KEYINPUT54), .B(G143), .Z(new_n1094));
  AOI211_X1 g0894(.A(new_n1090), .B(new_n1093), .C1(new_n768), .C2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n770), .A2(G128), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n773), .A2(G132), .B1(new_n784), .B2(G137), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n764), .A2(new_n406), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n1098), .B(KEYINPUT53), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n1095), .A2(new_n1096), .A3(new_n1097), .A4(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(G294), .ZN(new_n1101));
  OAI221_X1 g0901(.A(new_n1064), .B1(new_n1101), .B2(new_n746), .C1(new_n837), .C2(new_n1021), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(G68), .B2(new_n761), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n292), .A2(new_n764), .B1(new_n754), .B2(new_n391), .ZN(new_n1104));
  AOI211_X1 g0904(.A(new_n316), .B(new_n1104), .C1(G97), .C2(new_n768), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n1103), .B(new_n1105), .C1(new_n473), .C2(new_n772), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n743), .B1(new_n1100), .B2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(new_n252), .B2(new_n820), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1089), .A2(new_n791), .A3(new_n1108), .ZN(new_n1109));
  AND3_X1   g0909(.A1(new_n916), .A2(new_n907), .A3(G330), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n850), .A2(new_n851), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(new_n847), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n1112), .A2(new_n893), .B1(new_n892), .B2(new_n896), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n890), .A2(new_n893), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n705), .A2(new_n676), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n812), .A2(new_n813), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n811), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1114), .B1(new_n1117), .B2(new_n847), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1110), .B1(new_n1113), .B2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1088), .B1(new_n894), .B2(new_n852), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n811), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n672), .B1(new_n712), .B2(new_n704), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1116), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1121), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n893), .B(new_n890), .C1(new_n1124), .C2(new_n848), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n734), .A2(new_n916), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1120), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1119), .A2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1109), .B1(new_n1128), .B2(new_n789), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n642), .A2(G330), .A3(new_n907), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n900), .A2(new_n663), .A3(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n847), .B1(new_n734), .B2(new_n849), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1111), .B1(new_n1132), .B2(new_n1110), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n907), .A2(G330), .A3(new_n849), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(new_n848), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1124), .A2(new_n1135), .A3(new_n1126), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1131), .B1(new_n1133), .B2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1119), .A2(new_n1127), .A3(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1133), .A2(new_n1136), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1131), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n697), .B1(new_n1128), .B2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1129), .B1(new_n1138), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(G378));
  XOR2_X1   g0944(.A(KEYINPUT115), .B(KEYINPUT56), .Z(new_n1145));
  INV_X1    g0945(.A(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n424), .A2(new_n853), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n442), .A2(new_n444), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT55), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n442), .A2(KEYINPUT55), .A3(new_n444), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1147), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(KEYINPUT55), .B1(new_n442), .B2(new_n444), .ZN(new_n1153));
  AOI211_X1 g0953(.A(new_n1149), .B(new_n658), .C1(new_n435), .C2(new_n441), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1147), .ZN(new_n1155));
  NOR3_X1   g0955(.A1(new_n1153), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1146), .B1(new_n1152), .B2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1150), .A2(new_n1147), .A3(new_n1151), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1155), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1158), .A2(new_n1159), .A3(new_n1145), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1157), .A2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(new_n920), .B2(G330), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n872), .A2(new_n873), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n910), .B1(new_n1163), .B2(new_n917), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n890), .A2(KEYINPUT40), .A3(new_n907), .A4(new_n916), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1164), .A2(G330), .A3(new_n1165), .ZN(new_n1166));
  AND3_X1   g0966(.A1(new_n1158), .A2(new_n1159), .A3(new_n1145), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1145), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1166), .A2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n899), .B1(new_n1162), .B2(new_n1170), .ZN(new_n1171));
  AND3_X1   g0971(.A1(new_n874), .A2(new_n897), .A3(new_n898), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n920), .A2(new_n1161), .A3(G330), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1166), .A2(new_n1169), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1172), .A2(new_n1173), .A3(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1171), .A2(KEYINPUT117), .A3(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT117), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1178), .B(new_n899), .C1(new_n1162), .C2(new_n1170), .ZN(new_n1179));
  NAND4_X1  g0979(.A1(new_n1176), .A2(new_n1177), .A3(KEYINPUT57), .A4(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT116), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1171), .A2(new_n1181), .A3(new_n1175), .ZN(new_n1182));
  OAI211_X1 g0982(.A(KEYINPUT116), .B(new_n899), .C1(new_n1162), .C2(new_n1170), .ZN(new_n1183));
  AND3_X1   g0983(.A1(new_n1182), .A2(new_n1183), .A3(new_n1177), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n696), .B(new_n1180), .C1(new_n1184), .C2(KEYINPUT57), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1182), .A2(new_n1014), .A3(new_n1183), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n792), .B1(new_n1169), .B2(new_n818), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n201), .B1(new_n263), .B2(G41), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n837), .A2(new_n1091), .B1(new_n756), .B2(new_n406), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n773), .A2(G128), .ZN(new_n1190));
  INV_X1    g0990(.A(G132), .ZN(new_n1191));
  OAI221_X1 g0991(.A(new_n1190), .B1(new_n754), .B2(new_n1191), .C1(new_n836), .C2(new_n767), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n1189), .B(new_n1192), .C1(new_n780), .C2(new_n1094), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT59), .ZN(new_n1194));
  AOI21_X1  g0994(.A(G33), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n761), .A2(new_n748), .ZN(new_n1196));
  AOI21_X1  g0996(.A(G41), .B1(new_n747), .B2(G124), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1195), .A2(new_n1196), .A3(new_n1197), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1188), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n761), .A2(G58), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n1201), .B(new_n948), .C1(new_n385), .C2(new_n767), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n316), .B(new_n1202), .C1(G116), .C2(new_n770), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n754), .A2(new_n479), .B1(new_n746), .B2(new_n1021), .ZN(new_n1204));
  AOI211_X1 g1004(.A(new_n1028), .B(new_n1204), .C1(G107), .C2(new_n773), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1203), .A2(new_n1205), .A3(new_n286), .ZN(new_n1206));
  XOR2_X1   g1006(.A(new_n1206), .B(KEYINPUT58), .Z(new_n1207));
  OAI21_X1  g1007(.A(new_n793), .B1(new_n1200), .B2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n820), .A2(new_n201), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1187), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1210));
  AND2_X1   g1010(.A1(new_n1186), .A2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1185), .A2(new_n1211), .ZN(G375));
  OAI22_X1  g1012(.A1(new_n837), .A2(new_n1101), .B1(new_n385), .B2(new_n756), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n772), .A2(new_n1021), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n767), .A2(new_n391), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n760), .A2(new_n212), .ZN(new_n1216));
  NOR4_X1   g1016(.A1(new_n1213), .A2(new_n1214), .A3(new_n1215), .A4(new_n1216), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n265), .B1(new_n764), .B2(new_n479), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(G116), .B2(new_n784), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1217), .B(new_n1219), .C1(new_n1017), .C2(new_n746), .ZN(new_n1220));
  XOR2_X1   g1020(.A(new_n1220), .B(KEYINPUT118), .Z(new_n1221));
  NOR2_X1   g1021(.A1(new_n767), .A2(new_n406), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(G159), .A2(new_n780), .B1(new_n747), .B2(G128), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1223), .B(new_n316), .C1(new_n1191), .C2(new_n837), .ZN(new_n1224));
  AOI211_X1 g1024(.A(new_n1222), .B(new_n1224), .C1(G137), .C2(new_n773), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n782), .A2(G50), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n784), .A2(new_n1094), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1225), .A2(new_n1201), .A3(new_n1226), .A4(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n743), .B1(new_n1221), .B2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n818), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n791), .B1(new_n847), .B2(new_n1230), .ZN(new_n1231));
  AOI211_X1 g1031(.A(new_n1229), .B(new_n1231), .C1(new_n203), .C2(new_n820), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(new_n1139), .B2(new_n1014), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1131), .A2(new_n1133), .A3(new_n1136), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(new_n985), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1233), .B1(new_n1235), .B2(new_n1137), .ZN(G381));
  NOR3_X1   g1036(.A1(G390), .A2(G384), .A3(G381), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1046), .A2(new_n809), .A3(new_n1048), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1237), .A2(new_n1006), .A3(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT119), .ZN(new_n1241));
  AND2_X1   g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(G375), .A2(G378), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1243), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1244));
  OR2_X1    g1044(.A1(new_n1242), .A2(new_n1244), .ZN(G407));
  INV_X1    g1045(.A(G213), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1246), .B1(new_n1243), .B2(new_n671), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1247), .B1(new_n1242), .B2(new_n1244), .ZN(G409));
  INV_X1    g1048(.A(KEYINPUT127), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1246), .A2(G343), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(G2897), .ZN(new_n1251));
  AND2_X1   g1051(.A1(new_n1133), .A2(new_n1136), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT121), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1252), .A2(new_n1253), .A3(KEYINPUT60), .A4(new_n1131), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT60), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n697), .B1(new_n1234), .B2(new_n1255), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1131), .A2(new_n1133), .A3(new_n1136), .A4(KEYINPUT60), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1257), .A2(KEYINPUT121), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1254), .A2(new_n1256), .A3(new_n1141), .A4(new_n1258), .ZN(new_n1259));
  AND3_X1   g1059(.A1(new_n1259), .A2(G384), .A3(new_n1233), .ZN(new_n1260));
  AOI21_X1  g1060(.A(G384), .B1(new_n1259), .B2(new_n1233), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT122), .ZN(new_n1262));
  NOR3_X1   g1062(.A1(new_n1260), .A2(new_n1261), .A3(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1254), .A2(new_n1258), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1234), .A2(new_n1255), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1265), .A2(new_n696), .A3(new_n1141), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1233), .B1(new_n1264), .B2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(G384), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1259), .A2(G384), .A3(new_n1233), .ZN(new_n1270));
  AOI21_X1  g1070(.A(KEYINPUT122), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1251), .B1(new_n1263), .B2(new_n1271), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1273), .A2(new_n1251), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1272), .A2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1250), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1185), .A2(G378), .A3(new_n1211), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1182), .A2(new_n1177), .A3(new_n985), .A4(new_n1183), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1176), .A2(new_n1014), .A3(new_n1179), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1279), .A2(new_n1210), .A3(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(new_n1143), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(KEYINPUT120), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT120), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1281), .A2(new_n1284), .A3(new_n1143), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1278), .A2(new_n1283), .A3(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1276), .B1(new_n1277), .B2(new_n1286), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1249), .B1(new_n1287), .B2(KEYINPUT61), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT61), .ZN(new_n1289));
  AND3_X1   g1089(.A1(new_n1281), .A2(new_n1284), .A3(new_n1143), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1284), .B1(new_n1281), .B2(new_n1143), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1250), .B1(new_n1292), .B2(new_n1278), .ZN(new_n1293));
  OAI211_X1 g1093(.A(KEYINPUT127), .B(new_n1289), .C1(new_n1293), .C2(new_n1276), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1262), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1269), .A2(KEYINPUT122), .A3(new_n1270), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1286), .A2(new_n1277), .A3(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(KEYINPUT62), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT62), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1293), .A2(new_n1300), .A3(new_n1297), .ZN(new_n1301));
  NAND4_X1  g1101(.A1(new_n1288), .A2(new_n1294), .A3(new_n1299), .A4(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT125), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n809), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1304));
  OAI22_X1  g1104(.A1(new_n1006), .A2(new_n1303), .B1(new_n1239), .B2(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(G393), .A2(G396), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n985), .B1(new_n1059), .B2(new_n736), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1004), .B1(new_n1307), .B2(new_n789), .ZN(new_n1308));
  OAI211_X1 g1108(.A(new_n1306), .B(new_n1238), .C1(new_n1308), .C2(new_n966), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1305), .A2(new_n1309), .ZN(new_n1310));
  XNOR2_X1  g1110(.A(new_n1310), .B(G390), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1302), .A2(new_n1311), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1272), .A2(new_n1275), .A3(KEYINPUT123), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT123), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1251), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1315), .B1(new_n1295), .B2(new_n1296), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1314), .B1(new_n1316), .B2(new_n1274), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1313), .A2(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1286), .A2(new_n1277), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1320), .A2(KEYINPUT124), .ZN(new_n1321));
  INV_X1    g1121(.A(KEYINPUT124), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1318), .A2(new_n1322), .A3(new_n1319), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1321), .A2(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT126), .ZN(new_n1325));
  NAND4_X1  g1125(.A1(new_n1293), .A2(new_n1325), .A3(KEYINPUT63), .A4(new_n1297), .ZN(new_n1326));
  NAND4_X1  g1126(.A1(new_n1286), .A2(KEYINPUT63), .A3(new_n1277), .A4(new_n1297), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1327), .A2(KEYINPUT126), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1311), .B1(new_n1326), .B2(new_n1328), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT63), .ZN(new_n1330));
  AOI21_X1  g1130(.A(KEYINPUT61), .B1(new_n1298), .B2(new_n1330), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1324), .A2(new_n1329), .A3(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1312), .A2(new_n1332), .ZN(G405));
  INV_X1    g1133(.A(new_n1278), .ZN(new_n1334));
  AOI21_X1  g1134(.A(G378), .B1(new_n1185), .B2(new_n1211), .ZN(new_n1335));
  OAI21_X1  g1135(.A(new_n1297), .B1(new_n1334), .B2(new_n1335), .ZN(new_n1336));
  OR2_X1    g1136(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1337));
  OAI21_X1  g1137(.A(new_n1336), .B1(new_n1337), .B2(new_n1273), .ZN(new_n1338));
  XNOR2_X1  g1138(.A(new_n1338), .B(new_n1311), .ZN(G402));
endmodule


