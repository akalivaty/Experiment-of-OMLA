//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 1 0 1 1 0 0 1 1 1 1 1 0 1 1 0 1 1 1 1 0 1 0 0 0 0 0 0 1 0 0 0 0 0 0 0 1 0 1 0 1 0 0 0 0 0 1 1 1 0 1 1 1 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:47 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n667, new_n668,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n893, new_n894, new_n895, new_n896, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983;
  XOR2_X1   g000(.A(KEYINPUT73), .B(KEYINPUT27), .Z(new_n187));
  INV_X1    g001(.A(G237), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n188), .A2(new_n189), .A3(G210), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n187), .B(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT26), .B(G101), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n191), .B(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(KEYINPUT2), .A2(G113), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT69), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT69), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n197), .A2(KEYINPUT2), .A3(G113), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  NOR2_X1   g013(.A1(KEYINPUT2), .A2(G113), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  XNOR2_X1  g015(.A(G116), .B(G119), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n199), .A2(new_n201), .A3(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(KEYINPUT71), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n200), .B1(new_n196), .B2(new_n198), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT71), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(new_n206), .A3(new_n202), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n204), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT70), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n202), .B1(new_n205), .B2(new_n209), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n197), .B1(KEYINPUT2), .B2(G113), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n195), .A2(KEYINPUT69), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n201), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(KEYINPUT70), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n210), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n208), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT66), .ZN(new_n217));
  INV_X1    g031(.A(G134), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n217), .B1(new_n218), .B2(G137), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(KEYINPUT11), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n218), .A2(G137), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT11), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n217), .B(new_n222), .C1(new_n218), .C2(G137), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n220), .A2(new_n221), .A3(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G131), .ZN(new_n225));
  INV_X1    g039(.A(G131), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n220), .A2(new_n226), .A3(new_n221), .A4(new_n223), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n225), .A2(KEYINPUT67), .A3(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT67), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n224), .A2(new_n229), .A3(G131), .ZN(new_n230));
  NAND2_X1  g044(.A1(KEYINPUT0), .A2(G128), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G143), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(KEYINPUT64), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT64), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G143), .ZN(new_n236));
  INV_X1    g050(.A(G146), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n234), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n237), .A2(G143), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n232), .B1(new_n238), .B2(new_n240), .ZN(new_n241));
  NOR2_X1   g055(.A1(KEYINPUT0), .A2(G128), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n233), .A2(G146), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n234), .A2(new_n236), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n244), .B1(new_n245), .B2(G146), .ZN(new_n246));
  AOI22_X1  g060(.A1(new_n241), .A2(new_n243), .B1(new_n246), .B2(new_n232), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n228), .A2(new_n230), .A3(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n238), .A2(new_n240), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT1), .ZN(new_n250));
  OAI21_X1  g064(.A(G128), .B1(new_n244), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n244), .ZN(new_n253));
  INV_X1    g067(.A(G128), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n254), .A2(KEYINPUT1), .ZN(new_n255));
  XNOR2_X1  g069(.A(KEYINPUT64), .B(G143), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n253), .B(new_n255), .C1(new_n256), .C2(new_n237), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n252), .A2(new_n257), .ZN(new_n258));
  OR2_X1    g072(.A1(new_n218), .A2(G137), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n259), .A2(KEYINPUT68), .A3(new_n221), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n260), .B(G131), .C1(KEYINPUT68), .C2(new_n221), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n258), .A2(new_n261), .A3(new_n227), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n248), .A2(KEYINPUT30), .A3(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n262), .ZN(new_n264));
  AOI211_X1 g078(.A(new_n232), .B(new_n242), .C1(new_n238), .C2(new_n240), .ZN(new_n265));
  AOI211_X1 g079(.A(new_n244), .B(new_n231), .C1(new_n245), .C2(G146), .ZN(new_n266));
  NOR3_X1   g080(.A1(new_n265), .A2(new_n266), .A3(KEYINPUT65), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT65), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n249), .A2(new_n231), .A3(new_n243), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n246), .A2(new_n232), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n268), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  AND2_X1   g086(.A1(new_n228), .A2(new_n230), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n264), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n216), .B(new_n263), .C1(new_n274), .C2(KEYINPUT30), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  AND3_X1   g090(.A1(new_n208), .A2(KEYINPUT72), .A3(new_n215), .ZN(new_n277));
  AOI21_X1  g091(.A(KEYINPUT72), .B1(new_n208), .B2(new_n215), .ZN(new_n278));
  OAI211_X1 g092(.A(new_n262), .B(new_n248), .C1(new_n277), .C2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n194), .B1(new_n276), .B2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT28), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n279), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n248), .A2(new_n262), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n278), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n208), .A2(new_n215), .A3(KEYINPUT72), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(KEYINPUT65), .B1(new_n265), .B2(new_n266), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n269), .A2(new_n270), .A3(new_n268), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n228), .A2(new_n230), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n262), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  AOI22_X1  g108(.A1(new_n286), .A2(new_n289), .B1(new_n294), .B2(new_n216), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n284), .B1(new_n295), .B2(new_n283), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n296), .A2(new_n194), .ZN(new_n297));
  NOR3_X1   g111(.A1(new_n282), .A2(new_n297), .A3(KEYINPUT29), .ZN(new_n298));
  XNOR2_X1  g112(.A(KEYINPUT77), .B(G902), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n277), .A2(new_n278), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(new_n285), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(new_n279), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(KEYINPUT28), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n279), .A2(KEYINPUT76), .A3(new_n283), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT76), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n284), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n304), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n193), .A2(KEYINPUT29), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n300), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(G472), .B1(new_n298), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT32), .ZN(new_n312));
  AND3_X1   g126(.A1(new_n279), .A2(KEYINPUT74), .A3(new_n193), .ZN(new_n313));
  AOI21_X1  g127(.A(KEYINPUT74), .B1(new_n279), .B2(new_n193), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT75), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT31), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n315), .A2(new_n316), .A3(new_n317), .A4(new_n275), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n193), .B1(new_n301), .B2(new_n285), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT74), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n279), .A2(KEYINPUT74), .A3(new_n193), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n321), .A2(new_n275), .A3(new_n317), .A4(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(KEYINPUT75), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n318), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n321), .A2(new_n275), .A3(new_n322), .ZN(new_n326));
  AOI22_X1  g140(.A1(KEYINPUT31), .A2(new_n326), .B1(new_n296), .B2(new_n194), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  NOR2_X1   g142(.A1(G472), .A2(G902), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n312), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n329), .ZN(new_n331));
  AOI211_X1 g145(.A(KEYINPUT32), .B(new_n331), .C1(new_n325), .C2(new_n327), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n311), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  XOR2_X1   g147(.A(KEYINPUT9), .B(G234), .Z(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(G221), .B1(new_n335), .B2(G902), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(G902), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n253), .B1(new_n256), .B2(new_n237), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n250), .B1(new_n256), .B2(new_n237), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n339), .B1(new_n340), .B2(new_n254), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT83), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n246), .A2(new_n342), .A3(new_n255), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n257), .A2(KEYINPUT83), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n341), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(G104), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n346), .A2(G107), .ZN(new_n347));
  INV_X1    g161(.A(G107), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n348), .A2(G104), .ZN(new_n349));
  OAI21_X1  g163(.A(G101), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(KEYINPUT3), .B1(new_n346), .B2(G107), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT82), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n352), .B1(new_n348), .B2(G104), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT3), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n354), .A2(new_n348), .A3(G104), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n346), .A2(KEYINPUT82), .A3(G107), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n351), .A2(new_n353), .A3(new_n355), .A4(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n350), .B1(new_n357), .B2(G101), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(KEYINPUT10), .B1(new_n345), .B2(new_n359), .ZN(new_n360));
  AND2_X1   g174(.A1(new_n353), .A2(new_n356), .ZN(new_n361));
  INV_X1    g175(.A(G101), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n361), .A2(new_n362), .A3(new_n351), .A4(new_n355), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n357), .A2(G101), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n363), .A2(KEYINPUT4), .A3(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT4), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n357), .A2(new_n366), .A3(G101), .ZN(new_n367));
  AND3_X1   g181(.A1(new_n365), .A2(new_n247), .A3(new_n367), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n360), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n358), .A2(KEYINPUT84), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT84), .ZN(new_n371));
  OAI211_X1 g185(.A(new_n371), .B(new_n350), .C1(new_n357), .C2(G101), .ZN(new_n372));
  AND2_X1   g186(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n373), .A2(KEYINPUT85), .A3(KEYINPUT10), .A4(new_n258), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n370), .A2(new_n258), .A3(KEYINPUT10), .A4(new_n372), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT85), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n369), .A2(new_n293), .A3(new_n374), .A4(new_n377), .ZN(new_n378));
  XNOR2_X1  g192(.A(G110), .B(G140), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n189), .A2(G227), .ZN(new_n380));
  XNOR2_X1  g194(.A(new_n379), .B(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n375), .B(KEYINPUT85), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n293), .B1(new_n383), .B2(new_n369), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT12), .ZN(new_n386));
  AND3_X1   g200(.A1(new_n358), .A2(new_n252), .A3(new_n257), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n387), .B1(new_n359), .B2(new_n345), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n386), .B1(new_n388), .B2(new_n293), .ZN(new_n389));
  AND2_X1   g203(.A1(new_n345), .A2(new_n359), .ZN(new_n390));
  OAI211_X1 g204(.A(KEYINPUT12), .B(new_n273), .C1(new_n390), .C2(new_n387), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n381), .B1(new_n392), .B2(new_n378), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n338), .B1(new_n385), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(G469), .ZN(new_n395));
  XOR2_X1   g209(.A(KEYINPUT86), .B(G469), .Z(new_n396));
  NAND3_X1  g210(.A1(new_n369), .A2(new_n377), .A3(new_n374), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(new_n273), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n381), .B1(new_n398), .B2(new_n378), .ZN(new_n399));
  AND3_X1   g213(.A1(new_n392), .A2(new_n378), .A3(new_n381), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n300), .B(new_n396), .C1(new_n399), .C2(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n337), .B1(new_n395), .B2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(G475), .ZN(new_n403));
  XNOR2_X1  g217(.A(G125), .B(G140), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(KEYINPUT16), .ZN(new_n405));
  INV_X1    g219(.A(G140), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(G125), .ZN(new_n407));
  OAI21_X1  g221(.A(KEYINPUT80), .B1(new_n407), .B2(KEYINPUT16), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT80), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT16), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n409), .A2(new_n410), .A3(new_n406), .A4(G125), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n405), .A2(new_n408), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(new_n237), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n405), .A2(G146), .A3(new_n408), .A4(new_n411), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n413), .A2(KEYINPUT81), .A3(new_n414), .ZN(new_n415));
  OR3_X1    g229(.A1(new_n412), .A2(KEYINPUT81), .A3(new_n237), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n188), .A2(new_n189), .A3(G214), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n418), .A2(new_n234), .A3(new_n236), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n233), .A2(new_n188), .A3(new_n189), .A4(G214), .ZN(new_n420));
  AND3_X1   g234(.A1(new_n419), .A2(G131), .A3(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(G131), .B1(new_n419), .B2(new_n420), .ZN(new_n422));
  OR3_X1    g236(.A1(new_n421), .A2(new_n422), .A3(KEYINPUT17), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n421), .A2(KEYINPUT17), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n417), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT89), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT18), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n426), .B1(new_n427), .B2(new_n226), .ZN(new_n428));
  INV_X1    g242(.A(G214), .ZN(new_n429));
  NOR3_X1   g243(.A1(new_n429), .A2(G237), .A3(G953), .ZN(new_n430));
  OAI211_X1 g244(.A(new_n428), .B(new_n420), .C1(new_n245), .C2(new_n430), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n427), .A2(new_n226), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(KEYINPUT89), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(G125), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(G140), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n407), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(G146), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n404), .A2(new_n237), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n419), .A2(KEYINPUT89), .A3(new_n432), .A4(new_n420), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n434), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT90), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND4_X1  g258(.A1(new_n434), .A2(new_n440), .A3(KEYINPUT90), .A4(new_n441), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n425), .A2(new_n446), .ZN(new_n447));
  XNOR2_X1  g261(.A(G113), .B(G122), .ZN(new_n448));
  XNOR2_X1  g262(.A(new_n448), .B(new_n346), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n425), .A2(new_n449), .A3(new_n446), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n403), .B1(new_n453), .B2(new_n338), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n437), .A2(KEYINPUT19), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT19), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n404), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n455), .A2(new_n457), .A3(new_n237), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n414), .B(new_n458), .C1(new_n421), .C2(new_n422), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n446), .A2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT91), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n460), .A2(new_n461), .A3(new_n450), .ZN(new_n462));
  INV_X1    g276(.A(new_n459), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n463), .B1(new_n444), .B2(new_n445), .ZN(new_n464));
  OAI21_X1  g278(.A(KEYINPUT91), .B1(new_n464), .B2(new_n449), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n462), .A2(new_n465), .A3(new_n452), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT20), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n466), .A2(new_n467), .A3(new_n403), .A4(new_n338), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n466), .A2(new_n403), .A3(new_n338), .ZN(new_n469));
  XOR2_X1   g283(.A(KEYINPUT88), .B(KEYINPUT20), .Z(new_n470));
  AOI22_X1  g284(.A1(KEYINPUT92), .A2(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  OR2_X1    g285(.A1(new_n468), .A2(KEYINPUT92), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n454), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  XNOR2_X1  g287(.A(G116), .B(G122), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(new_n348), .ZN(new_n475));
  XOR2_X1   g289(.A(new_n475), .B(KEYINPUT94), .Z(new_n476));
  INV_X1    g290(.A(KEYINPUT14), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(G116), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n479), .A2(KEYINPUT14), .A3(G122), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n478), .A2(G107), .A3(new_n480), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n233), .A2(G128), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n483), .B1(new_n256), .B2(new_n254), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n484), .A2(G134), .ZN(new_n485));
  AND2_X1   g299(.A1(new_n484), .A2(G134), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n476), .B(new_n481), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(G217), .ZN(new_n488));
  NOR3_X1   g302(.A1(new_n335), .A2(new_n488), .A3(G953), .ZN(new_n489));
  OR3_X1    g303(.A1(new_n484), .A2(KEYINPUT93), .A3(G134), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n474), .B(new_n348), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT13), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n245), .A2(new_n492), .A3(G128), .ZN(new_n493));
  OAI211_X1 g307(.A(G134), .B(new_n493), .C1(new_n484), .C2(new_n492), .ZN(new_n494));
  OAI21_X1  g308(.A(KEYINPUT93), .B1(new_n484), .B2(G134), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n490), .A2(new_n491), .A3(new_n494), .A4(new_n495), .ZN(new_n496));
  AND3_X1   g310(.A1(new_n487), .A2(new_n489), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n489), .B1(new_n487), .B2(new_n496), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n499), .A2(new_n299), .ZN(new_n500));
  INV_X1    g314(.A(G478), .ZN(new_n501));
  NOR2_X1   g315(.A1(KEYINPUT95), .A2(KEYINPUT15), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(KEYINPUT95), .A2(KEYINPUT15), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n501), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n500), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n505), .B1(new_n499), .B2(new_n299), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(G234), .A2(G237), .ZN(new_n511));
  AND3_X1   g325(.A1(new_n511), .A2(G952), .A3(new_n189), .ZN(new_n512));
  XNOR2_X1  g326(.A(KEYINPUT21), .B(G898), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n513), .B(KEYINPUT96), .ZN(new_n514));
  AND3_X1   g328(.A1(new_n299), .A2(G953), .A3(new_n511), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n512), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  AND4_X1   g331(.A1(new_n402), .A2(new_n473), .A3(new_n510), .A4(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n254), .A2(G119), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(KEYINPUT79), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT78), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n254), .A2(G119), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT23), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT79), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n519), .A2(new_n526), .ZN(new_n527));
  OAI211_X1 g341(.A(KEYINPUT78), .B(KEYINPUT23), .C1(new_n254), .C2(G119), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n521), .A2(new_n525), .A3(new_n527), .A4(new_n528), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n529), .B1(new_n524), .B2(new_n519), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n520), .A2(new_n523), .ZN(new_n531));
  XOR2_X1   g345(.A(KEYINPUT24), .B(G110), .Z(new_n532));
  OAI22_X1  g346(.A1(new_n530), .A2(G110), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n533), .A2(new_n414), .A3(new_n439), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n530), .A2(G110), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n531), .A2(new_n532), .ZN(new_n536));
  NAND4_X1  g350(.A1(new_n535), .A2(new_n415), .A3(new_n416), .A4(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n189), .A2(G221), .A3(G234), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n539), .B(KEYINPUT22), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n540), .B(G137), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n538), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n534), .A2(new_n537), .A3(new_n541), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n543), .A2(new_n300), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(KEYINPUT25), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n488), .B1(new_n300), .B2(G234), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT25), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n543), .A2(new_n548), .A3(new_n300), .A4(new_n544), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n546), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  AND2_X1   g364(.A1(new_n543), .A2(new_n544), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n547), .A2(G902), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AND2_X1   g367(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  OAI21_X1  g368(.A(G214), .B1(G237), .B2(G902), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n202), .A2(KEYINPUT5), .ZN(new_n557));
  OR2_X1    g371(.A1(new_n479), .A2(G119), .ZN(new_n558));
  OAI211_X1 g372(.A(new_n557), .B(G113), .C1(KEYINPUT5), .C2(new_n558), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n370), .A2(new_n208), .A3(new_n372), .A4(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n216), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n365), .A2(new_n367), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  XOR2_X1   g377(.A(G110), .B(G122), .Z(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n564), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n560), .B(new_n566), .C1(new_n561), .C2(new_n562), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n565), .A2(KEYINPUT6), .A3(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT6), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n563), .A2(new_n569), .A3(new_n564), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n252), .A2(new_n435), .A3(new_n257), .ZN(new_n571));
  OAI211_X1 g385(.A(KEYINPUT87), .B(new_n571), .C1(new_n247), .C2(new_n435), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n189), .A2(G224), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT87), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n574), .B(G125), .C1(new_n265), .C2(new_n266), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n572), .A2(new_n573), .A3(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n573), .B1(new_n572), .B2(new_n575), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n568), .A2(new_n570), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n208), .A2(new_n559), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n581), .B(new_n358), .ZN(new_n582));
  XOR2_X1   g396(.A(new_n564), .B(KEYINPUT8), .Z(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n573), .A2(KEYINPUT7), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n572), .A2(new_n575), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n572), .A2(new_n575), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n587), .A2(KEYINPUT7), .A3(new_n573), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n584), .A2(new_n586), .A3(new_n567), .A4(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n580), .A2(new_n338), .A3(new_n589), .ZN(new_n590));
  OAI21_X1  g404(.A(G210), .B1(G237), .B2(G902), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n580), .A2(new_n338), .A3(new_n591), .A4(new_n589), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n556), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n333), .A2(new_n518), .A3(new_n554), .A4(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n596), .B(G101), .ZN(G3));
  INV_X1    g411(.A(G472), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n598), .B1(new_n328), .B2(new_n300), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n392), .A2(new_n378), .ZN(new_n600));
  INV_X1    g414(.A(new_n381), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n398), .A2(new_n378), .A3(new_n381), .ZN(new_n603));
  AOI21_X1  g417(.A(G902), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(G469), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n401), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n606), .A2(new_n554), .A3(new_n336), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n331), .B1(new_n325), .B2(new_n327), .ZN(new_n608));
  NOR3_X1   g422(.A1(new_n599), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n595), .A2(new_n517), .ZN(new_n610));
  INV_X1    g424(.A(new_n499), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n487), .A2(new_n496), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(KEYINPUT97), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(KEYINPUT33), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n499), .A2(KEYINPUT33), .A3(new_n613), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n615), .A2(new_n300), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(G478), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n500), .A2(new_n501), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NOR3_X1   g434(.A1(new_n610), .A2(new_n473), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n609), .A2(new_n621), .ZN(new_n622));
  XOR2_X1   g436(.A(KEYINPUT34), .B(G104), .Z(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(G6));
  OR2_X1    g438(.A1(new_n469), .A2(new_n470), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n469), .A2(new_n470), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n454), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(new_n509), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n628), .A2(new_n610), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n609), .A2(new_n629), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT35), .B(G107), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G9));
  NOR2_X1   g446(.A1(new_n599), .A2(new_n608), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n542), .A2(KEYINPUT36), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n538), .B(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(new_n552), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n550), .A2(new_n636), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n518), .A2(new_n595), .A3(new_n633), .A4(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(new_n638), .B(KEYINPUT37), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(G110), .ZN(G12));
  NAND2_X1  g454(.A1(new_n606), .A2(new_n336), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n593), .A2(new_n594), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n555), .ZN(new_n643));
  INV_X1    g457(.A(new_n637), .ZN(new_n644));
  NOR3_X1   g458(.A1(new_n641), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(G900), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n512), .B1(new_n515), .B2(new_n646), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n628), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n333), .A2(new_n645), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(G128), .ZN(G30));
  XNOR2_X1  g464(.A(new_n642), .B(KEYINPUT98), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(KEYINPUT38), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n652), .A2(new_n637), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n647), .B(KEYINPUT39), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n402), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(new_n656), .B(KEYINPUT40), .Z(new_n657));
  AOI22_X1  g471(.A1(new_n315), .A2(new_n275), .B1(new_n194), .B2(new_n303), .ZN(new_n658));
  OAI21_X1  g472(.A(G472), .B1(new_n658), .B2(G902), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n659), .B1(new_n330), .B2(new_n332), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n473), .A2(new_n510), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n555), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n653), .A2(new_n657), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(new_n256), .ZN(G45));
  NOR3_X1   g480(.A1(new_n473), .A2(new_n620), .A3(new_n647), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n333), .A2(new_n645), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G146), .ZN(G48));
  INV_X1    g483(.A(new_n554), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n326), .A2(KEYINPUT31), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n296), .A2(new_n194), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n673), .B1(new_n318), .B2(new_n324), .ZN(new_n674));
  OAI21_X1  g488(.A(KEYINPUT32), .B1(new_n674), .B2(new_n331), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n608), .A2(new_n312), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n670), .B1(new_n677), .B2(new_n311), .ZN(new_n678));
  INV_X1    g492(.A(new_n378), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n601), .B1(new_n679), .B2(new_n384), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n392), .A2(new_n378), .A3(new_n381), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n299), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  OAI211_X1 g496(.A(new_n401), .B(new_n336), .C1(new_n682), .C2(new_n605), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n678), .A2(KEYINPUT99), .A3(new_n621), .A4(new_n684), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n333), .A2(new_n621), .A3(new_n554), .A4(new_n684), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT99), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(KEYINPUT41), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G113), .ZN(G15));
  NAND4_X1  g505(.A1(new_n333), .A2(new_n629), .A3(new_n554), .A4(new_n684), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G116), .ZN(G18));
  INV_X1    g507(.A(KEYINPUT100), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n684), .A2(new_n694), .A3(new_n595), .ZN(new_n695));
  OAI21_X1  g509(.A(KEYINPUT100), .B1(new_n643), .B2(new_n683), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(new_n454), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n468), .A2(KEYINPUT92), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(new_n626), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n468), .A2(KEYINPUT92), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n698), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NOR3_X1   g516(.A1(new_n702), .A2(new_n516), .A3(new_n509), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n697), .A2(new_n333), .A3(new_n703), .A4(new_n637), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G119), .ZN(G21));
  XOR2_X1   g519(.A(new_n329), .B(KEYINPUT101), .Z(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  AOI22_X1  g521(.A1(new_n318), .A2(new_n324), .B1(new_n194), .B2(new_n308), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n707), .B1(new_n708), .B2(new_n671), .ZN(new_n709));
  NOR3_X1   g523(.A1(new_n599), .A2(new_n709), .A3(new_n670), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n662), .A2(new_n595), .A3(new_n517), .A4(new_n684), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  XOR2_X1   g527(.A(new_n713), .B(G122), .Z(G24));
  NOR3_X1   g528(.A1(new_n599), .A2(new_n709), .A3(new_n644), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n697), .A2(new_n667), .A3(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G125), .ZN(G27));
  INV_X1    g531(.A(KEYINPUT102), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n593), .A2(new_n555), .A3(new_n594), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n718), .B1(new_n641), .B2(new_n719), .ZN(new_n720));
  AND3_X1   g534(.A1(new_n593), .A2(new_n555), .A3(new_n594), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n402), .A2(KEYINPUT102), .A3(new_n721), .ZN(new_n722));
  AND4_X1   g536(.A1(KEYINPUT42), .A2(new_n720), .A3(new_n667), .A4(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT103), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n675), .A2(new_n724), .A3(new_n676), .ZN(new_n725));
  OAI21_X1  g539(.A(KEYINPUT103), .B1(new_n330), .B2(new_n332), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n725), .A2(new_n726), .A3(new_n311), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n723), .A2(new_n554), .A3(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT42), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n333), .A2(new_n554), .A3(new_n720), .A4(new_n722), .ZN(new_n730));
  INV_X1    g544(.A(new_n667), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n729), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n728), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(KEYINPUT104), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT104), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n728), .A2(new_n732), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G131), .ZN(G33));
  INV_X1    g552(.A(new_n730), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(new_n648), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G134), .ZN(G36));
  AND2_X1   g555(.A1(new_n618), .A2(new_n619), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n473), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(KEYINPUT43), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n644), .B1(new_n744), .B2(KEYINPUT106), .ZN(new_n745));
  INV_X1    g559(.A(new_n633), .ZN(new_n746));
  OAI211_X1 g560(.A(new_n745), .B(new_n746), .C1(KEYINPUT106), .C2(new_n744), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT44), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n719), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n602), .A2(new_n603), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(KEYINPUT45), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(G469), .ZN(new_n752));
  NAND2_X1  g566(.A1(G469), .A2(G902), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n752), .A2(KEYINPUT46), .A3(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT46), .ZN(new_n755));
  OAI211_X1 g569(.A(new_n755), .B(G469), .C1(new_n751), .C2(G902), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n754), .A2(new_n401), .A3(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n757), .A2(new_n336), .A3(new_n655), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT105), .ZN(new_n759));
  OR2_X1    g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n758), .A2(new_n759), .ZN(new_n761));
  AND2_X1   g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  OAI211_X1 g576(.A(new_n749), .B(new_n762), .C1(new_n748), .C2(new_n747), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G137), .ZN(G39));
  INV_X1    g578(.A(KEYINPUT47), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT107), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n757), .A2(new_n766), .A3(new_n336), .ZN(new_n767));
  INV_X1    g581(.A(new_n767), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n766), .B1(new_n757), .B2(new_n336), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n765), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(new_n769), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n771), .A2(KEYINPUT47), .A3(new_n767), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n731), .A2(new_n333), .A3(new_n719), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n770), .A2(new_n772), .A3(new_n670), .A4(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(KEYINPUT108), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G140), .ZN(G42));
  XOR2_X1   g590(.A(new_n743), .B(KEYINPUT43), .Z(new_n777));
  NAND3_X1  g591(.A1(new_n777), .A2(new_n512), .A3(new_n710), .ZN(new_n778));
  INV_X1    g592(.A(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(new_n697), .ZN(new_n780));
  AND3_X1   g594(.A1(new_n684), .A2(new_n512), .A3(new_n721), .ZN(new_n781));
  AND3_X1   g595(.A1(new_n661), .A2(new_n554), .A3(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n782), .A2(new_n702), .A3(new_n742), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n780), .A2(G952), .A3(new_n189), .A4(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(KEYINPUT117), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n777), .A2(new_n781), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n727), .A2(new_n554), .ZN(new_n787));
  INV_X1    g601(.A(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(KEYINPUT48), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n785), .A2(new_n790), .ZN(new_n791));
  XOR2_X1   g605(.A(new_n791), .B(KEYINPUT118), .Z(new_n792));
  INV_X1    g606(.A(KEYINPUT50), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n683), .A2(new_n555), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(KEYINPUT114), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n652), .A2(new_n795), .ZN(new_n796));
  XOR2_X1   g610(.A(new_n796), .B(KEYINPUT115), .Z(new_n797));
  AOI21_X1  g611(.A(new_n793), .B1(new_n797), .B2(new_n779), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n793), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n401), .B1(new_n682), .B2(new_n605), .ZN(new_n800));
  INV_X1    g614(.A(new_n800), .ZN(new_n801));
  AOI22_X1  g615(.A1(new_n770), .A2(new_n772), .B1(new_n337), .B2(new_n801), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n799), .B1(new_n802), .B2(new_n719), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n798), .B1(new_n803), .B2(new_n779), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n786), .A2(new_n715), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n782), .A2(new_n473), .A3(new_n620), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(KEYINPUT116), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n804), .A2(new_n805), .A3(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT51), .ZN(new_n809));
  OR2_X1    g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT54), .ZN(new_n811));
  OAI21_X1  g625(.A(KEYINPUT109), .B1(new_n473), .B2(new_n620), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT109), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n702), .A2(new_n742), .A3(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT110), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n509), .B(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(new_n473), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n812), .A2(new_n814), .A3(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(new_n610), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n818), .A2(new_n609), .A3(new_n819), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n715), .A2(new_n667), .A3(new_n720), .A4(new_n722), .ZN(new_n821));
  AND4_X1   g635(.A1(new_n596), .A2(new_n820), .A3(new_n638), .A4(new_n821), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n644), .B1(new_n677), .B2(new_n311), .ZN(new_n823));
  INV_X1    g637(.A(new_n816), .ZN(new_n824));
  INV_X1    g638(.A(new_n647), .ZN(new_n825));
  AND4_X1   g639(.A1(new_n402), .A2(new_n627), .A3(new_n721), .A4(new_n825), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n823), .A2(KEYINPUT111), .A3(new_n824), .A4(new_n826), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n333), .A2(new_n826), .A3(new_n637), .A4(new_n824), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT111), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n827), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n822), .A2(new_n831), .A3(new_n740), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n832), .B(KEYINPUT113), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n704), .A2(new_n692), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n713), .B1(new_n685), .B2(new_n688), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n702), .A2(new_n555), .A3(new_n642), .A4(new_n509), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n836), .A2(new_n637), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n837), .A2(new_n402), .A3(new_n825), .A4(new_n660), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n333), .B(new_n645), .C1(new_n648), .C2(new_n667), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n838), .A2(new_n716), .A3(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT52), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n840), .A2(new_n841), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n834), .B(new_n835), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n833), .A2(KEYINPUT53), .A3(new_n733), .A4(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT53), .ZN(new_n847));
  AOI22_X1  g661(.A1(new_n827), .A2(new_n830), .B1(new_n739), .B2(new_n648), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n728), .A2(new_n732), .A3(new_n735), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n735), .B1(new_n728), .B2(new_n732), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n822), .B(new_n848), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  OAI211_X1 g665(.A(KEYINPUT112), .B(new_n847), .C1(new_n851), .C2(new_n844), .ZN(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n840), .B(new_n841), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n822), .A2(new_n740), .A3(new_n831), .ZN(new_n855));
  INV_X1    g669(.A(new_n713), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n689), .A2(new_n856), .A3(new_n834), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n737), .A2(new_n854), .A3(new_n855), .A4(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(KEYINPUT112), .B1(new_n858), .B2(new_n847), .ZN(new_n859));
  OAI211_X1 g673(.A(new_n811), .B(new_n846), .C1(new_n853), .C2(new_n859), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n858), .A2(new_n847), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n858), .A2(new_n847), .ZN(new_n862));
  OAI21_X1  g676(.A(KEYINPUT54), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n808), .A2(new_n809), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n792), .A2(new_n810), .A3(new_n864), .A4(new_n865), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n866), .B1(G952), .B2(G953), .ZN(new_n867));
  XOR2_X1   g681(.A(new_n800), .B(KEYINPUT49), .Z(new_n868));
  NAND3_X1  g682(.A1(new_n652), .A2(new_n554), .A3(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n869), .A2(new_n743), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n870), .A2(new_n555), .A3(new_n336), .A4(new_n661), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n867), .A2(new_n871), .ZN(G75));
  OAI21_X1  g686(.A(new_n846), .B1(new_n853), .B2(new_n859), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(new_n299), .ZN(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(new_n592), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT56), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n568), .A2(new_n570), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n878), .B(new_n579), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n879), .B(KEYINPUT55), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n876), .A2(new_n877), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n880), .B1(new_n876), .B2(new_n877), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n189), .A2(G952), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(G51));
  NAND2_X1  g698(.A1(new_n873), .A2(KEYINPUT54), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(new_n860), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n753), .A2(KEYINPUT57), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n753), .A2(KEYINPUT57), .ZN(new_n889));
  OAI22_X1  g703(.A1(new_n888), .A2(new_n889), .B1(new_n399), .B2(new_n400), .ZN(new_n890));
  OR2_X1    g704(.A1(new_n874), .A2(new_n752), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n883), .B1(new_n890), .B2(new_n891), .ZN(G54));
  NAND3_X1  g706(.A1(new_n875), .A2(KEYINPUT58), .A3(G475), .ZN(new_n893));
  INV_X1    g707(.A(new_n466), .ZN(new_n894));
  AND2_X1   g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n893), .A2(new_n894), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n895), .A2(new_n896), .A3(new_n883), .ZN(G60));
  XOR2_X1   g711(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n898));
  NOR2_X1   g712(.A1(new_n501), .A2(new_n338), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n898), .B(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n901), .B1(new_n860), .B2(new_n863), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n615), .A2(new_n616), .ZN(new_n903));
  INV_X1    g717(.A(new_n903), .ZN(new_n904));
  OAI21_X1  g718(.A(KEYINPUT121), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT120), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n903), .A2(new_n901), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n906), .B1(new_n886), .B2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(new_n907), .ZN(new_n909));
  AOI211_X1 g723(.A(KEYINPUT120), .B(new_n909), .C1(new_n885), .C2(new_n860), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n905), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(new_n883), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n903), .B1(new_n864), .B2(new_n901), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n912), .B1(new_n913), .B2(KEYINPUT121), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n911), .A2(new_n914), .ZN(G63));
  NAND2_X1  g729(.A1(G217), .A2(G902), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n916), .B(KEYINPUT60), .Z(new_n917));
  NAND3_X1  g731(.A1(new_n873), .A2(new_n635), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(new_n912), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n551), .B1(new_n873), .B2(new_n917), .ZN(new_n920));
  OAI21_X1  g734(.A(KEYINPUT122), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  XNOR2_X1  g735(.A(KEYINPUT123), .B(KEYINPUT61), .ZN(new_n922));
  INV_X1    g736(.A(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  OAI211_X1 g738(.A(KEYINPUT122), .B(new_n922), .C1(new_n919), .C2(new_n920), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(G66));
  AND3_X1   g740(.A1(new_n820), .A2(new_n596), .A3(new_n638), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n857), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(new_n189), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT124), .ZN(new_n930));
  INV_X1    g744(.A(G224), .ZN(new_n931));
  OAI21_X1  g745(.A(G953), .B1(new_n514), .B2(new_n931), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n932), .B(KEYINPUT125), .Z(new_n933));
  NAND2_X1  g747(.A1(new_n930), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n878), .B1(G898), .B2(new_n189), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n934), .B(new_n935), .ZN(G69));
  AOI21_X1  g750(.A(new_n189), .B1(G227), .B2(G900), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n747), .A2(new_n748), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n721), .ZN(new_n939));
  OAI211_X1 g753(.A(new_n761), .B(new_n760), .C1(new_n747), .C2(new_n748), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n774), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  AND2_X1   g756(.A1(new_n716), .A2(new_n839), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n665), .A2(new_n943), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(KEYINPUT62), .Z(new_n945));
  NOR2_X1   g759(.A1(new_n656), .A2(new_n719), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n678), .A2(new_n818), .A3(new_n946), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n942), .A2(new_n945), .A3(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n263), .B1(new_n274), .B2(KEYINPUT30), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n455), .A2(new_n457), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n950), .B(new_n951), .ZN(new_n952));
  NOR3_X1   g766(.A1(new_n949), .A2(G953), .A3(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(new_n737), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n941), .A2(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT126), .ZN(new_n956));
  INV_X1    g770(.A(new_n836), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n762), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n943), .B1(new_n958), .B2(new_n787), .ZN(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n955), .A2(new_n956), .A3(new_n740), .A4(new_n960), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n763), .A2(new_n737), .A3(new_n740), .A4(new_n774), .ZN(new_n962));
  OAI21_X1  g776(.A(KEYINPUT126), .B1(new_n962), .B2(new_n959), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n961), .A2(new_n963), .A3(new_n189), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n964), .B1(new_n646), .B2(new_n189), .ZN(new_n965));
  AOI211_X1 g779(.A(new_n937), .B(new_n953), .C1(new_n965), .C2(new_n952), .ZN(new_n966));
  NAND2_X1  g780(.A1(G227), .A2(G900), .ZN(new_n967));
  AND4_X1   g781(.A1(G953), .A2(new_n965), .A3(new_n967), .A4(new_n952), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n966), .A2(new_n968), .ZN(G72));
  NAND2_X1  g783(.A1(G472), .A2(G902), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n970), .B(KEYINPUT63), .Z(new_n971));
  OAI21_X1  g785(.A(new_n971), .B1(new_n948), .B2(new_n928), .ZN(new_n972));
  OAI211_X1 g786(.A(new_n972), .B(new_n193), .C1(new_n276), .C2(new_n280), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n281), .A2(new_n326), .ZN(new_n974));
  OAI211_X1 g788(.A(new_n971), .B(new_n974), .C1(new_n861), .C2(new_n862), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n973), .A2(new_n912), .A3(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(new_n928), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n961), .A2(new_n963), .A3(new_n977), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n978), .A2(KEYINPUT127), .A3(new_n971), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n276), .A2(new_n280), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g795(.A(KEYINPUT127), .B1(new_n978), .B2(new_n971), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n976), .B1(new_n983), .B2(new_n194), .ZN(G57));
endmodule


