

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737;

  XNOR2_X2 U376 ( .A(n546), .B(KEYINPUT104), .ZN(n735) );
  XNOR2_X1 U377 ( .A(n536), .B(KEYINPUT40), .ZN(n734) );
  NOR2_X1 U378 ( .A1(n643), .A2(n571), .ZN(n536) );
  XNOR2_X2 U379 ( .A(n432), .B(n479), .ZN(n568) );
  NOR2_X2 U380 ( .A1(n592), .A2(n591), .ZN(n593) );
  BUF_X1 U381 ( .A(n658), .Z(n355) );
  BUF_X2 U382 ( .A(n658), .Z(n356) );
  XNOR2_X1 U383 ( .A(n495), .B(n494), .ZN(n658) );
  XNOR2_X2 U384 ( .A(n390), .B(KEYINPUT22), .ZN(n436) );
  NOR2_X2 U385 ( .A1(n605), .A2(n420), .ZN(n390) );
  NOR2_X1 U386 ( .A1(n734), .A2(n731), .ZN(n425) );
  AND2_X2 U387 ( .A1(n417), .A2(n414), .ZN(n698) );
  NAND2_X1 U388 ( .A1(n415), .A2(n368), .ZN(n414) );
  XNOR2_X1 U389 ( .A(n425), .B(KEYINPUT46), .ZN(n422) );
  XNOR2_X1 U390 ( .A(n444), .B(KEYINPUT32), .ZN(n737) );
  XNOR2_X1 U391 ( .A(n550), .B(KEYINPUT74), .ZN(n641) );
  XNOR2_X1 U392 ( .A(n395), .B(n365), .ZN(n592) );
  XNOR2_X1 U393 ( .A(n397), .B(n589), .ZN(n676) );
  NOR2_X1 U394 ( .A1(n588), .A2(n601), .ZN(n397) );
  XNOR2_X1 U395 ( .A(n555), .B(KEYINPUT19), .ZN(n577) );
  XNOR2_X1 U396 ( .A(n500), .B(n447), .ZN(n527) );
  XNOR2_X1 U397 ( .A(n398), .B(n519), .ZN(n693) );
  XNOR2_X1 U398 ( .A(n718), .B(G146), .ZN(n519) );
  XNOR2_X1 U399 ( .A(n721), .B(n430), .ZN(n429) );
  XNOR2_X1 U400 ( .A(n475), .B(KEYINPUT4), .ZN(n485) );
  XNOR2_X1 U401 ( .A(n435), .B(G110), .ZN(n421) );
  INV_X1 U402 ( .A(G119), .ZN(n435) );
  XNOR2_X1 U403 ( .A(G104), .B(G122), .ZN(n470) );
  INV_X2 U404 ( .A(G128), .ZN(n376) );
  XNOR2_X1 U405 ( .A(n429), .B(n426), .ZN(n619) );
  XNOR2_X2 U406 ( .A(n615), .B(n614), .ZN(n709) );
  NOR2_X1 U407 ( .A1(G237), .A2(G953), .ZN(n455) );
  XNOR2_X1 U408 ( .A(n474), .B(KEYINPUT10), .ZN(n452) );
  INV_X1 U409 ( .A(n722), .ZN(n403) );
  XNOR2_X1 U410 ( .A(n544), .B(n480), .ZN(n667) );
  INV_X1 U411 ( .A(KEYINPUT38), .ZN(n480) );
  INV_X1 U412 ( .A(G469), .ZN(n521) );
  OR2_X1 U413 ( .A1(n527), .A2(n411), .ZN(n552) );
  XNOR2_X1 U414 ( .A(G140), .B(G137), .ZN(n514) );
  NAND2_X1 U415 ( .A1(n423), .A2(n422), .ZN(n424) );
  OR2_X1 U416 ( .A1(G902), .A2(G237), .ZN(n481) );
  INV_X1 U417 ( .A(n600), .ZN(n588) );
  NOR2_X1 U418 ( .A1(n552), .A2(n356), .ZN(n410) );
  AND2_X1 U419 ( .A1(n527), .A2(n359), .ZN(n653) );
  XNOR2_X1 U420 ( .A(n519), .B(n493), .ZN(n623) );
  XNOR2_X1 U421 ( .A(n613), .B(KEYINPUT80), .ZN(n614) );
  XNOR2_X1 U422 ( .A(n448), .B(KEYINPUT24), .ZN(n431) );
  XNOR2_X1 U423 ( .A(G128), .B(KEYINPUT23), .ZN(n448) );
  XNOR2_X1 U424 ( .A(n452), .B(n514), .ZN(n721) );
  XNOR2_X1 U425 ( .A(n428), .B(n427), .ZN(n463) );
  INV_X1 U426 ( .A(KEYINPUT8), .ZN(n427) );
  NAND2_X1 U427 ( .A1(n476), .A2(G234), .ZN(n428) );
  XNOR2_X1 U428 ( .A(G140), .B(G143), .ZN(n449) );
  XNOR2_X1 U429 ( .A(KEYINPUT11), .B(KEYINPUT95), .ZN(n451) );
  XNOR2_X1 U430 ( .A(n520), .B(n518), .ZN(n398) );
  XNOR2_X1 U431 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U432 ( .A(KEYINPUT82), .B(KEYINPUT39), .ZN(n534) );
  NAND2_X1 U433 ( .A1(n568), .A2(n563), .ZN(n555) );
  NAND2_X1 U434 ( .A1(n676), .A2(n602), .ZN(n395) );
  NOR2_X1 U435 ( .A1(n442), .A2(n527), .ZN(n441) );
  NOR2_X1 U436 ( .A1(n579), .A2(KEYINPUT65), .ZN(n442) );
  NAND2_X1 U437 ( .A1(n698), .A2(G472), .ZN(n386) );
  XNOR2_X1 U438 ( .A(n623), .B(KEYINPUT62), .ZN(n624) );
  NOR2_X1 U439 ( .A1(n476), .A2(G952), .ZN(n708) );
  NOR2_X1 U440 ( .A1(n686), .A2(n685), .ZN(n375) );
  NOR2_X1 U441 ( .A1(n641), .A2(n551), .ZN(n371) );
  NAND2_X1 U442 ( .A1(n650), .A2(n560), .ZN(n408) );
  XNOR2_X1 U443 ( .A(n583), .B(KEYINPUT84), .ZN(n584) );
  AND2_X1 U444 ( .A1(n407), .A2(n405), .ZN(n423) );
  NOR2_X1 U445 ( .A1(n408), .A2(n370), .ZN(n407) );
  XNOR2_X1 U446 ( .A(n406), .B(KEYINPUT77), .ZN(n405) );
  XNOR2_X1 U447 ( .A(n371), .B(KEYINPUT68), .ZN(n370) );
  XOR2_X1 U448 ( .A(KEYINPUT5), .B(G116), .Z(n487) );
  XNOR2_X1 U449 ( .A(G137), .B(G119), .ZN(n486) );
  XOR2_X1 U450 ( .A(G104), .B(G101), .Z(n513) );
  INV_X1 U451 ( .A(G107), .ZN(n516) );
  XNOR2_X1 U452 ( .A(G101), .B(KEYINPUT66), .ZN(n472) );
  XOR2_X1 U453 ( .A(G113), .B(KEYINPUT3), .Z(n473) );
  XNOR2_X1 U454 ( .A(G107), .B(G116), .ZN(n471) );
  AND2_X1 U455 ( .A1(n399), .A2(n402), .ZN(n387) );
  NAND2_X1 U456 ( .A1(n400), .A2(n416), .ZN(n401) );
  NAND2_X1 U457 ( .A1(n403), .A2(n404), .ZN(n400) );
  XNOR2_X1 U458 ( .A(n478), .B(KEYINPUT86), .ZN(n384) );
  XOR2_X1 U459 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n478) );
  NAND2_X1 U460 ( .A1(n378), .A2(n377), .ZN(n380) );
  INV_X1 U461 ( .A(KEYINPUT2), .ZN(n377) );
  XNOR2_X1 U462 ( .A(n418), .B(n379), .ZN(n417) );
  NOR2_X1 U463 ( .A1(n688), .A2(n616), .ZN(n432) );
  XNOR2_X1 U464 ( .A(n483), .B(KEYINPUT41), .ZN(n666) );
  XNOR2_X1 U465 ( .A(n562), .B(n393), .ZN(n554) );
  INV_X1 U466 ( .A(KEYINPUT107), .ZN(n393) );
  XNOR2_X1 U467 ( .A(n604), .B(KEYINPUT102), .ZN(n531) );
  XNOR2_X1 U468 ( .A(n410), .B(n409), .ZN(n524) );
  INV_X1 U469 ( .A(KEYINPUT28), .ZN(n409) );
  XNOR2_X1 U470 ( .A(n446), .B(KEYINPUT0), .ZN(n605) );
  NAND2_X1 U471 ( .A1(n557), .A2(n653), .ZN(n604) );
  XNOR2_X1 U472 ( .A(n355), .B(KEYINPUT6), .ZN(n600) );
  XNOR2_X1 U473 ( .A(n385), .B(n491), .ZN(n412) );
  XNOR2_X1 U474 ( .A(n434), .B(n433), .ZN(n385) );
  XNOR2_X1 U475 ( .A(n471), .B(KEYINPUT16), .ZN(n433) );
  XNOR2_X1 U476 ( .A(n421), .B(n470), .ZN(n434) );
  AND2_X1 U477 ( .A1(n463), .A2(G221), .ZN(n426) );
  XNOR2_X1 U478 ( .A(n464), .B(n394), .ZN(n704) );
  XNOR2_X1 U479 ( .A(n466), .B(n465), .ZN(n394) );
  XNOR2_X1 U480 ( .A(n457), .B(n456), .ZN(n700) );
  XNOR2_X1 U481 ( .A(n453), .B(n396), .ZN(n457) );
  XNOR2_X1 U482 ( .A(n362), .B(n454), .ZN(n396) );
  XNOR2_X1 U483 ( .A(n412), .B(n381), .ZN(n688) );
  XNOR2_X1 U484 ( .A(n383), .B(n382), .ZN(n381) );
  XNOR2_X1 U485 ( .A(n485), .B(n384), .ZN(n383) );
  XNOR2_X1 U486 ( .A(n477), .B(n474), .ZN(n382) );
  NAND2_X1 U487 ( .A1(n436), .A2(n445), .ZN(n444) );
  AND2_X1 U488 ( .A1(n582), .A2(n360), .ZN(n445) );
  NAND2_X1 U489 ( .A1(n439), .A2(n438), .ZN(n437) );
  AND2_X1 U490 ( .A1(n443), .A2(n441), .ZN(n440) );
  INV_X1 U491 ( .A(KEYINPUT65), .ZN(n438) );
  XNOR2_X1 U492 ( .A(n386), .B(n624), .ZN(n625) );
  INV_X1 U493 ( .A(n708), .ZN(n391) );
  INV_X1 U494 ( .A(KEYINPUT53), .ZN(n372) );
  XNOR2_X1 U495 ( .A(n375), .B(KEYINPUT118), .ZN(n374) );
  AND2_X1 U496 ( .A1(n363), .A2(n358), .ZN(n357) );
  AND2_X1 U497 ( .A1(n652), .A2(n367), .ZN(n358) );
  XOR2_X1 U498 ( .A(n503), .B(n502), .Z(n359) );
  XOR2_X1 U499 ( .A(n588), .B(KEYINPUT73), .Z(n360) );
  XNOR2_X1 U500 ( .A(KEYINPUT76), .B(n617), .ZN(n361) );
  AND2_X1 U501 ( .A1(G214), .A2(n488), .ZN(n362) );
  AND2_X1 U502 ( .A1(n570), .A2(n732), .ZN(n363) );
  AND2_X1 U503 ( .A1(n579), .A2(KEYINPUT65), .ZN(n364) );
  XOR2_X1 U504 ( .A(n586), .B(KEYINPUT67), .Z(n365) );
  XOR2_X1 U505 ( .A(G902), .B(KEYINPUT15), .Z(n616) );
  XNOR2_X1 U506 ( .A(n485), .B(n484), .ZN(n718) );
  XOR2_X1 U507 ( .A(n561), .B(KEYINPUT81), .Z(n366) );
  AND2_X1 U508 ( .A1(n404), .A2(KEYINPUT79), .ZN(n367) );
  NAND2_X1 U509 ( .A1(n616), .A2(KEYINPUT2), .ZN(n368) );
  INV_X1 U510 ( .A(KEYINPUT79), .ZN(n416) );
  NOR2_X1 U511 ( .A1(n412), .A2(n716), .ZN(n369) );
  INV_X1 U512 ( .A(G953), .ZN(n572) );
  XNOR2_X1 U513 ( .A(n373), .B(n372), .ZN(G75) );
  NAND2_X1 U514 ( .A1(n374), .A2(n572), .ZN(n373) );
  XNOR2_X2 U515 ( .A(n376), .B(G143), .ZN(n475) );
  NAND2_X1 U516 ( .A1(n403), .A2(n388), .ZN(n378) );
  AND2_X1 U517 ( .A1(n380), .A2(n417), .ZN(n686) );
  INV_X1 U518 ( .A(KEYINPUT71), .ZN(n379) );
  OR2_X1 U519 ( .A1(n733), .A2(KEYINPUT44), .ZN(n595) );
  NOR2_X2 U520 ( .A1(n691), .A2(n708), .ZN(n692) );
  NAND2_X1 U521 ( .A1(n737), .A2(n413), .ZN(n585) );
  NAND2_X1 U522 ( .A1(n698), .A2(G217), .ZN(n618) );
  NAND2_X1 U523 ( .A1(n401), .A2(n387), .ZN(n415) );
  NOR2_X2 U524 ( .A1(n620), .A2(n708), .ZN(n622) );
  NAND2_X1 U525 ( .A1(n440), .A2(n437), .ZN(n413) );
  NOR2_X2 U526 ( .A1(n625), .A2(n708), .ZN(n627) );
  NAND2_X1 U527 ( .A1(n388), .A2(n357), .ZN(n399) );
  INV_X1 U528 ( .A(n709), .ZN(n388) );
  XNOR2_X1 U529 ( .A(n389), .B(KEYINPUT60), .ZN(G60) );
  NOR2_X2 U530 ( .A1(n703), .A2(n708), .ZN(n389) );
  AND2_X1 U531 ( .A1(n392), .A2(n391), .ZN(G54) );
  XNOR2_X1 U532 ( .A(n696), .B(n697), .ZN(n392) );
  XNOR2_X1 U533 ( .A(n424), .B(n366), .ZN(n570) );
  NAND2_X1 U534 ( .A1(n553), .A2(n600), .ZN(n562) );
  XNOR2_X1 U535 ( .A(n593), .B(KEYINPUT35), .ZN(n733) );
  NAND2_X1 U536 ( .A1(n670), .A2(n359), .ZN(n420) );
  XNOR2_X2 U537 ( .A(G125), .B(G146), .ZN(n474) );
  NAND2_X1 U538 ( .A1(n363), .A2(n652), .ZN(n722) );
  NAND2_X1 U539 ( .A1(n709), .A2(n416), .ZN(n402) );
  INV_X1 U540 ( .A(n496), .ZN(n404) );
  NAND2_X1 U541 ( .A1(n735), .A2(n547), .ZN(n406) );
  NAND2_X1 U542 ( .A1(n559), .A2(n558), .ZN(n650) );
  NAND2_X1 U543 ( .A1(n541), .A2(n359), .ZN(n411) );
  XNOR2_X1 U544 ( .A(n413), .B(G110), .ZN(G12) );
  NAND2_X1 U545 ( .A1(n419), .A2(n363), .ZN(n418) );
  NOR2_X1 U546 ( .A1(n709), .A2(n361), .ZN(n419) );
  XNOR2_X1 U547 ( .A(n421), .B(n431), .ZN(n430) );
  INV_X1 U548 ( .A(n527), .ZN(n580) );
  INV_X1 U549 ( .A(n436), .ZN(n439) );
  NAND2_X1 U550 ( .A1(n436), .A2(n364), .ZN(n443) );
  NAND2_X1 U551 ( .A1(n577), .A2(n576), .ZN(n446) );
  XNOR2_X1 U552 ( .A(n690), .B(n689), .ZN(n691) );
  XOR2_X1 U553 ( .A(n499), .B(n498), .Z(n447) );
  INV_X1 U554 ( .A(KEYINPUT48), .ZN(n561) );
  XNOR2_X1 U555 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U556 ( .A(n470), .B(KEYINPUT12), .ZN(n456) );
  XNOR2_X1 U557 ( .A(n688), .B(n687), .ZN(n689) );
  XNOR2_X1 U558 ( .A(n535), .B(n534), .ZN(n571) );
  XNOR2_X1 U559 ( .A(KEYINPUT63), .B(KEYINPUT89), .ZN(n626) );
  INV_X1 U560 ( .A(KEYINPUT121), .ZN(n621) );
  XOR2_X2 U561 ( .A(KEYINPUT64), .B(G953), .Z(n476) );
  XOR2_X1 U562 ( .A(KEYINPUT42), .B(KEYINPUT106), .Z(n526) );
  XOR2_X1 U563 ( .A(G131), .B(G113), .Z(n450) );
  XNOR2_X1 U564 ( .A(n450), .B(n449), .ZN(n454) );
  XNOR2_X1 U565 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U566 ( .A(n455), .B(KEYINPUT70), .ZN(n488) );
  NOR2_X1 U567 ( .A1(G902), .A2(n700), .ZN(n459) );
  XNOR2_X1 U568 ( .A(KEYINPUT13), .B(G475), .ZN(n458) );
  XNOR2_X1 U569 ( .A(n459), .B(n458), .ZN(n537) );
  INV_X1 U570 ( .A(n537), .ZN(n539) );
  XOR2_X1 U571 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n462) );
  INV_X1 U572 ( .A(n471), .ZN(n460) );
  XNOR2_X1 U573 ( .A(n475), .B(n460), .ZN(n461) );
  XNOR2_X1 U574 ( .A(n462), .B(n461), .ZN(n466) );
  XOR2_X1 U575 ( .A(G122), .B(G134), .Z(n465) );
  NAND2_X1 U576 ( .A1(G217), .A2(n463), .ZN(n464) );
  NOR2_X1 U577 ( .A1(G902), .A2(n704), .ZN(n468) );
  XNOR2_X1 U578 ( .A(KEYINPUT96), .B(G478), .ZN(n467) );
  XNOR2_X1 U579 ( .A(n468), .B(n467), .ZN(n540) );
  NAND2_X1 U580 ( .A1(n539), .A2(n540), .ZN(n469) );
  XNOR2_X1 U581 ( .A(n469), .B(KEYINPUT98), .ZN(n578) );
  XNOR2_X1 U582 ( .A(n473), .B(n472), .ZN(n491) );
  NAND2_X1 U583 ( .A1(G224), .A2(n476), .ZN(n477) );
  NAND2_X1 U584 ( .A1(G210), .A2(n481), .ZN(n479) );
  INV_X1 U585 ( .A(n568), .ZN(n544) );
  NOR2_X1 U586 ( .A1(n578), .A2(n667), .ZN(n674) );
  NAND2_X1 U587 ( .A1(G214), .A2(n481), .ZN(n482) );
  XNOR2_X1 U588 ( .A(KEYINPUT90), .B(n482), .ZN(n563) );
  NAND2_X1 U589 ( .A1(n674), .A2(n563), .ZN(n483) );
  XNOR2_X1 U590 ( .A(G131), .B(G134), .ZN(n484) );
  XNOR2_X1 U591 ( .A(n487), .B(n486), .ZN(n490) );
  NAND2_X1 U592 ( .A1(n488), .A2(G210), .ZN(n489) );
  XOR2_X1 U593 ( .A(n490), .B(n489), .Z(n492) );
  NOR2_X1 U594 ( .A1(G902), .A2(n623), .ZN(n495) );
  XNOR2_X1 U595 ( .A(KEYINPUT94), .B(G472), .ZN(n494) );
  NOR2_X1 U596 ( .A1(G902), .A2(n619), .ZN(n500) );
  XOR2_X1 U597 ( .A(KEYINPUT92), .B(KEYINPUT25), .Z(n499) );
  INV_X1 U598 ( .A(n616), .ZN(n496) );
  NAND2_X1 U599 ( .A1(n496), .A2(G234), .ZN(n497) );
  XNOR2_X1 U600 ( .A(n497), .B(KEYINPUT20), .ZN(n501) );
  NAND2_X1 U601 ( .A1(n501), .A2(G217), .ZN(n498) );
  XOR2_X1 U602 ( .A(KEYINPUT93), .B(KEYINPUT21), .Z(n503) );
  NAND2_X1 U603 ( .A1(n501), .A2(G221), .ZN(n502) );
  NAND2_X1 U604 ( .A1(G237), .A2(G234), .ZN(n504) );
  XNOR2_X1 U605 ( .A(n504), .B(KEYINPUT14), .ZN(n505) );
  AND2_X1 U606 ( .A1(G952), .A2(n505), .ZN(n680) );
  NAND2_X1 U607 ( .A1(n572), .A2(n680), .ZN(n574) );
  INV_X1 U608 ( .A(n574), .ZN(n510) );
  INV_X1 U609 ( .A(n476), .ZN(n507) );
  NAND2_X1 U610 ( .A1(n505), .A2(G902), .ZN(n506) );
  XNOR2_X1 U611 ( .A(n506), .B(KEYINPUT91), .ZN(n573) );
  NAND2_X1 U612 ( .A1(n507), .A2(n573), .ZN(n508) );
  NOR2_X1 U613 ( .A1(G900), .A2(n508), .ZN(n509) );
  NOR2_X1 U614 ( .A1(n510), .A2(n509), .ZN(n511) );
  XNOR2_X1 U615 ( .A(KEYINPUT75), .B(n511), .ZN(n541) );
  NAND2_X1 U616 ( .A1(G227), .A2(n476), .ZN(n512) );
  XOR2_X1 U617 ( .A(n513), .B(n512), .Z(n520) );
  INV_X1 U618 ( .A(n514), .ZN(n515) );
  XNOR2_X1 U619 ( .A(n515), .B(G110), .ZN(n517) );
  NOR2_X1 U620 ( .A1(n693), .A2(G902), .ZN(n522) );
  XNOR2_X2 U621 ( .A(n522), .B(n521), .ZN(n557) );
  XNOR2_X1 U622 ( .A(n557), .B(KEYINPUT105), .ZN(n523) );
  NOR2_X1 U623 ( .A1(n524), .A2(n523), .ZN(n549) );
  NAND2_X1 U624 ( .A1(n666), .A2(n549), .ZN(n525) );
  XNOR2_X1 U625 ( .A(n526), .B(n525), .ZN(n731) );
  NAND2_X1 U626 ( .A1(n537), .A2(n540), .ZN(n643) );
  XNOR2_X1 U627 ( .A(KEYINPUT103), .B(KEYINPUT30), .ZN(n529) );
  INV_X1 U628 ( .A(n563), .ZN(n672) );
  NOR2_X1 U629 ( .A1(n672), .A2(n356), .ZN(n528) );
  XNOR2_X1 U630 ( .A(n529), .B(n528), .ZN(n530) );
  NOR2_X1 U631 ( .A1(n531), .A2(n530), .ZN(n542) );
  INV_X1 U632 ( .A(n541), .ZN(n532) );
  NOR2_X1 U633 ( .A1(n667), .A2(n532), .ZN(n533) );
  AND2_X1 U634 ( .A1(n542), .A2(n533), .ZN(n535) );
  OR2_X1 U635 ( .A1(n537), .A2(n540), .ZN(n646) );
  NAND2_X1 U636 ( .A1(n643), .A2(n646), .ZN(n607) );
  INV_X1 U637 ( .A(n607), .ZN(n668) );
  NAND2_X1 U638 ( .A1(KEYINPUT47), .A2(n668), .ZN(n538) );
  XNOR2_X1 U639 ( .A(KEYINPUT78), .B(n538), .ZN(n547) );
  NOR2_X1 U640 ( .A1(n540), .A2(n539), .ZN(n590) );
  NAND2_X1 U641 ( .A1(n542), .A2(n541), .ZN(n543) );
  NOR2_X1 U642 ( .A1(n544), .A2(n543), .ZN(n545) );
  NAND2_X1 U643 ( .A1(n590), .A2(n545), .ZN(n546) );
  NOR2_X1 U644 ( .A1(KEYINPUT47), .A2(n668), .ZN(n548) );
  XNOR2_X1 U645 ( .A(KEYINPUT69), .B(n548), .ZN(n551) );
  NAND2_X1 U646 ( .A1(n549), .A2(n577), .ZN(n550) );
  NOR2_X1 U647 ( .A1(n643), .A2(n552), .ZN(n553) );
  NOR2_X1 U648 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U649 ( .A(KEYINPUT36), .B(n556), .ZN(n559) );
  XNOR2_X2 U650 ( .A(n557), .B(KEYINPUT1), .ZN(n587) );
  XNOR2_X1 U651 ( .A(n587), .B(KEYINPUT87), .ZN(n581) );
  INV_X1 U652 ( .A(n581), .ZN(n558) );
  NAND2_X1 U653 ( .A1(n641), .A2(KEYINPUT47), .ZN(n560) );
  XOR2_X1 U654 ( .A(KEYINPUT100), .B(KEYINPUT43), .Z(n566) );
  NOR2_X1 U655 ( .A1(n587), .A2(n562), .ZN(n564) );
  NAND2_X1 U656 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U657 ( .A(n566), .B(n565), .ZN(n567) );
  NOR2_X1 U658 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U659 ( .A(KEYINPUT101), .B(n569), .ZN(n732) );
  OR2_X1 U660 ( .A1(n646), .A2(n571), .ZN(n652) );
  NOR2_X1 U661 ( .A1(G898), .A2(n572), .ZN(n716) );
  NAND2_X1 U662 ( .A1(n716), .A2(n573), .ZN(n575) );
  NAND2_X1 U663 ( .A1(n575), .A2(n574), .ZN(n576) );
  INV_X1 U664 ( .A(n578), .ZN(n670) );
  INV_X1 U665 ( .A(n587), .ZN(n597) );
  AND2_X1 U666 ( .A1(n356), .A2(n597), .ZN(n579) );
  XNOR2_X1 U667 ( .A(KEYINPUT99), .B(n580), .ZN(n656) );
  NOR2_X1 U668 ( .A1(n581), .A2(n656), .ZN(n582) );
  NOR2_X1 U669 ( .A1(KEYINPUT44), .A2(KEYINPUT83), .ZN(n583) );
  XNOR2_X1 U670 ( .A(n585), .B(n584), .ZN(n594) );
  XNOR2_X1 U671 ( .A(KEYINPUT34), .B(KEYINPUT72), .ZN(n586) );
  INV_X1 U672 ( .A(n605), .ZN(n602) );
  NAND2_X1 U673 ( .A1(n653), .A2(n587), .ZN(n601) );
  XNOR2_X1 U674 ( .A(KEYINPUT85), .B(KEYINPUT33), .ZN(n589) );
  INV_X1 U675 ( .A(n590), .ZN(n591) );
  NAND2_X1 U676 ( .A1(n594), .A2(n733), .ZN(n596) );
  NAND2_X1 U677 ( .A1(n596), .A2(n595), .ZN(n612) );
  AND2_X1 U678 ( .A1(n436), .A2(n597), .ZN(n598) );
  NAND2_X1 U679 ( .A1(n656), .A2(n598), .ZN(n599) );
  NOR2_X1 U680 ( .A1(n600), .A2(n599), .ZN(n628) );
  NOR2_X1 U681 ( .A1(n356), .A2(n601), .ZN(n663) );
  NAND2_X1 U682 ( .A1(n602), .A2(n663), .ZN(n603) );
  XOR2_X1 U683 ( .A(KEYINPUT31), .B(n603), .Z(n645) );
  NOR2_X1 U684 ( .A1(n605), .A2(n604), .ZN(n606) );
  NAND2_X1 U685 ( .A1(n356), .A2(n606), .ZN(n633) );
  NAND2_X1 U686 ( .A1(n645), .A2(n633), .ZN(n608) );
  NAND2_X1 U687 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U688 ( .A(n609), .B(KEYINPUT97), .ZN(n610) );
  NOR2_X1 U689 ( .A1(n628), .A2(n610), .ZN(n611) );
  NAND2_X1 U690 ( .A1(n612), .A2(n611), .ZN(n615) );
  INV_X1 U691 ( .A(KEYINPUT45), .ZN(n613) );
  NAND2_X1 U692 ( .A1(KEYINPUT2), .A2(n652), .ZN(n617) );
  XNOR2_X1 U693 ( .A(n618), .B(n619), .ZN(n620) );
  XNOR2_X1 U694 ( .A(n622), .B(n621), .ZN(G66) );
  XNOR2_X1 U695 ( .A(n627), .B(n626), .ZN(G57) );
  XOR2_X1 U696 ( .A(G101), .B(n628), .Z(n629) );
  XNOR2_X1 U697 ( .A(KEYINPUT108), .B(n629), .ZN(G3) );
  NOR2_X1 U698 ( .A1(n643), .A2(n633), .ZN(n630) );
  XOR2_X1 U699 ( .A(G104), .B(n630), .Z(G6) );
  XOR2_X1 U700 ( .A(KEYINPUT111), .B(KEYINPUT110), .Z(n632) );
  XNOR2_X1 U701 ( .A(KEYINPUT26), .B(KEYINPUT27), .ZN(n631) );
  XNOR2_X1 U702 ( .A(n632), .B(n631), .ZN(n637) );
  NOR2_X1 U703 ( .A1(n646), .A2(n633), .ZN(n635) );
  XNOR2_X1 U704 ( .A(G107), .B(KEYINPUT109), .ZN(n634) );
  XNOR2_X1 U705 ( .A(n635), .B(n634), .ZN(n636) );
  XOR2_X1 U706 ( .A(n637), .B(n636), .Z(G9) );
  NOR2_X1 U707 ( .A1(n641), .A2(n646), .ZN(n639) );
  XNOR2_X1 U708 ( .A(KEYINPUT112), .B(KEYINPUT29), .ZN(n638) );
  XNOR2_X1 U709 ( .A(n639), .B(n638), .ZN(n640) );
  XNOR2_X1 U710 ( .A(G128), .B(n640), .ZN(G30) );
  NOR2_X1 U711 ( .A1(n641), .A2(n643), .ZN(n642) );
  XOR2_X1 U712 ( .A(G146), .B(n642), .Z(G48) );
  NOR2_X1 U713 ( .A1(n643), .A2(n645), .ZN(n644) );
  XOR2_X1 U714 ( .A(G113), .B(n644), .Z(G15) );
  NOR2_X1 U715 ( .A1(n646), .A2(n645), .ZN(n647) );
  XOR2_X1 U716 ( .A(KEYINPUT114), .B(n647), .Z(n648) );
  XNOR2_X1 U717 ( .A(G116), .B(n648), .ZN(G18) );
  XOR2_X1 U718 ( .A(G125), .B(KEYINPUT37), .Z(n649) );
  XNOR2_X1 U719 ( .A(n650), .B(n649), .ZN(G27) );
  XOR2_X1 U720 ( .A(G134), .B(KEYINPUT115), .Z(n651) );
  XNOR2_X1 U721 ( .A(n652), .B(n651), .ZN(G36) );
  NAND2_X1 U722 ( .A1(n676), .A2(n666), .ZN(n683) );
  XOR2_X1 U723 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n655) );
  OR2_X1 U724 ( .A1(n587), .A2(n653), .ZN(n654) );
  XNOR2_X1 U725 ( .A(n655), .B(n654), .ZN(n661) );
  NOR2_X1 U726 ( .A1(n656), .A2(n359), .ZN(n657) );
  XNOR2_X1 U727 ( .A(KEYINPUT49), .B(n657), .ZN(n659) );
  NAND2_X1 U728 ( .A1(n659), .A2(n356), .ZN(n660) );
  NOR2_X1 U729 ( .A1(n661), .A2(n660), .ZN(n662) );
  NOR2_X1 U730 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U731 ( .A(KEYINPUT51), .B(n664), .ZN(n665) );
  NAND2_X1 U732 ( .A1(n666), .A2(n665), .ZN(n678) );
  NOR2_X1 U733 ( .A1(n668), .A2(n667), .ZN(n669) );
  NOR2_X1 U734 ( .A1(n670), .A2(n669), .ZN(n671) );
  NOR2_X1 U735 ( .A1(n672), .A2(n671), .ZN(n673) );
  OR2_X1 U736 ( .A1(n674), .A2(n673), .ZN(n675) );
  NAND2_X1 U737 ( .A1(n676), .A2(n675), .ZN(n677) );
  NAND2_X1 U738 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U739 ( .A(KEYINPUT52), .B(n679), .ZN(n681) );
  NAND2_X1 U740 ( .A1(n681), .A2(n680), .ZN(n682) );
  NAND2_X1 U741 ( .A1(n683), .A2(n682), .ZN(n684) );
  XOR2_X1 U742 ( .A(KEYINPUT117), .B(n684), .Z(n685) );
  NAND2_X1 U743 ( .A1(n698), .A2(G210), .ZN(n690) );
  XOR2_X1 U744 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n687) );
  XNOR2_X1 U745 ( .A(n692), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U746 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n695) );
  XNOR2_X1 U747 ( .A(n693), .B(KEYINPUT119), .ZN(n694) );
  XNOR2_X1 U748 ( .A(n695), .B(n694), .ZN(n697) );
  NAND2_X1 U749 ( .A1(n698), .A2(G469), .ZN(n696) );
  NAND2_X1 U750 ( .A1(n698), .A2(G475), .ZN(n702) );
  XOR2_X1 U751 ( .A(KEYINPUT59), .B(KEYINPUT88), .Z(n699) );
  XNOR2_X1 U752 ( .A(n700), .B(n699), .ZN(n701) );
  XNOR2_X1 U753 ( .A(n702), .B(n701), .ZN(n703) );
  XNOR2_X1 U754 ( .A(n704), .B(KEYINPUT120), .ZN(n706) );
  NAND2_X1 U755 ( .A1(G478), .A2(n698), .ZN(n705) );
  XNOR2_X1 U756 ( .A(n706), .B(n705), .ZN(n707) );
  NOR2_X1 U757 ( .A1(n708), .A2(n707), .ZN(G63) );
  OR2_X1 U758 ( .A1(G953), .A2(n709), .ZN(n714) );
  NAND2_X1 U759 ( .A1(G224), .A2(G953), .ZN(n710) );
  XNOR2_X1 U760 ( .A(n710), .B(KEYINPUT122), .ZN(n711) );
  XNOR2_X1 U761 ( .A(KEYINPUT61), .B(n711), .ZN(n712) );
  NAND2_X1 U762 ( .A1(n712), .A2(G898), .ZN(n713) );
  NAND2_X1 U763 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U764 ( .A(n715), .B(KEYINPUT123), .ZN(n717) );
  XOR2_X1 U765 ( .A(n717), .B(n369), .Z(G69) );
  XOR2_X1 U766 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n719) );
  XNOR2_X1 U767 ( .A(n718), .B(n719), .ZN(n720) );
  XNOR2_X1 U768 ( .A(n721), .B(n720), .ZN(n724) );
  XNOR2_X1 U769 ( .A(n722), .B(n724), .ZN(n723) );
  NAND2_X1 U770 ( .A1(n723), .A2(n476), .ZN(n730) );
  XNOR2_X1 U771 ( .A(n724), .B(G227), .ZN(n725) );
  XNOR2_X1 U772 ( .A(n725), .B(KEYINPUT126), .ZN(n726) );
  NAND2_X1 U773 ( .A1(n726), .A2(G900), .ZN(n727) );
  NAND2_X1 U774 ( .A1(G953), .A2(n727), .ZN(n728) );
  XOR2_X1 U775 ( .A(KEYINPUT127), .B(n728), .Z(n729) );
  NAND2_X1 U776 ( .A1(n730), .A2(n729), .ZN(G72) );
  XOR2_X1 U777 ( .A(n731), .B(G137), .Z(G39) );
  XNOR2_X1 U778 ( .A(G140), .B(n732), .ZN(G42) );
  XNOR2_X1 U779 ( .A(n733), .B(G122), .ZN(G24) );
  XOR2_X1 U780 ( .A(G131), .B(n734), .Z(G33) );
  XOR2_X1 U781 ( .A(G143), .B(n735), .Z(n736) );
  XNOR2_X1 U782 ( .A(KEYINPUT113), .B(n736), .ZN(G45) );
  XNOR2_X1 U783 ( .A(n737), .B(G119), .ZN(G21) );
endmodule

