//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 1 1 1 1 1 1 1 1 0 0 0 1 1 0 1 0 0 0 1 0 0 0 0 1 1 0 0 0 0 0 1 0 0 1 1 0 0 1 1 0 1 1 0 0 1 1 1 0 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:35 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n748, new_n749, new_n751, new_n752, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013;
  INV_X1    g000(.A(KEYINPUT85), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT12), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT64), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n189), .B1(new_n190), .B2(G146), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(KEYINPUT64), .A3(G143), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n190), .A2(G146), .ZN(new_n194));
  NAND4_X1  g008(.A1(new_n191), .A2(new_n193), .A3(G128), .A4(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT1), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(KEYINPUT66), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT66), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(KEYINPUT1), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n195), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT67), .ZN(new_n202));
  XNOR2_X1  g016(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n190), .A2(G146), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n202), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n192), .A2(G143), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n200), .A2(KEYINPUT67), .A3(new_n206), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n205), .A2(new_n207), .A3(G128), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n194), .A2(new_n206), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n201), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G107), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n211), .A2(G104), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT3), .ZN(new_n213));
  INV_X1    g027(.A(G104), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n214), .A2(G107), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n212), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G101), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT79), .ZN(new_n218));
  OAI211_X1 g032(.A(new_n218), .B(KEYINPUT3), .C1(new_n214), .C2(G107), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n211), .A2(G104), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n218), .B1(new_n221), .B2(KEYINPUT3), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n216), .B(new_n217), .C1(new_n220), .C2(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(G101), .B1(new_n215), .B2(new_n212), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n210), .A2(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n191), .A2(new_n194), .A3(new_n193), .ZN(new_n227));
  OAI21_X1  g041(.A(G128), .B1(new_n204), .B2(new_n196), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT80), .ZN(new_n230));
  OAI22_X1  g044(.A1(new_n229), .A2(new_n230), .B1(new_n195), .B2(new_n200), .ZN(new_n231));
  AOI21_X1  g045(.A(KEYINPUT80), .B1(new_n227), .B2(new_n228), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n223), .B(new_n224), .C1(new_n231), .C2(new_n232), .ZN(new_n233));
  AND2_X1   g047(.A1(new_n226), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(G131), .ZN(new_n235));
  INV_X1    g049(.A(G137), .ZN(new_n236));
  OAI21_X1  g050(.A(KEYINPUT65), .B1(new_n236), .B2(G134), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT65), .ZN(new_n238));
  INV_X1    g052(.A(G134), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n238), .A2(new_n239), .A3(G137), .ZN(new_n240));
  AND2_X1   g054(.A1(new_n237), .A2(new_n240), .ZN(new_n241));
  AND3_X1   g055(.A1(new_n236), .A2(KEYINPUT11), .A3(G134), .ZN(new_n242));
  AOI21_X1  g056(.A(KEYINPUT11), .B1(new_n236), .B2(G134), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n235), .B1(new_n241), .B2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT11), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n246), .B1(new_n239), .B2(G137), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n236), .A2(KEYINPUT11), .A3(G134), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n237), .A2(new_n247), .A3(new_n240), .A4(new_n248), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n249), .A2(G131), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n245), .A2(new_n250), .ZN(new_n251));
  OAI211_X1 g065(.A(KEYINPUT84), .B(new_n188), .C1(new_n234), .C2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT84), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n251), .B1(new_n226), .B2(new_n233), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n253), .B1(new_n254), .B2(KEYINPUT12), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(KEYINPUT12), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n252), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT10), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n233), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n195), .ZN(new_n260));
  XOR2_X1   g074(.A(KEYINPUT0), .B(G128), .Z(new_n261));
  AOI22_X1  g075(.A1(new_n260), .A2(KEYINPUT0), .B1(new_n209), .B2(new_n261), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n216), .B1(new_n220), .B2(new_n222), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n263), .A2(new_n264), .A3(G101), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n223), .A2(KEYINPUT4), .ZN(new_n266));
  OAI21_X1  g080(.A(KEYINPUT79), .B1(new_n215), .B2(new_n213), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(new_n219), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n217), .B1(new_n268), .B2(new_n216), .ZN(new_n269));
  OAI211_X1 g083(.A(new_n262), .B(new_n265), .C1(new_n266), .C2(new_n269), .ZN(new_n270));
  AND2_X1   g084(.A1(new_n259), .A2(new_n270), .ZN(new_n271));
  XOR2_X1   g085(.A(new_n251), .B(KEYINPUT83), .Z(new_n272));
  INV_X1    g086(.A(KEYINPUT81), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n225), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n223), .A2(KEYINPUT81), .A3(new_n224), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(G128), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n198), .A2(KEYINPUT1), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n196), .A2(KEYINPUT66), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n206), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n277), .B1(new_n280), .B2(new_n202), .ZN(new_n281));
  AOI22_X1  g095(.A1(new_n281), .A2(new_n207), .B1(new_n194), .B2(new_n206), .ZN(new_n282));
  OAI21_X1  g096(.A(KEYINPUT10), .B1(new_n282), .B2(new_n201), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT82), .ZN(new_n284));
  NOR3_X1   g098(.A1(new_n276), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(new_n275), .ZN(new_n286));
  AOI21_X1  g100(.A(KEYINPUT81), .B1(new_n223), .B2(new_n224), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n210), .A2(new_n258), .ZN(new_n289));
  AOI21_X1  g103(.A(KEYINPUT82), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n271), .B(new_n272), .C1(new_n285), .C2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n257), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g106(.A(G110), .B(G140), .ZN(new_n293));
  INV_X1    g107(.A(G227), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n294), .A2(G953), .ZN(new_n295));
  XOR2_X1   g109(.A(new_n293), .B(new_n295), .Z(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n229), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n201), .B1(new_n298), .B2(KEYINPUT80), .ZN(new_n299));
  INV_X1    g113(.A(new_n232), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n225), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n270), .B1(new_n301), .B2(KEYINPUT10), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n284), .B1(new_n276), .B2(new_n283), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n288), .A2(new_n289), .A3(KEYINPUT82), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n297), .B1(new_n305), .B2(new_n272), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n271), .B1(new_n285), .B2(new_n290), .ZN(new_n307));
  INV_X1    g121(.A(new_n251), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  AOI22_X1  g123(.A1(new_n292), .A2(new_n297), .B1(new_n306), .B2(new_n309), .ZN(new_n310));
  OAI211_X1 g124(.A(new_n187), .B(G469), .C1(new_n310), .C2(G902), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G902), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n303), .A2(new_n304), .ZN(new_n314));
  AND3_X1   g128(.A1(new_n314), .A2(new_n271), .A3(new_n272), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n251), .B1(new_n314), .B2(new_n271), .ZN(new_n316));
  NOR3_X1   g130(.A1(new_n315), .A2(new_n316), .A3(new_n297), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n296), .B1(new_n257), .B2(new_n291), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n313), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n187), .B1(new_n319), .B2(G469), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n297), .B1(new_n315), .B2(new_n316), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n306), .A2(new_n257), .ZN(new_n322));
  AOI21_X1  g136(.A(G902), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(G469), .ZN(new_n324));
  AOI21_X1  g138(.A(KEYINPUT86), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n291), .B1(new_n251), .B2(new_n305), .ZN(new_n326));
  AOI22_X1  g140(.A1(new_n326), .A2(new_n297), .B1(new_n306), .B2(new_n257), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT86), .ZN(new_n328));
  NOR4_X1   g142(.A1(new_n327), .A2(new_n328), .A3(G469), .A4(G902), .ZN(new_n329));
  OAI22_X1  g143(.A1(new_n312), .A2(new_n320), .B1(new_n325), .B2(new_n329), .ZN(new_n330));
  OAI21_X1  g144(.A(G214), .B1(G237), .B2(G902), .ZN(new_n331));
  INV_X1    g145(.A(G116), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(KEYINPUT69), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT69), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(G116), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n333), .A2(new_n335), .A3(G119), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n336), .B1(new_n332), .B2(G119), .ZN(new_n337));
  XNOR2_X1  g151(.A(KEYINPUT2), .B(G113), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n338), .ZN(new_n340));
  OAI211_X1 g154(.A(new_n340), .B(new_n336), .C1(new_n332), .C2(G119), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n342), .B(new_n265), .C1(new_n266), .C2(new_n269), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT87), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n263), .A2(G101), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n346), .A2(KEYINPUT4), .A3(new_n223), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n347), .A2(KEYINPUT87), .A3(new_n342), .A4(new_n265), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n332), .A2(G119), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT5), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  OAI211_X1 g165(.A(G113), .B(new_n351), .C1(new_n337), .C2(new_n350), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n274), .A2(new_n341), .A3(new_n275), .A4(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n345), .A2(new_n348), .A3(new_n353), .ZN(new_n354));
  XNOR2_X1  g168(.A(G110), .B(G122), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n345), .A2(new_n353), .A3(new_n348), .A4(new_n355), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n357), .A2(KEYINPUT6), .A3(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT6), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n354), .A2(new_n360), .A3(new_n356), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n262), .A2(G125), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n362), .B1(new_n210), .B2(G125), .ZN(new_n363));
  INV_X1    g177(.A(G953), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(G224), .ZN(new_n365));
  XNOR2_X1  g179(.A(new_n363), .B(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n359), .A2(new_n361), .A3(new_n366), .ZN(new_n367));
  XNOR2_X1  g181(.A(new_n355), .B(KEYINPUT8), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n352), .A2(new_n341), .ZN(new_n369));
  AND2_X1   g183(.A1(new_n369), .A2(new_n225), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n369), .A2(new_n225), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n368), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  AND2_X1   g186(.A1(new_n365), .A2(KEYINPUT7), .ZN(new_n373));
  OR2_X1    g187(.A1(new_n363), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n363), .A2(new_n373), .ZN(new_n375));
  AND3_X1   g189(.A1(new_n372), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(G902), .B1(new_n376), .B2(new_n358), .ZN(new_n377));
  OAI21_X1  g191(.A(G210), .B1(G237), .B2(G902), .ZN(new_n378));
  AND3_X1   g192(.A1(new_n367), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n378), .B(KEYINPUT88), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n381), .B1(new_n367), .B2(new_n377), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n331), .B1(new_n379), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(KEYINPUT89), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n367), .A2(new_n377), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(new_n380), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n367), .A2(new_n377), .A3(new_n378), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT89), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n388), .A2(new_n389), .A3(new_n331), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n384), .A2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(G221), .ZN(new_n392));
  XNOR2_X1  g206(.A(KEYINPUT9), .B(G234), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n392), .B1(new_n394), .B2(new_n313), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  NOR2_X1   g210(.A1(G475), .A2(G902), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT92), .ZN(new_n399));
  INV_X1    g213(.A(G125), .ZN(new_n400));
  OAI21_X1  g214(.A(KEYINPUT76), .B1(new_n400), .B2(G140), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT76), .ZN(new_n402));
  INV_X1    g216(.A(G140), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n402), .A2(new_n403), .A3(G125), .ZN(new_n404));
  AOI21_X1  g218(.A(KEYINPUT16), .B1(new_n401), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(KEYINPUT76), .A2(KEYINPUT16), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n403), .A2(G125), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n400), .A2(G140), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n406), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  OAI21_X1  g223(.A(G146), .B1(new_n405), .B2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT77), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  OR2_X1    g226(.A1(KEYINPUT90), .A2(G143), .ZN(new_n413));
  NOR2_X1   g227(.A1(G237), .A2(G953), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n413), .B1(G214), .B2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(G237), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n416), .A2(new_n364), .A3(G214), .ZN(new_n417));
  NOR2_X1   g231(.A1(KEYINPUT90), .A2(G143), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(G131), .B1(new_n415), .B2(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n413), .A2(G214), .A3(new_n414), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n417), .A2(new_n418), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n421), .A2(new_n422), .A3(new_n235), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n420), .A2(new_n423), .ZN(new_n424));
  OAI211_X1 g238(.A(KEYINPUT77), .B(G146), .C1(new_n405), .C2(new_n409), .ZN(new_n425));
  AND3_X1   g239(.A1(new_n407), .A2(new_n408), .A3(KEYINPUT19), .ZN(new_n426));
  AOI21_X1  g240(.A(KEYINPUT19), .B1(new_n407), .B2(new_n408), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n192), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n412), .A2(new_n424), .A3(new_n425), .A4(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n421), .A2(new_n422), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n430), .A2(KEYINPUT18), .A3(G131), .ZN(new_n431));
  NAND2_X1  g245(.A1(KEYINPUT18), .A2(G131), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n421), .A2(new_n422), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n407), .A2(new_n408), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(G146), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT91), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n407), .A2(new_n408), .A3(new_n192), .ZN(new_n437));
  AND3_X1   g251(.A1(new_n435), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n436), .B1(new_n435), .B2(new_n437), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n431), .B(new_n433), .C1(new_n438), .C2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n429), .A2(new_n440), .ZN(new_n441));
  XNOR2_X1  g255(.A(G113), .B(G122), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n442), .B(new_n214), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n399), .B1(new_n441), .B2(new_n444), .ZN(new_n445));
  AOI211_X1 g259(.A(KEYINPUT92), .B(new_n443), .C1(new_n429), .C2(new_n440), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n401), .A2(new_n404), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT16), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(new_n409), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n450), .A2(new_n451), .A3(new_n192), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(new_n410), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT17), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n420), .A2(new_n454), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(KEYINPUT93), .B1(new_n424), .B2(KEYINPUT17), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT93), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n420), .A2(new_n458), .A3(new_n454), .A4(new_n423), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n456), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n460), .A2(new_n443), .A3(new_n440), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n398), .B1(new_n447), .B2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT20), .ZN(new_n463));
  OAI21_X1  g277(.A(KEYINPUT94), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n441), .A2(new_n444), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(KEYINPUT92), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n441), .A2(new_n399), .A3(new_n444), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n466), .A2(new_n461), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(new_n397), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT94), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n469), .A2(new_n470), .A3(KEYINPUT20), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n462), .A2(new_n463), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n464), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n461), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n443), .B1(new_n460), .B2(new_n440), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n313), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(G475), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n473), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(G478), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n479), .A2(KEYINPUT15), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n190), .A2(G128), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n277), .A2(G143), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(G134), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n481), .A2(new_n482), .A3(new_n239), .ZN(new_n485));
  AND3_X1   g299(.A1(new_n484), .A2(KEYINPUT97), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(KEYINPUT97), .B1(new_n484), .B2(new_n485), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n333), .A2(new_n335), .A3(G122), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT95), .ZN(new_n490));
  OR2_X1    g304(.A1(new_n332), .A2(G122), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n489), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n490), .B1(new_n489), .B2(new_n491), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n211), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  AND2_X1   g309(.A1(new_n489), .A2(KEYINPUT14), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n491), .B1(new_n489), .B2(KEYINPUT14), .ZN(new_n497));
  OAI21_X1  g311(.A(G107), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  AND3_X1   g312(.A1(new_n488), .A2(new_n495), .A3(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT13), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n481), .A2(KEYINPUT96), .A3(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n190), .A2(KEYINPUT13), .A3(G128), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n501), .A2(new_n482), .A3(new_n502), .ZN(new_n503));
  AOI21_X1  g317(.A(KEYINPUT96), .B1(new_n481), .B2(new_n500), .ZN(new_n504));
  OAI21_X1  g318(.A(G134), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n485), .ZN(new_n506));
  INV_X1    g320(.A(new_n494), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n507), .A2(G107), .A3(new_n492), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n506), .B1(new_n495), .B2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(G217), .ZN(new_n510));
  NOR3_X1   g324(.A1(new_n393), .A2(new_n510), .A3(G953), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  OR3_X1    g326(.A1(new_n499), .A2(new_n509), .A3(new_n512), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n512), .B1(new_n499), .B2(new_n509), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n480), .B1(new_n516), .B2(G902), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n515), .B(new_n313), .C1(KEYINPUT15), .C2(new_n479), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(G952), .ZN(new_n520));
  AOI211_X1 g334(.A(G953), .B(new_n520), .C1(G234), .C2(G237), .ZN(new_n521));
  INV_X1    g335(.A(G234), .ZN(new_n522));
  OAI211_X1 g336(.A(G902), .B(G953), .C1(new_n522), .C2(new_n416), .ZN(new_n523));
  XNOR2_X1  g337(.A(new_n523), .B(KEYINPUT98), .ZN(new_n524));
  XNOR2_X1  g338(.A(KEYINPUT21), .B(G898), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n521), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NOR3_X1   g340(.A1(new_n478), .A2(new_n519), .A3(new_n526), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n330), .A2(new_n391), .A3(new_n396), .A4(new_n527), .ZN(new_n528));
  XNOR2_X1  g342(.A(KEYINPUT68), .B(KEYINPUT30), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n241), .A2(new_n244), .A3(new_n235), .ZN(new_n531));
  XOR2_X1   g345(.A(G134), .B(G137), .Z(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(G131), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n535), .B1(new_n282), .B2(new_n201), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n261), .A2(new_n209), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n260), .A2(KEYINPUT0), .ZN(new_n538));
  OAI211_X1 g352(.A(new_n537), .B(new_n538), .C1(new_n245), .C2(new_n250), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n530), .B1(new_n536), .B2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT68), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n541), .A2(KEYINPUT30), .ZN(new_n542));
  OAI211_X1 g356(.A(new_n539), .B(new_n542), .C1(new_n210), .C2(new_n534), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n342), .B1(new_n540), .B2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT31), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n414), .A2(G210), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n547), .B(KEYINPUT27), .ZN(new_n548));
  XNOR2_X1  g362(.A(KEYINPUT26), .B(G101), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n548), .B(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n342), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n551), .B(new_n539), .C1(new_n210), .C2(new_n534), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n545), .A2(new_n546), .A3(new_n550), .A4(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT71), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n552), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n539), .B1(new_n210), .B2(new_n534), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(new_n529), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(new_n543), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n556), .B1(new_n559), .B2(new_n342), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n560), .A2(KEYINPUT71), .A3(new_n546), .A4(new_n550), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n555), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n560), .A2(new_n550), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n563), .A2(KEYINPUT70), .A3(KEYINPUT31), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT70), .ZN(new_n565));
  INV_X1    g379(.A(new_n550), .ZN(new_n566));
  AOI211_X1 g380(.A(new_n566), .B(new_n556), .C1(new_n559), .C2(new_n342), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n565), .B1(new_n567), .B2(new_n546), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n551), .B1(new_n536), .B2(new_n539), .ZN(new_n569));
  OAI21_X1  g383(.A(KEYINPUT28), .B1(new_n569), .B2(new_n556), .ZN(new_n570));
  OAI21_X1  g384(.A(KEYINPUT72), .B1(new_n556), .B2(KEYINPUT28), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT72), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT28), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n552), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n570), .A2(new_n571), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(new_n566), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n562), .A2(new_n564), .A3(new_n568), .A4(new_n576), .ZN(new_n577));
  NOR2_X1   g391(.A1(G472), .A2(G902), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT32), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n577), .A2(KEYINPUT32), .A3(new_n578), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n570), .A2(new_n571), .A3(new_n550), .A4(new_n574), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(G902), .B1(new_n584), .B2(KEYINPUT29), .ZN(new_n585));
  INV_X1    g399(.A(new_n560), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(new_n566), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT29), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT73), .ZN(new_n589));
  OAI211_X1 g403(.A(new_n587), .B(new_n588), .C1(new_n589), .C2(new_n583), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n584), .A2(KEYINPUT73), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n585), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(G472), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n581), .A2(new_n582), .A3(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n437), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n277), .A2(G119), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT23), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n277), .A2(KEYINPUT23), .A3(G119), .ZN(new_n599));
  INV_X1    g413(.A(G110), .ZN(new_n600));
  INV_X1    g414(.A(G119), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(G128), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n598), .A2(new_n599), .A3(new_n600), .A4(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n596), .A2(new_n602), .ZN(new_n604));
  XNOR2_X1  g418(.A(KEYINPUT24), .B(G110), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n595), .B1(new_n603), .B2(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n412), .A2(new_n425), .A3(new_n607), .ZN(new_n608));
  XOR2_X1   g422(.A(KEYINPUT24), .B(G110), .Z(new_n609));
  INV_X1    g423(.A(KEYINPUT75), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n609), .A2(new_n610), .A3(new_n596), .A4(new_n602), .ZN(new_n611));
  OAI21_X1  g425(.A(KEYINPUT75), .B1(new_n604), .B2(new_n605), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n598), .A2(new_n602), .A3(new_n599), .ZN(new_n613));
  AOI22_X1  g427(.A1(new_n611), .A2(new_n612), .B1(G110), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n453), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n608), .A2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT78), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(KEYINPUT22), .B(G137), .ZN(new_n619));
  NOR3_X1   g433(.A1(new_n392), .A2(new_n522), .A3(G953), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n608), .A2(new_n615), .A3(KEYINPUT78), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n618), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  OR2_X1    g437(.A1(new_n616), .A2(new_n621), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n623), .A2(new_n313), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(KEYINPUT25), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT25), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n623), .A2(new_n627), .A3(new_n313), .A4(new_n624), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n510), .B1(G234), .B2(new_n313), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(KEYINPUT74), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n626), .A2(new_n628), .A3(new_n630), .ZN(new_n631));
  AND2_X1   g445(.A1(new_n623), .A2(new_n624), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n630), .A2(G902), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n594), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n528), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(KEYINPUT99), .B(G101), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G3));
  OAI21_X1  g454(.A(G469), .B1(new_n310), .B2(G902), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(KEYINPUT85), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n311), .ZN(new_n643));
  AND2_X1   g457(.A1(new_n306), .A2(new_n257), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n296), .B1(new_n309), .B2(new_n291), .ZN(new_n645));
  OAI211_X1 g459(.A(new_n324), .B(new_n313), .C1(new_n644), .C2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(new_n328), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n323), .A2(KEYINPUT86), .A3(new_n324), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n395), .B1(new_n643), .B2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n579), .ZN(new_n651));
  INV_X1    g465(.A(G472), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n652), .B1(new_n577), .B2(new_n313), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n651), .A2(new_n653), .A3(new_n635), .ZN(new_n654));
  AND2_X1   g468(.A1(new_n650), .A2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n331), .ZN(new_n656));
  INV_X1    g470(.A(new_n378), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n385), .A2(new_n657), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n656), .B1(new_n658), .B2(new_n387), .ZN(new_n659));
  INV_X1    g473(.A(new_n526), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NOR3_X1   g475(.A1(new_n516), .A2(G478), .A3(G902), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n515), .A2(KEYINPUT33), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT33), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n664), .B1(new_n513), .B2(new_n514), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n313), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n662), .B1(new_n666), .B2(G478), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n478), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n661), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n655), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT34), .B(G104), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G6));
  NAND2_X1  g486(.A1(new_n519), .A2(new_n477), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT101), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n464), .A2(KEYINPUT100), .A3(new_n471), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n472), .ZN(new_n676));
  AOI21_X1  g490(.A(KEYINPUT100), .B1(new_n464), .B2(new_n471), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n674), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n464), .A2(new_n471), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT100), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n681), .A2(KEYINPUT101), .A3(new_n472), .A4(new_n675), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n673), .B1(new_n678), .B2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT102), .ZN(new_n684));
  INV_X1    g498(.A(new_n661), .ZN(new_n685));
  AND3_X1   g499(.A1(new_n683), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n684), .B1(new_n683), .B2(new_n685), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n655), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  XOR2_X1   g502(.A(KEYINPUT35), .B(G107), .Z(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(G9));
  NAND2_X1  g504(.A1(new_n618), .A2(new_n622), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n621), .A2(KEYINPUT36), .ZN(new_n692));
  OR2_X1    g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n691), .A2(new_n692), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n693), .A2(new_n633), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n631), .A2(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NOR3_X1   g511(.A1(new_n651), .A2(new_n653), .A3(new_n697), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n650), .A2(new_n391), .A3(new_n527), .A4(new_n698), .ZN(new_n699));
  XOR2_X1   g513(.A(KEYINPUT37), .B(G110), .Z(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(G12));
  NAND2_X1  g515(.A1(new_n659), .A2(new_n696), .ZN(new_n702));
  AND3_X1   g516(.A1(new_n577), .A2(KEYINPUT32), .A3(new_n578), .ZN(new_n703));
  AOI21_X1  g517(.A(KEYINPUT32), .B1(new_n577), .B2(new_n578), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n702), .B1(new_n705), .B2(new_n593), .ZN(new_n706));
  INV_X1    g520(.A(G900), .ZN(new_n707));
  AND2_X1   g521(.A1(new_n524), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(KEYINPUT103), .ZN(new_n709));
  INV_X1    g523(.A(new_n521), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n708), .A2(KEYINPUT103), .ZN(new_n712));
  OR2_X1    g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(new_n713), .ZN(new_n714));
  AOI211_X1 g528(.A(new_n673), .B(new_n714), .C1(new_n678), .C2(new_n682), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n706), .A2(new_n715), .A3(new_n650), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G128), .ZN(G30));
  XOR2_X1   g531(.A(new_n388), .B(KEYINPUT38), .Z(new_n718));
  NAND2_X1  g532(.A1(new_n478), .A2(new_n519), .ZN(new_n719));
  NOR4_X1   g533(.A1(new_n718), .A2(new_n656), .A3(new_n696), .A4(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n713), .B(KEYINPUT39), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n650), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(KEYINPUT40), .ZN(new_n723));
  AND2_X1   g537(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n566), .B1(new_n569), .B2(new_n556), .ZN(new_n725));
  AND2_X1   g539(.A1(new_n563), .A2(new_n725), .ZN(new_n726));
  OAI21_X1  g540(.A(G472), .B1(new_n726), .B2(G902), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n581), .A2(new_n582), .A3(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT104), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n728), .B(new_n729), .ZN(new_n730));
  OAI211_X1 g544(.A(new_n724), .B(new_n730), .C1(KEYINPUT40), .C2(new_n722), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G143), .ZN(G45));
  AOI21_X1  g546(.A(new_n697), .B1(new_n705), .B2(new_n593), .ZN(new_n733));
  AND3_X1   g547(.A1(new_n478), .A2(new_n667), .A3(new_n713), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n734), .A2(KEYINPUT105), .A3(new_n659), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT105), .ZN(new_n736));
  INV_X1    g550(.A(new_n659), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n478), .A2(new_n667), .A3(new_n713), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n736), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n733), .A2(new_n650), .A3(new_n735), .A4(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G146), .ZN(G48));
  NAND2_X1  g555(.A1(new_n321), .A2(new_n322), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n324), .B1(new_n742), .B2(new_n313), .ZN(new_n743));
  AOI211_X1 g557(.A(new_n395), .B(new_n743), .C1(new_n647), .C2(new_n648), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n744), .A2(new_n669), .A3(new_n594), .A4(new_n636), .ZN(new_n745));
  XNOR2_X1  g559(.A(KEYINPUT41), .B(G113), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n745), .B(new_n746), .ZN(G15));
  INV_X1    g561(.A(new_n637), .ZN(new_n748));
  OAI211_X1 g562(.A(new_n748), .B(new_n744), .C1(new_n686), .C2(new_n687), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G116), .ZN(G18));
  INV_X1    g564(.A(new_n702), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n744), .A2(new_n594), .A3(new_n527), .A4(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G119), .ZN(G21));
  NAND3_X1  g567(.A1(new_n631), .A2(KEYINPUT106), .A3(new_n634), .ZN(new_n754));
  INV_X1    g568(.A(new_n754), .ZN(new_n755));
  AOI21_X1  g569(.A(KEYINPUT106), .B1(new_n631), .B2(new_n634), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  AOI22_X1  g571(.A1(new_n563), .A2(KEYINPUT31), .B1(new_n575), .B2(new_n566), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n562), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(new_n578), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  NOR3_X1   g575(.A1(new_n653), .A2(new_n757), .A3(new_n761), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n737), .A2(new_n719), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n744), .A2(new_n762), .A3(new_n660), .A4(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G122), .ZN(G24));
  NAND2_X1  g579(.A1(new_n577), .A2(new_n313), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(G472), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n734), .A2(new_n767), .A3(new_n696), .A4(new_n760), .ZN(new_n768));
  INV_X1    g582(.A(new_n743), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n649), .A2(new_n396), .A3(new_n659), .A4(new_n769), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(new_n400), .ZN(G27));
  NOR2_X1   g586(.A1(new_n388), .A2(new_n656), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n396), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n641), .B1(new_n325), .B2(new_n329), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(KEYINPUT107), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT107), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n649), .A2(new_n777), .A3(new_n641), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n774), .B1(new_n776), .B2(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n779), .A2(new_n748), .A3(new_n734), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT42), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n478), .A2(KEYINPUT42), .A3(new_n667), .A4(new_n713), .ZN(new_n782));
  AOI211_X1 g596(.A(new_n774), .B(new_n782), .C1(new_n776), .C2(new_n778), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n593), .A2(new_n582), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n784), .B1(KEYINPUT108), .B2(new_n581), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT108), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n704), .A2(new_n786), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n757), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  AOI22_X1  g602(.A1(new_n780), .A2(new_n781), .B1(new_n783), .B2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(new_n235), .ZN(G33));
  NAND3_X1  g604(.A1(new_n779), .A2(new_n748), .A3(new_n715), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G134), .ZN(G36));
  AOI21_X1  g606(.A(new_n697), .B1(new_n767), .B2(new_n579), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(KEYINPUT109), .ZN(new_n794));
  AND3_X1   g608(.A1(new_n667), .A2(new_n473), .A3(new_n477), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT43), .ZN(new_n796));
  OR2_X1    g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n795), .A2(new_n796), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n794), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n793), .A2(KEYINPUT109), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  OR2_X1    g615(.A1(new_n801), .A2(KEYINPUT44), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(KEYINPUT44), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT45), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n310), .B(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(G469), .ZN(new_n806));
  NAND2_X1  g620(.A1(G469), .A2(G902), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n806), .A2(KEYINPUT46), .A3(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT46), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n809), .B(G469), .C1(new_n805), .C2(G902), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n808), .A2(new_n649), .A3(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n811), .A2(new_n396), .A3(new_n721), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n802), .A2(new_n773), .A3(new_n803), .A4(new_n813), .ZN(new_n814));
  XNOR2_X1  g628(.A(KEYINPUT110), .B(G137), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n814), .B(new_n815), .ZN(G39));
  NAND2_X1  g630(.A1(new_n811), .A2(new_n396), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT47), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n811), .A2(KEYINPUT47), .A3(new_n396), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n734), .A2(new_n635), .A3(new_n773), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n822), .A2(new_n594), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g638(.A(KEYINPUT111), .B(G140), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n824), .B(new_n825), .ZN(G42));
  AOI21_X1  g640(.A(new_n743), .B1(new_n647), .B2(new_n648), .ZN(new_n827));
  XOR2_X1   g641(.A(new_n827), .B(KEYINPUT49), .Z(new_n828));
  NOR3_X1   g642(.A1(new_n757), .A2(new_n656), .A3(new_n395), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n718), .A2(new_n829), .A3(new_n795), .ZN(new_n830));
  OR3_X1    g644(.A1(new_n730), .A2(new_n828), .A3(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n797), .A2(new_n521), .A3(new_n798), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT118), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n827), .A2(new_n396), .A3(new_n773), .ZN(new_n834));
  OR3_X1    g648(.A1(new_n832), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n833), .B1(new_n832), .B2(new_n834), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(new_n788), .ZN(new_n838));
  OAI21_X1  g652(.A(KEYINPUT48), .B1(new_n838), .B2(KEYINPUT119), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n839), .B1(KEYINPUT119), .B2(new_n838), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT48), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n838), .A2(KEYINPUT119), .A3(new_n841), .ZN(new_n842));
  NOR4_X1   g656(.A1(new_n730), .A2(new_n834), .A3(new_n635), .A4(new_n710), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n843), .A2(new_n478), .A3(new_n667), .ZN(new_n844));
  AND4_X1   g658(.A1(new_n521), .A2(new_n797), .A3(new_n762), .A4(new_n798), .ZN(new_n845));
  INV_X1    g659(.A(new_n770), .ZN(new_n846));
  AOI211_X1 g660(.A(new_n520), .B(G953), .C1(new_n845), .C2(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n842), .A2(new_n844), .A3(new_n847), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n840), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n827), .A2(new_n395), .ZN(new_n850));
  INV_X1    g664(.A(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT116), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n851), .B1(new_n821), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n853), .B1(new_n852), .B2(new_n821), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n845), .A2(new_n773), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT51), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n837), .A2(new_n767), .A3(new_n696), .A4(new_n760), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n718), .A2(new_n656), .A3(new_n744), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n845), .A2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT50), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n861), .A2(KEYINPUT117), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n860), .B(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n478), .A2(new_n667), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n843), .A2(new_n864), .ZN(new_n865));
  AND3_X1   g679(.A1(new_n858), .A2(new_n863), .A3(new_n865), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n856), .A2(new_n857), .A3(new_n866), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n855), .B1(new_n821), .B2(new_n851), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n857), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n849), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT53), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n473), .A2(new_n477), .A3(new_n519), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT113), .ZN(new_n873));
  OR2_X1    g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n668), .A2(KEYINPUT112), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT112), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n478), .A2(new_n876), .A3(new_n667), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n872), .A2(new_n873), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n874), .A2(new_n875), .A3(new_n877), .A4(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n526), .B1(new_n384), .B2(new_n390), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n879), .A2(new_n650), .A3(new_n654), .A4(new_n880), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n881), .A2(new_n699), .A3(new_n745), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n764), .A2(new_n752), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n883), .A2(new_n638), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n882), .A2(new_n884), .A3(new_n749), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n477), .A2(new_n713), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n697), .A2(new_n519), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n773), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n888), .B1(new_n678), .B2(new_n682), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n889), .A2(new_n594), .A3(new_n650), .ZN(new_n890));
  INV_X1    g704(.A(new_n768), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n779), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n791), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n789), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n885), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n891), .A2(new_n846), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n713), .B(KEYINPUT114), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n631), .A2(new_n695), .A3(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT115), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n631), .A2(KEYINPUT115), .A3(new_n695), .A4(new_n897), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n900), .A2(new_n396), .A3(new_n901), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n737), .A2(new_n902), .A3(new_n719), .ZN(new_n903));
  AND3_X1   g717(.A1(new_n649), .A2(new_n777), .A3(new_n641), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n777), .B1(new_n649), .B2(new_n641), .ZN(new_n905));
  OAI211_X1 g719(.A(new_n728), .B(new_n903), .C1(new_n904), .C2(new_n905), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n740), .A2(new_n716), .A3(new_n896), .A4(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT52), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  AND4_X1   g723(.A1(new_n594), .A2(new_n330), .A3(new_n396), .A4(new_n751), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n771), .B1(new_n910), .B2(new_n715), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n911), .A2(KEYINPUT52), .A3(new_n740), .A4(new_n906), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n909), .A2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n871), .B1(new_n895), .B2(new_n914), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n882), .A2(new_n884), .A3(new_n749), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n916), .A2(new_n789), .A3(new_n893), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n917), .A2(KEYINPUT53), .A3(new_n913), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n915), .A2(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT54), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n915), .A2(new_n918), .A3(KEYINPUT54), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n870), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NOR2_X1   g737(.A1(G952), .A2(G953), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n831), .B1(new_n923), .B2(new_n924), .ZN(G75));
  NOR2_X1   g739(.A1(new_n364), .A2(G952), .ZN(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n313), .B1(new_n915), .B2(new_n918), .ZN(new_n928));
  AOI21_X1  g742(.A(KEYINPUT56), .B1(new_n928), .B2(new_n657), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n359), .A2(new_n361), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(new_n366), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(KEYINPUT121), .ZN(new_n932));
  XOR2_X1   g746(.A(KEYINPUT120), .B(KEYINPUT55), .Z(new_n933));
  XNOR2_X1  g747(.A(new_n932), .B(new_n933), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n927), .B1(new_n929), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(KEYINPUT53), .B1(new_n917), .B2(new_n913), .ZN(new_n936));
  AND4_X1   g750(.A1(KEYINPUT53), .A2(new_n913), .A3(new_n885), .A4(new_n894), .ZN(new_n937));
  OAI21_X1  g751(.A(G902), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(KEYINPUT122), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT122), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n919), .A2(new_n940), .A3(G902), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n939), .A2(new_n380), .A3(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT56), .ZN(new_n943));
  AND2_X1   g757(.A1(new_n934), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n935), .B1(new_n942), .B2(new_n944), .ZN(G51));
  XOR2_X1   g759(.A(new_n807), .B(KEYINPUT57), .Z(new_n946));
  NAND3_X1  g760(.A1(new_n921), .A2(new_n922), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(new_n742), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n939), .A2(new_n941), .A3(G469), .A4(new_n805), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n926), .B1(new_n948), .B2(new_n949), .ZN(G54));
  AND2_X1   g764(.A1(KEYINPUT58), .A2(G475), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n939), .A2(new_n941), .A3(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(new_n468), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n939), .A2(new_n941), .A3(new_n468), .A4(new_n951), .ZN(new_n955));
  AND3_X1   g769(.A1(new_n954), .A2(new_n927), .A3(new_n955), .ZN(G60));
  NAND2_X1  g770(.A1(G478), .A2(G902), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n957), .B(KEYINPUT59), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n921), .A2(new_n922), .A3(new_n958), .ZN(new_n959));
  OR2_X1    g773(.A1(new_n663), .A2(new_n665), .ZN(new_n960));
  INV_X1    g774(.A(new_n960), .ZN(new_n961));
  AND2_X1   g775(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n959), .A2(new_n961), .ZN(new_n963));
  NOR3_X1   g777(.A1(new_n962), .A2(new_n963), .A3(new_n926), .ZN(G63));
  XNOR2_X1  g778(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n510), .A2(new_n313), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n965), .B(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n968), .B1(new_n915), .B2(new_n918), .ZN(new_n969));
  OR2_X1    g783(.A1(new_n969), .A2(new_n632), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n969), .A2(new_n694), .A3(new_n693), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n970), .A2(new_n927), .A3(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT61), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n970), .A2(new_n971), .A3(KEYINPUT61), .A4(new_n927), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n974), .A2(new_n975), .ZN(G66));
  NAND2_X1  g790(.A1(G224), .A2(G953), .ZN(new_n977));
  OAI22_X1  g791(.A1(new_n916), .A2(G953), .B1(new_n525), .B2(new_n977), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n978), .B(KEYINPUT124), .ZN(new_n979));
  INV_X1    g793(.A(G898), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n930), .B1(new_n980), .B2(G953), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n979), .B(new_n981), .ZN(G69));
  INV_X1    g796(.A(new_n722), .ZN(new_n983));
  NAND4_X1  g797(.A1(new_n983), .A2(new_n748), .A3(new_n773), .A4(new_n879), .ZN(new_n984));
  AND3_X1   g798(.A1(new_n814), .A2(new_n824), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n911), .A2(new_n740), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n986), .B(KEYINPUT125), .ZN(new_n987));
  AND3_X1   g801(.A1(new_n987), .A2(KEYINPUT62), .A3(new_n731), .ZN(new_n988));
  AOI21_X1  g802(.A(KEYINPUT62), .B1(new_n987), .B2(new_n731), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n985), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n426), .A2(new_n427), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n559), .B(new_n991), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n990), .A2(new_n364), .A3(new_n992), .ZN(new_n993));
  AND2_X1   g807(.A1(new_n992), .A2(new_n294), .ZN(new_n994));
  OAI21_X1  g808(.A(G953), .B1(new_n994), .B2(new_n707), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n788), .A2(new_n763), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n791), .B1(new_n996), .B2(new_n812), .ZN(new_n997));
  AOI211_X1 g811(.A(new_n789), .B(new_n997), .C1(new_n821), .C2(new_n823), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n998), .A2(new_n814), .A3(new_n987), .ZN(new_n999));
  MUX2_X1   g813(.A(new_n294), .B(new_n999), .S(new_n364), .Z(new_n1000));
  OAI211_X1 g814(.A(new_n993), .B(new_n995), .C1(new_n1000), .C2(new_n992), .ZN(G72));
  NAND2_X1  g815(.A1(G472), .A2(G902), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1002), .B(KEYINPUT63), .ZN(new_n1003));
  XOR2_X1   g817(.A(new_n1003), .B(KEYINPUT126), .Z(new_n1004));
  OAI21_X1  g818(.A(new_n1004), .B1(new_n990), .B2(new_n916), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n1005), .A2(new_n550), .A3(new_n586), .ZN(new_n1006));
  NAND4_X1  g820(.A1(new_n998), .A2(new_n814), .A3(new_n885), .A4(new_n987), .ZN(new_n1007));
  INV_X1    g821(.A(KEYINPUT127), .ZN(new_n1008));
  AND3_X1   g822(.A1(new_n1007), .A2(new_n1008), .A3(new_n1004), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n1008), .B1(new_n1007), .B2(new_n1004), .ZN(new_n1010));
  OAI211_X1 g824(.A(new_n566), .B(new_n560), .C1(new_n1009), .C2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n1003), .B1(new_n587), .B2(new_n563), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n926), .B1(new_n919), .B2(new_n1012), .ZN(new_n1013));
  AND3_X1   g827(.A1(new_n1006), .A2(new_n1011), .A3(new_n1013), .ZN(G57));
endmodule


