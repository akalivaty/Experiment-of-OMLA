

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581;

  XNOR2_X1 U322 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U323 ( .A(KEYINPUT82), .B(KEYINPUT0), .Z(n290) );
  OR2_X1 U324 ( .A1(n456), .A2(n572), .ZN(n457) );
  XNOR2_X1 U325 ( .A(n335), .B(n334), .ZN(n337) );
  NOR2_X1 U326 ( .A1(n576), .A2(n458), .ZN(n459) );
  XOR2_X1 U327 ( .A(n339), .B(n338), .Z(n544) );
  XNOR2_X1 U328 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n447) );
  XOR2_X1 U329 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n292) );
  XNOR2_X1 U330 ( .A(KEYINPUT90), .B(KEYINPUT91), .ZN(n291) );
  XNOR2_X1 U331 ( .A(n292), .B(n291), .ZN(n297) );
  XNOR2_X1 U332 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n293) );
  XNOR2_X1 U333 ( .A(n293), .B(KEYINPUT2), .ZN(n348) );
  XOR2_X1 U334 ( .A(n348), .B(G1GAT), .Z(n295) );
  NAND2_X1 U335 ( .A1(G225GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U336 ( .A(n295), .B(n294), .ZN(n296) );
  XNOR2_X1 U337 ( .A(n297), .B(n296), .ZN(n311) );
  XOR2_X1 U338 ( .A(G148GAT), .B(G120GAT), .Z(n299) );
  XNOR2_X1 U339 ( .A(G141GAT), .B(G127GAT), .ZN(n298) );
  XNOR2_X1 U340 ( .A(n299), .B(n298), .ZN(n303) );
  XOR2_X1 U341 ( .A(G57GAT), .B(KEYINPUT1), .Z(n301) );
  XNOR2_X1 U342 ( .A(KEYINPUT89), .B(KEYINPUT6), .ZN(n300) );
  XNOR2_X1 U343 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U344 ( .A(n303), .B(n302), .Z(n309) );
  XOR2_X1 U345 ( .A(G85GAT), .B(G162GAT), .Z(n306) );
  XNOR2_X1 U346 ( .A(G113GAT), .B(KEYINPUT81), .ZN(n304) );
  XNOR2_X1 U347 ( .A(n290), .B(n304), .ZN(n329) );
  XNOR2_X1 U348 ( .A(G29GAT), .B(n329), .ZN(n305) );
  XNOR2_X1 U349 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U350 ( .A(G134GAT), .B(n307), .ZN(n308) );
  XNOR2_X1 U351 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U352 ( .A(n311), .B(n310), .ZN(n534) );
  XOR2_X1 U353 ( .A(KEYINPUT83), .B(KEYINPUT17), .Z(n313) );
  XNOR2_X1 U354 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n312) );
  XNOR2_X1 U355 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U356 ( .A(n314), .B(G183GAT), .Z(n316) );
  XNOR2_X1 U357 ( .A(G169GAT), .B(G176GAT), .ZN(n315) );
  XNOR2_X1 U358 ( .A(n316), .B(n315), .ZN(n339) );
  XNOR2_X1 U359 ( .A(G204GAT), .B(G92GAT), .ZN(n317) );
  XNOR2_X1 U360 ( .A(n317), .B(G64GAT), .ZN(n440) );
  XOR2_X1 U361 ( .A(n440), .B(KEYINPUT93), .Z(n319) );
  NAND2_X1 U362 ( .A1(G226GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U363 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U364 ( .A(n339), .B(n320), .ZN(n328) );
  XOR2_X1 U365 ( .A(G36GAT), .B(G190GAT), .Z(n390) );
  XOR2_X1 U366 ( .A(KEYINPUT92), .B(n390), .Z(n326) );
  XNOR2_X1 U367 ( .A(G211GAT), .B(KEYINPUT87), .ZN(n321) );
  XNOR2_X1 U368 ( .A(n321), .B(KEYINPUT21), .ZN(n322) );
  XOR2_X1 U369 ( .A(n322), .B(KEYINPUT86), .Z(n324) );
  XNOR2_X1 U370 ( .A(G197GAT), .B(G218GAT), .ZN(n323) );
  XNOR2_X1 U371 ( .A(n324), .B(n323), .ZN(n352) );
  XNOR2_X1 U372 ( .A(G8GAT), .B(n352), .ZN(n325) );
  XNOR2_X1 U373 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U374 ( .A(n328), .B(n327), .Z(n536) );
  XNOR2_X1 U375 ( .A(n536), .B(KEYINPUT27), .ZN(n362) );
  NAND2_X1 U376 ( .A1(n534), .A2(n362), .ZN(n506) );
  XOR2_X1 U377 ( .A(G43GAT), .B(G134GAT), .Z(n401) );
  XOR2_X1 U378 ( .A(n401), .B(n329), .Z(n335) );
  XOR2_X1 U379 ( .A(KEYINPUT20), .B(KEYINPUT64), .Z(n331) );
  XNOR2_X1 U380 ( .A(G99GAT), .B(G190GAT), .ZN(n330) );
  XNOR2_X1 U381 ( .A(n331), .B(n330), .ZN(n333) );
  NAND2_X1 U382 ( .A1(G227GAT), .A2(G233GAT), .ZN(n332) );
  XOR2_X1 U383 ( .A(G15GAT), .B(G127GAT), .Z(n369) );
  XOR2_X1 U384 ( .A(G120GAT), .B(G71GAT), .Z(n428) );
  XOR2_X1 U385 ( .A(n369), .B(n428), .Z(n336) );
  XNOR2_X1 U386 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U387 ( .A(KEYINPUT84), .B(n544), .ZN(n355) );
  XOR2_X1 U388 ( .A(KEYINPUT23), .B(KEYINPUT22), .Z(n341) );
  XNOR2_X1 U389 ( .A(G204GAT), .B(KEYINPUT88), .ZN(n340) );
  XNOR2_X1 U390 ( .A(n341), .B(n340), .ZN(n345) );
  XOR2_X1 U391 ( .A(KEYINPUT85), .B(KEYINPUT24), .Z(n343) );
  XOR2_X1 U392 ( .A(G141GAT), .B(G22GAT), .Z(n422) );
  XOR2_X1 U393 ( .A(G50GAT), .B(G162GAT), .Z(n391) );
  XNOR2_X1 U394 ( .A(n422), .B(n391), .ZN(n342) );
  XNOR2_X1 U395 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U396 ( .A(n345), .B(n344), .Z(n347) );
  NAND2_X1 U397 ( .A1(G228GAT), .A2(G233GAT), .ZN(n346) );
  XNOR2_X1 U398 ( .A(n347), .B(n346), .ZN(n349) );
  XOR2_X1 U399 ( .A(n349), .B(n348), .Z(n354) );
  XOR2_X1 U400 ( .A(G78GAT), .B(G148GAT), .Z(n351) );
  XNOR2_X1 U401 ( .A(G106GAT), .B(KEYINPUT73), .ZN(n350) );
  XNOR2_X1 U402 ( .A(n351), .B(n350), .ZN(n441) );
  XNOR2_X1 U403 ( .A(n352), .B(n441), .ZN(n353) );
  XNOR2_X1 U404 ( .A(n354), .B(n353), .ZN(n535) );
  XNOR2_X1 U405 ( .A(n535), .B(KEYINPUT28), .ZN(n507) );
  NAND2_X1 U406 ( .A1(n355), .A2(n507), .ZN(n356) );
  NOR2_X1 U407 ( .A1(n506), .A2(n356), .ZN(n357) );
  XNOR2_X1 U408 ( .A(KEYINPUT94), .B(n357), .ZN(n368) );
  INV_X1 U409 ( .A(n544), .ZN(n487) );
  NAND2_X1 U410 ( .A1(n487), .A2(n536), .ZN(n358) );
  NAND2_X1 U411 ( .A1(n358), .A2(n535), .ZN(n359) );
  XNOR2_X1 U412 ( .A(n359), .B(KEYINPUT95), .ZN(n360) );
  XOR2_X1 U413 ( .A(KEYINPUT25), .B(n360), .Z(n364) );
  NOR2_X1 U414 ( .A1(n535), .A2(n487), .ZN(n361) );
  XNOR2_X1 U415 ( .A(KEYINPUT26), .B(n361), .ZN(n561) );
  AND2_X1 U416 ( .A1(n362), .A2(n561), .ZN(n363) );
  NOR2_X1 U417 ( .A1(n364), .A2(n363), .ZN(n365) );
  NOR2_X1 U418 ( .A1(n534), .A2(n365), .ZN(n366) );
  XNOR2_X1 U419 ( .A(KEYINPUT96), .B(n366), .ZN(n367) );
  NOR2_X1 U420 ( .A1(n368), .A2(n367), .ZN(n456) );
  XOR2_X1 U421 ( .A(G155GAT), .B(G78GAT), .Z(n371) );
  XOR2_X1 U422 ( .A(G1GAT), .B(G8GAT), .Z(n417) );
  XNOR2_X1 U423 ( .A(n417), .B(n369), .ZN(n370) );
  XNOR2_X1 U424 ( .A(n371), .B(n370), .ZN(n376) );
  XNOR2_X1 U425 ( .A(G57GAT), .B(KEYINPUT70), .ZN(n372) );
  XNOR2_X1 U426 ( .A(n372), .B(KEYINPUT13), .ZN(n429) );
  XOR2_X1 U427 ( .A(n429), .B(KEYINPUT79), .Z(n374) );
  NAND2_X1 U428 ( .A1(G231GAT), .A2(G233GAT), .ZN(n373) );
  XNOR2_X1 U429 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U430 ( .A(n376), .B(n375), .Z(n378) );
  XNOR2_X1 U431 ( .A(G22GAT), .B(G211GAT), .ZN(n377) );
  XNOR2_X1 U432 ( .A(n378), .B(n377), .ZN(n386) );
  XOR2_X1 U433 ( .A(KEYINPUT15), .B(G64GAT), .Z(n380) );
  XNOR2_X1 U434 ( .A(G183GAT), .B(G71GAT), .ZN(n379) );
  XNOR2_X1 U435 ( .A(n380), .B(n379), .ZN(n384) );
  XOR2_X1 U436 ( .A(KEYINPUT78), .B(KEYINPUT12), .Z(n382) );
  XNOR2_X1 U437 ( .A(KEYINPUT80), .B(KEYINPUT14), .ZN(n381) );
  XNOR2_X1 U438 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U439 ( .A(n384), .B(n383), .Z(n385) );
  XNOR2_X1 U440 ( .A(n386), .B(n385), .ZN(n572) );
  INV_X1 U441 ( .A(n572), .ZN(n527) );
  XOR2_X1 U442 ( .A(G29GAT), .B(KEYINPUT7), .Z(n388) );
  XNOR2_X1 U443 ( .A(KEYINPUT68), .B(KEYINPUT8), .ZN(n387) );
  XNOR2_X1 U444 ( .A(n388), .B(n387), .ZN(n419) );
  XNOR2_X1 U445 ( .A(G99GAT), .B(G85GAT), .ZN(n389) );
  XNOR2_X1 U446 ( .A(n389), .B(KEYINPUT74), .ZN(n433) );
  XNOR2_X1 U447 ( .A(n419), .B(n433), .ZN(n405) );
  XOR2_X1 U448 ( .A(n391), .B(n390), .Z(n393) );
  NAND2_X1 U449 ( .A1(G232GAT), .A2(G233GAT), .ZN(n392) );
  XNOR2_X1 U450 ( .A(n393), .B(n392), .ZN(n397) );
  XOR2_X1 U451 ( .A(G92GAT), .B(KEYINPUT76), .Z(n395) );
  XNOR2_X1 U452 ( .A(G106GAT), .B(KEYINPUT9), .ZN(n394) );
  XNOR2_X1 U453 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U454 ( .A(n397), .B(n396), .Z(n403) );
  XOR2_X1 U455 ( .A(KEYINPUT10), .B(KEYINPUT77), .Z(n399) );
  XNOR2_X1 U456 ( .A(G218GAT), .B(KEYINPUT11), .ZN(n398) );
  XNOR2_X1 U457 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U458 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U459 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U460 ( .A(n405), .B(n404), .ZN(n531) );
  INV_X1 U461 ( .A(n531), .ZN(n555) );
  NOR2_X1 U462 ( .A1(n527), .A2(n555), .ZN(n406) );
  XOR2_X1 U463 ( .A(KEYINPUT16), .B(n406), .Z(n407) );
  NOR2_X1 U464 ( .A1(n456), .A2(n407), .ZN(n408) );
  XNOR2_X1 U465 ( .A(KEYINPUT97), .B(n408), .ZN(n473) );
  XOR2_X1 U466 ( .A(KEYINPUT66), .B(G15GAT), .Z(n410) );
  XNOR2_X1 U467 ( .A(G169GAT), .B(G113GAT), .ZN(n409) );
  XNOR2_X1 U468 ( .A(n410), .B(n409), .ZN(n414) );
  XOR2_X1 U469 ( .A(KEYINPUT69), .B(KEYINPUT65), .Z(n412) );
  XNOR2_X1 U470 ( .A(KEYINPUT30), .B(KEYINPUT29), .ZN(n411) );
  XNOR2_X1 U471 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U472 ( .A(n414), .B(n413), .ZN(n427) );
  XOR2_X1 U473 ( .A(G197GAT), .B(G43GAT), .Z(n416) );
  XNOR2_X1 U474 ( .A(G50GAT), .B(G36GAT), .ZN(n415) );
  XNOR2_X1 U475 ( .A(n416), .B(n415), .ZN(n418) );
  XOR2_X1 U476 ( .A(n418), .B(n417), .Z(n425) );
  XOR2_X1 U477 ( .A(n419), .B(KEYINPUT67), .Z(n421) );
  NAND2_X1 U478 ( .A1(G229GAT), .A2(G233GAT), .ZN(n420) );
  XNOR2_X1 U479 ( .A(n421), .B(n420), .ZN(n423) );
  XNOR2_X1 U480 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U481 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U482 ( .A(n427), .B(n426), .ZN(n545) );
  INV_X1 U483 ( .A(n545), .ZN(n563) );
  XNOR2_X1 U484 ( .A(n429), .B(n428), .ZN(n431) );
  AND2_X1 U485 ( .A1(G230GAT), .A2(G233GAT), .ZN(n430) );
  XNOR2_X1 U486 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U487 ( .A(n432), .B(KEYINPUT71), .Z(n435) );
  XNOR2_X1 U488 ( .A(n433), .B(KEYINPUT33), .ZN(n434) );
  XOR2_X1 U489 ( .A(n435), .B(n434), .Z(n439) );
  XOR2_X1 U490 ( .A(KEYINPUT72), .B(KEYINPUT32), .Z(n437) );
  XNOR2_X1 U491 ( .A(G176GAT), .B(KEYINPUT31), .ZN(n436) );
  XNOR2_X1 U492 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U493 ( .A(n439), .B(n438), .ZN(n443) );
  XNOR2_X1 U494 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U495 ( .A(n443), .B(n442), .ZN(n567) );
  NOR2_X1 U496 ( .A1(n563), .A2(n567), .ZN(n444) );
  XNOR2_X1 U497 ( .A(n444), .B(KEYINPUT75), .ZN(n460) );
  NOR2_X1 U498 ( .A1(n473), .A2(n460), .ZN(n445) );
  XNOR2_X1 U499 ( .A(n445), .B(KEYINPUT98), .ZN(n453) );
  NAND2_X1 U500 ( .A1(n534), .A2(n453), .ZN(n446) );
  XNOR2_X1 U501 ( .A(n447), .B(n446), .ZN(G1324GAT) );
  XOR2_X1 U502 ( .A(G8GAT), .B(KEYINPUT99), .Z(n449) );
  NAND2_X1 U503 ( .A1(n453), .A2(n536), .ZN(n448) );
  XNOR2_X1 U504 ( .A(n449), .B(n448), .ZN(G1325GAT) );
  XOR2_X1 U505 ( .A(KEYINPUT35), .B(KEYINPUT100), .Z(n451) );
  NAND2_X1 U506 ( .A1(n453), .A2(n487), .ZN(n450) );
  XNOR2_X1 U507 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U508 ( .A(G15GAT), .B(n452), .ZN(G1326GAT) );
  XOR2_X1 U509 ( .A(G22GAT), .B(KEYINPUT101), .Z(n455) );
  INV_X1 U510 ( .A(n507), .ZN(n491) );
  NAND2_X1 U511 ( .A1(n491), .A2(n453), .ZN(n454) );
  XNOR2_X1 U512 ( .A(n455), .B(n454), .ZN(G1327GAT) );
  XNOR2_X1 U513 ( .A(n531), .B(KEYINPUT36), .ZN(n576) );
  XNOR2_X1 U514 ( .A(KEYINPUT102), .B(n457), .ZN(n458) );
  XNOR2_X1 U515 ( .A(KEYINPUT37), .B(n459), .ZN(n484) );
  NOR2_X1 U516 ( .A1(n484), .A2(n460), .ZN(n463) );
  XOR2_X1 U517 ( .A(KEYINPUT104), .B(KEYINPUT38), .Z(n461) );
  XNOR2_X1 U518 ( .A(KEYINPUT103), .B(n461), .ZN(n462) );
  XNOR2_X2 U519 ( .A(n463), .B(n462), .ZN(n471) );
  NAND2_X1 U520 ( .A1(n534), .A2(n471), .ZN(n465) );
  XOR2_X1 U521 ( .A(G29GAT), .B(KEYINPUT39), .Z(n464) );
  XNOR2_X1 U522 ( .A(n465), .B(n464), .ZN(G1328GAT) );
  NAND2_X1 U523 ( .A1(n536), .A2(n471), .ZN(n466) );
  XNOR2_X1 U524 ( .A(n466), .B(G36GAT), .ZN(G1329GAT) );
  XNOR2_X1 U525 ( .A(G43GAT), .B(KEYINPUT106), .ZN(n470) );
  XOR2_X1 U526 ( .A(KEYINPUT105), .B(KEYINPUT40), .Z(n468) );
  NAND2_X1 U527 ( .A1(n471), .A2(n487), .ZN(n467) );
  XNOR2_X1 U528 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U529 ( .A(n470), .B(n469), .ZN(G1330GAT) );
  NAND2_X1 U530 ( .A1(n491), .A2(n471), .ZN(n472) );
  XNOR2_X1 U531 ( .A(G50GAT), .B(n472), .ZN(G1331GAT) );
  XNOR2_X1 U532 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n476) );
  XNOR2_X1 U533 ( .A(KEYINPUT41), .B(n567), .ZN(n521) );
  INV_X1 U534 ( .A(n521), .ZN(n551) );
  NAND2_X1 U535 ( .A1(n551), .A2(n563), .ZN(n483) );
  NOR2_X1 U536 ( .A1(n483), .A2(n473), .ZN(n474) );
  XOR2_X1 U537 ( .A(KEYINPUT107), .B(n474), .Z(n479) );
  NAND2_X1 U538 ( .A1(n534), .A2(n479), .ZN(n475) );
  XNOR2_X1 U539 ( .A(n476), .B(n475), .ZN(G1332GAT) );
  NAND2_X1 U540 ( .A1(n536), .A2(n479), .ZN(n477) );
  XNOR2_X1 U541 ( .A(n477), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U542 ( .A1(n487), .A2(n479), .ZN(n478) );
  XNOR2_X1 U543 ( .A(n478), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U544 ( .A(KEYINPUT108), .B(KEYINPUT43), .Z(n481) );
  NAND2_X1 U545 ( .A1(n479), .A2(n491), .ZN(n480) );
  XNOR2_X1 U546 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U547 ( .A(G78GAT), .B(n482), .ZN(G1335GAT) );
  NOR2_X1 U548 ( .A1(n484), .A2(n483), .ZN(n492) );
  NAND2_X1 U549 ( .A1(n534), .A2(n492), .ZN(n485) );
  XNOR2_X1 U550 ( .A(G85GAT), .B(n485), .ZN(G1336GAT) );
  NAND2_X1 U551 ( .A1(n536), .A2(n492), .ZN(n486) );
  XNOR2_X1 U552 ( .A(n486), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U553 ( .A(KEYINPUT109), .B(KEYINPUT110), .Z(n489) );
  NAND2_X1 U554 ( .A1(n492), .A2(n487), .ZN(n488) );
  XNOR2_X1 U555 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U556 ( .A(G99GAT), .B(n490), .ZN(G1338GAT) );
  NAND2_X1 U557 ( .A1(n492), .A2(n491), .ZN(n493) );
  XNOR2_X1 U558 ( .A(n493), .B(KEYINPUT44), .ZN(n494) );
  XNOR2_X1 U559 ( .A(G106GAT), .B(n494), .ZN(G1339GAT) );
  XOR2_X1 U560 ( .A(KEYINPUT47), .B(KEYINPUT111), .Z(n499) );
  NOR2_X1 U561 ( .A1(n563), .A2(n521), .ZN(n495) );
  XNOR2_X1 U562 ( .A(n495), .B(KEYINPUT46), .ZN(n496) );
  NOR2_X1 U563 ( .A1(n572), .A2(n496), .ZN(n497) );
  NAND2_X1 U564 ( .A1(n497), .A2(n531), .ZN(n498) );
  XNOR2_X1 U565 ( .A(n499), .B(n498), .ZN(n504) );
  NOR2_X1 U566 ( .A1(n527), .A2(n576), .ZN(n500) );
  XNOR2_X1 U567 ( .A(n500), .B(KEYINPUT45), .ZN(n501) );
  NAND2_X1 U568 ( .A1(n501), .A2(n563), .ZN(n502) );
  NOR2_X1 U569 ( .A1(n567), .A2(n502), .ZN(n503) );
  NOR2_X1 U570 ( .A1(n504), .A2(n503), .ZN(n505) );
  XNOR2_X1 U571 ( .A(KEYINPUT48), .B(n505), .ZN(n538) );
  NOR2_X1 U572 ( .A1(n538), .A2(n506), .ZN(n519) );
  NAND2_X1 U573 ( .A1(n519), .A2(n507), .ZN(n508) );
  NOR2_X1 U574 ( .A1(n544), .A2(n508), .ZN(n515) );
  NAND2_X1 U575 ( .A1(n545), .A2(n515), .ZN(n509) );
  XNOR2_X1 U576 ( .A(G113GAT), .B(n509), .ZN(G1340GAT) );
  XOR2_X1 U577 ( .A(G120GAT), .B(KEYINPUT49), .Z(n511) );
  NAND2_X1 U578 ( .A1(n515), .A2(n551), .ZN(n510) );
  XNOR2_X1 U579 ( .A(n511), .B(n510), .ZN(G1341GAT) );
  XOR2_X1 U580 ( .A(KEYINPUT50), .B(KEYINPUT112), .Z(n513) );
  NAND2_X1 U581 ( .A1(n515), .A2(n572), .ZN(n512) );
  XNOR2_X1 U582 ( .A(n513), .B(n512), .ZN(n514) );
  XOR2_X1 U583 ( .A(G127GAT), .B(n514), .Z(G1342GAT) );
  XOR2_X1 U584 ( .A(KEYINPUT51), .B(KEYINPUT113), .Z(n517) );
  NAND2_X1 U585 ( .A1(n515), .A2(n555), .ZN(n516) );
  XNOR2_X1 U586 ( .A(n517), .B(n516), .ZN(n518) );
  XOR2_X1 U587 ( .A(G134GAT), .B(n518), .Z(G1343GAT) );
  NAND2_X1 U588 ( .A1(n519), .A2(n561), .ZN(n530) );
  NOR2_X1 U589 ( .A1(n563), .A2(n530), .ZN(n520) );
  XOR2_X1 U590 ( .A(G141GAT), .B(n520), .Z(G1344GAT) );
  NOR2_X1 U591 ( .A1(n521), .A2(n530), .ZN(n526) );
  XOR2_X1 U592 ( .A(KEYINPUT53), .B(KEYINPUT115), .Z(n523) );
  XNOR2_X1 U593 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n522) );
  XNOR2_X1 U594 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U595 ( .A(KEYINPUT114), .B(n524), .ZN(n525) );
  XNOR2_X1 U596 ( .A(n526), .B(n525), .ZN(G1345GAT) );
  NOR2_X1 U597 ( .A1(n527), .A2(n530), .ZN(n528) );
  XOR2_X1 U598 ( .A(KEYINPUT116), .B(n528), .Z(n529) );
  XNOR2_X1 U599 ( .A(G155GAT), .B(n529), .ZN(G1346GAT) );
  NOR2_X1 U600 ( .A1(n531), .A2(n530), .ZN(n533) );
  XNOR2_X1 U601 ( .A(G162GAT), .B(KEYINPUT117), .ZN(n532) );
  XNOR2_X1 U602 ( .A(n533), .B(n532), .ZN(G1347GAT) );
  INV_X1 U603 ( .A(n534), .ZN(n560) );
  AND2_X1 U604 ( .A1(n560), .A2(n535), .ZN(n540) );
  XOR2_X1 U605 ( .A(n536), .B(KEYINPUT118), .Z(n537) );
  NOR2_X1 U606 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U607 ( .A(KEYINPUT54), .B(n539), .ZN(n559) );
  NAND2_X1 U608 ( .A1(n540), .A2(n559), .ZN(n541) );
  XNOR2_X1 U609 ( .A(n541), .B(KEYINPUT55), .ZN(n542) );
  XNOR2_X1 U610 ( .A(n542), .B(KEYINPUT119), .ZN(n543) );
  NOR2_X1 U611 ( .A1(n544), .A2(n543), .ZN(n556) );
  NAND2_X1 U612 ( .A1(n556), .A2(n545), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n546), .B(KEYINPUT120), .ZN(n547) );
  XNOR2_X1 U614 ( .A(G169GAT), .B(n547), .ZN(G1348GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n549) );
  XNOR2_X1 U616 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n548) );
  XNOR2_X1 U617 ( .A(n549), .B(n548), .ZN(n550) );
  XOR2_X1 U618 ( .A(KEYINPUT56), .B(n550), .Z(n553) );
  NAND2_X1 U619 ( .A1(n556), .A2(n551), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(G1349GAT) );
  NAND2_X1 U621 ( .A1(n572), .A2(n556), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n554), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U623 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n558) );
  NAND2_X1 U624 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n558), .B(n557), .ZN(G1351GAT) );
  AND2_X1 U626 ( .A1(n560), .A2(n559), .ZN(n562) );
  NAND2_X1 U627 ( .A1(n562), .A2(n561), .ZN(n575) );
  NOR2_X1 U628 ( .A1(n563), .A2(n575), .ZN(n565) );
  XNOR2_X1 U629 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U631 ( .A(G197GAT), .B(n566), .ZN(G1352GAT) );
  XOR2_X1 U632 ( .A(KEYINPUT61), .B(KEYINPUT123), .Z(n569) );
  INV_X1 U633 ( .A(n575), .ZN(n571) );
  NAND2_X1 U634 ( .A1(n571), .A2(n567), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(n570) );
  XOR2_X1 U636 ( .A(G204GAT), .B(n570), .Z(G1353GAT) );
  NAND2_X1 U637 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U638 ( .A(n573), .B(KEYINPUT124), .ZN(n574) );
  XNOR2_X1 U639 ( .A(G211GAT), .B(n574), .ZN(G1354GAT) );
  NOR2_X1 U640 ( .A1(n576), .A2(n575), .ZN(n581) );
  XOR2_X1 U641 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n578) );
  XNOR2_X1 U642 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U644 ( .A(KEYINPUT125), .B(n579), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n581), .B(n580), .ZN(G1355GAT) );
endmodule

