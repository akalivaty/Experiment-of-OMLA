//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 1 0 1 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 1 1 0 1 1 1 0 1 1 0 0 0 1 0 0 1 1 0 0 1 1 0 1 0 0 0 1 1 1 0 1 0 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:51 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n756, new_n757, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n917, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G143), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G128), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT1), .ZN(new_n193));
  AOI21_X1  g007(.A(new_n193), .B1(G143), .B2(new_n187), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n191), .B1(new_n192), .B2(new_n194), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n188), .A2(new_n190), .A3(new_n193), .A4(G128), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT11), .ZN(new_n198));
  INV_X1    g012(.A(G134), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n198), .B1(new_n199), .B2(G137), .ZN(new_n200));
  INV_X1    g014(.A(G137), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n201), .A2(KEYINPUT11), .A3(G134), .ZN(new_n202));
  INV_X1    g016(.A(G131), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n199), .A2(G137), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n200), .A2(new_n202), .A3(new_n203), .A4(new_n204), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n199), .A2(G137), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n201), .A2(G134), .ZN(new_n207));
  OAI21_X1  g021(.A(G131), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  AND3_X1   g022(.A1(new_n205), .A2(new_n208), .A3(KEYINPUT68), .ZN(new_n209));
  AOI21_X1  g023(.A(KEYINPUT68), .B1(new_n205), .B2(new_n208), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n197), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n189), .A2(G146), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n187), .A2(G143), .ZN(new_n213));
  NAND2_X1  g027(.A1(KEYINPUT0), .A2(G128), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  NOR2_X1   g029(.A1(KEYINPUT0), .A2(G128), .ZN(new_n216));
  OAI22_X1  g030(.A1(new_n212), .A2(new_n213), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n188), .A2(new_n190), .A3(new_n214), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n200), .A2(new_n202), .A3(new_n204), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G131), .ZN(new_n220));
  AOI221_X4 g034(.A(KEYINPUT67), .B1(new_n217), .B2(new_n218), .C1(new_n220), .C2(new_n205), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT67), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n220), .A2(new_n205), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n217), .A2(new_n218), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n222), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n211), .B1(new_n221), .B2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT66), .ZN(new_n227));
  INV_X1    g041(.A(G119), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n227), .B1(new_n228), .B2(G116), .ZN(new_n229));
  INV_X1    g043(.A(G116), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n230), .A2(KEYINPUT66), .A3(G119), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n230), .A2(G119), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(KEYINPUT2), .A2(G113), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(KEYINPUT65), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT65), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n238), .A2(KEYINPUT2), .A3(G113), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  NOR2_X1   g054(.A1(KEYINPUT2), .A2(G113), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n235), .A2(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n233), .B1(new_n229), .B2(new_n231), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n241), .B1(new_n237), .B2(new_n239), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  AND3_X1   g061(.A1(new_n244), .A2(KEYINPUT69), .A3(new_n247), .ZN(new_n248));
  AOI21_X1  g062(.A(KEYINPUT69), .B1(new_n244), .B2(new_n247), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n226), .A2(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(KEYINPUT11), .B1(new_n201), .B2(G134), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n252), .A2(new_n207), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n203), .B1(new_n253), .B2(new_n202), .ZN(new_n254));
  INV_X1    g068(.A(new_n205), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n224), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  AND2_X1   g070(.A1(new_n205), .A2(new_n208), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(new_n197), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT30), .ZN(new_n259));
  AND3_X1   g073(.A1(new_n256), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n256), .A2(KEYINPUT67), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n223), .A2(new_n222), .A3(new_n224), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n205), .A2(new_n208), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT68), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n205), .A2(new_n208), .A3(KEYINPUT68), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  AOI22_X1  g082(.A1(new_n262), .A2(new_n263), .B1(new_n197), .B2(new_n268), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n261), .B1(new_n269), .B2(new_n259), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n244), .A2(new_n247), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n251), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT72), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT31), .ZN(new_n274));
  INV_X1    g088(.A(G237), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(KEYINPUT70), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT70), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(G237), .ZN(new_n278));
  OR2_X1    g092(.A1(KEYINPUT71), .A2(G953), .ZN(new_n279));
  NAND2_X1  g093(.A1(KEYINPUT71), .A2(G953), .ZN(new_n280));
  AOI22_X1  g094(.A1(new_n276), .A2(new_n278), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(G210), .ZN(new_n282));
  XNOR2_X1  g096(.A(new_n282), .B(G101), .ZN(new_n283));
  XNOR2_X1  g097(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n284));
  XNOR2_X1  g098(.A(new_n283), .B(new_n284), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n272), .A2(new_n273), .A3(new_n274), .A4(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n250), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n269), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n260), .B1(new_n226), .B2(KEYINPUT30), .ZN(new_n289));
  INV_X1    g103(.A(new_n271), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n288), .B(new_n285), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(KEYINPUT72), .B1(new_n291), .B2(KEYINPUT31), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n286), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n290), .B1(new_n256), .B2(new_n258), .ZN(new_n294));
  OAI21_X1  g108(.A(KEYINPUT28), .B1(new_n251), .B2(new_n294), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n211), .B(new_n256), .C1(new_n248), .C2(new_n249), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT73), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT28), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n297), .B1(new_n296), .B2(new_n298), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n295), .A2(new_n299), .A3(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n285), .ZN(new_n303));
  AOI22_X1  g117(.A1(new_n302), .A2(new_n303), .B1(new_n291), .B2(KEYINPUT31), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n293), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(KEYINPUT74), .ZN(new_n306));
  NOR2_X1   g120(.A1(G472), .A2(G902), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT74), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n293), .A2(new_n308), .A3(new_n304), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n306), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT32), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(KEYINPUT75), .B1(new_n301), .B2(new_n299), .ZN(new_n313));
  INV_X1    g127(.A(new_n299), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT75), .ZN(new_n315));
  NOR3_X1   g129(.A1(new_n314), .A2(new_n315), .A3(new_n300), .ZN(new_n316));
  OR2_X1    g130(.A1(new_n313), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n226), .A2(new_n250), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n288), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(KEYINPUT28), .ZN(new_n320));
  NAND4_X1  g134(.A1(new_n317), .A2(KEYINPUT29), .A3(new_n285), .A4(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(G902), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n272), .A2(new_n303), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n324), .B1(new_n285), .B2(new_n302), .ZN(new_n325));
  OAI211_X1 g139(.A(new_n321), .B(new_n322), .C1(new_n325), .C2(KEYINPUT29), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(G472), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n306), .A2(KEYINPUT32), .A3(new_n307), .A4(new_n309), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n312), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  XOR2_X1   g143(.A(KEYINPUT9), .B(G234), .Z(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(G221), .B1(new_n331), .B2(G902), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n279), .A2(new_n280), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(G227), .ZN(new_n334));
  XNOR2_X1  g148(.A(G110), .B(G140), .ZN(new_n335));
  XNOR2_X1  g149(.A(new_n334), .B(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(new_n223), .ZN(new_n338));
  OAI21_X1  g152(.A(KEYINPUT80), .B1(new_n212), .B2(new_n193), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT80), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n188), .A2(new_n340), .A3(KEYINPUT1), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n339), .A2(G128), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(new_n191), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(new_n196), .ZN(new_n344));
  INV_X1    g158(.A(G107), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT3), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n345), .B1(new_n346), .B2(G104), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(G104), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(G101), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(KEYINPUT79), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT79), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(G101), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  XNOR2_X1  g168(.A(KEYINPUT78), .B(G107), .ZN(new_n355));
  OAI211_X1 g169(.A(new_n349), .B(new_n354), .C1(new_n348), .C2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(G104), .A2(G107), .ZN(new_n357));
  OAI211_X1 g171(.A(G101), .B(new_n357), .C1(new_n355), .C2(G104), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n344), .A2(new_n360), .A3(KEYINPUT81), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT81), .ZN(new_n362));
  INV_X1    g176(.A(new_n196), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n363), .B1(new_n342), .B2(new_n191), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n362), .B1(new_n364), .B2(new_n359), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n361), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT10), .ZN(new_n367));
  AOI21_X1  g181(.A(KEYINPUT82), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT82), .ZN(new_n369));
  AOI211_X1 g183(.A(new_n369), .B(KEYINPUT10), .C1(new_n361), .C2(new_n365), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n345), .A2(KEYINPUT78), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT78), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(G107), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n348), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(G104), .ZN(new_n376));
  AOI21_X1  g190(.A(G107), .B1(new_n376), .B2(KEYINPUT3), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n376), .A2(KEYINPUT3), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g193(.A(G101), .B1(new_n375), .B2(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n380), .A2(KEYINPUT4), .A3(new_n356), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT4), .ZN(new_n382));
  OAI211_X1 g196(.A(new_n382), .B(G101), .C1(new_n375), .C2(new_n379), .ZN(new_n383));
  AND3_X1   g197(.A1(new_n381), .A2(new_n224), .A3(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT83), .ZN(new_n385));
  AND3_X1   g199(.A1(new_n356), .A2(new_n385), .A3(new_n358), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n385), .B1(new_n356), .B2(new_n358), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n197), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n384), .B1(new_n390), .B2(KEYINPUT10), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n338), .B1(new_n371), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n366), .A2(new_n367), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n369), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n366), .A2(KEYINPUT82), .A3(new_n367), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n394), .A2(new_n391), .A3(new_n338), .A4(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n337), .B1(new_n392), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n389), .A2(new_n359), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n366), .A2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT84), .ZN(new_n401));
  AOI21_X1  g215(.A(KEYINPUT12), .B1(new_n223), .B2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n400), .A2(new_n223), .A3(new_n403), .ZN(new_n404));
  AOI22_X1  g218(.A1(new_n361), .A2(new_n365), .B1(new_n389), .B2(new_n359), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n402), .B1(new_n405), .B2(new_n338), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(KEYINPUT85), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT85), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n404), .A2(new_n406), .A3(new_n409), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n408), .A2(new_n396), .A3(new_n336), .A4(new_n410), .ZN(new_n411));
  AOI211_X1 g225(.A(G469), .B(G902), .C1(new_n398), .C2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(G469), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n394), .A2(new_n391), .A3(new_n395), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(new_n223), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n415), .A2(new_n396), .A3(new_n336), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n396), .A2(new_n407), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(new_n337), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n413), .B1(new_n419), .B2(new_n322), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n332), .B1(new_n412), .B2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(G475), .ZN(new_n422));
  INV_X1    g236(.A(G125), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n423), .A2(G140), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT16), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT76), .ZN(new_n428));
  INV_X1    g242(.A(G140), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n428), .B1(new_n429), .B2(G125), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n423), .A2(KEYINPUT76), .A3(G140), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n424), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n427), .B1(new_n432), .B2(new_n426), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n433), .B(G146), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n281), .A2(G214), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(new_n189), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n281), .A2(G143), .A3(G214), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n439), .A2(KEYINPUT17), .A3(G131), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(G131), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n437), .A2(new_n438), .A3(new_n203), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  OAI211_X1 g257(.A(new_n435), .B(new_n440), .C1(new_n443), .C2(KEYINPUT17), .ZN(new_n444));
  XNOR2_X1  g258(.A(G113), .B(G122), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n445), .B(new_n376), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n423), .A2(G140), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n425), .A2(new_n447), .A3(new_n187), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n448), .B1(new_n432), .B2(new_n187), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT18), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n450), .A2(new_n203), .ZN(new_n451));
  OAI221_X1 g265(.A(new_n449), .B1(new_n439), .B2(new_n451), .C1(new_n441), .C2(new_n450), .ZN(new_n452));
  AND3_X1   g266(.A1(new_n444), .A2(new_n446), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n433), .A2(G146), .ZN(new_n454));
  XOR2_X1   g268(.A(KEYINPUT94), .B(KEYINPUT19), .Z(new_n455));
  NAND3_X1  g269(.A1(new_n455), .A2(new_n425), .A3(new_n447), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT19), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n456), .B(new_n187), .C1(new_n457), .C2(new_n432), .ZN(new_n458));
  OR2_X1    g272(.A1(new_n458), .A2(KEYINPUT95), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(KEYINPUT95), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n443), .A2(new_n454), .A3(new_n459), .A4(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n446), .B1(new_n461), .B2(new_n452), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n422), .B(new_n322), .C1(new_n453), .C2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(KEYINPUT20), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n444), .A2(new_n446), .A3(new_n452), .ZN(new_n465));
  AND2_X1   g279(.A1(new_n461), .A2(new_n452), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n465), .B1(new_n466), .B2(new_n446), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT20), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n467), .A2(new_n468), .A3(new_n422), .A4(new_n322), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n446), .B1(new_n444), .B2(new_n452), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n322), .B1(new_n453), .B2(new_n470), .ZN(new_n471));
  XNOR2_X1  g285(.A(KEYINPUT96), .B(G475), .ZN(new_n472));
  AOI22_X1  g286(.A1(new_n464), .A2(new_n469), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(G953), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(G952), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n475), .B1(G234), .B2(G237), .ZN(new_n476));
  AOI211_X1 g290(.A(new_n322), .B(new_n333), .C1(G234), .C2(G237), .ZN(new_n477));
  XOR2_X1   g291(.A(KEYINPUT21), .B(G898), .Z(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n476), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  AND2_X1   g295(.A1(KEYINPUT64), .A2(G128), .ZN(new_n482));
  NOR2_X1   g296(.A1(KEYINPUT64), .A2(G128), .ZN(new_n483));
  OAI21_X1  g297(.A(G143), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n189), .A2(G128), .ZN(new_n485));
  AND3_X1   g299(.A1(new_n484), .A2(new_n199), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n199), .B1(new_n484), .B2(new_n485), .ZN(new_n487));
  OAI21_X1  g301(.A(KEYINPUT99), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n484), .A2(new_n485), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(G134), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n484), .A2(new_n199), .A3(new_n485), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT99), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  AND3_X1   g307(.A1(new_n230), .A2(KEYINPUT14), .A3(G122), .ZN(new_n494));
  XNOR2_X1  g308(.A(G116), .B(G122), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT14), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n372), .A2(new_n374), .ZN(new_n498));
  AOI22_X1  g312(.A1(new_n497), .A2(G107), .B1(new_n498), .B2(new_n495), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n488), .A2(new_n493), .A3(new_n499), .ZN(new_n500));
  XOR2_X1   g314(.A(G116), .B(G122), .Z(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(new_n355), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n498), .A2(new_n495), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT97), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  XNOR2_X1  g320(.A(KEYINPUT98), .B(KEYINPUT13), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n507), .A2(G128), .A3(new_n189), .ZN(new_n508));
  OAI211_X1 g322(.A(G134), .B(new_n508), .C1(new_n489), .C2(new_n507), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n502), .A2(KEYINPUT97), .A3(new_n503), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n506), .A2(new_n509), .A3(new_n491), .A4(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n500), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(KEYINPUT100), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT100), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n500), .A2(new_n511), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(G217), .ZN(new_n517));
  NOR3_X1   g331(.A1(new_n331), .A2(new_n517), .A3(G953), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n513), .A2(new_n518), .A3(new_n515), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n520), .A2(new_n521), .A3(new_n322), .ZN(new_n522));
  INV_X1    g336(.A(G478), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n523), .A2(KEYINPUT15), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n522), .B(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n473), .A2(new_n481), .A3(new_n526), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n421), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n517), .B1(G234), .B2(new_n322), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n333), .A2(G221), .A3(G234), .ZN(new_n531));
  XNOR2_X1  g345(.A(KEYINPUT22), .B(G137), .ZN(new_n532));
  XNOR2_X1  g346(.A(new_n531), .B(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT23), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n534), .B1(new_n228), .B2(G128), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n228), .A2(G128), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n192), .A2(G119), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n535), .B(new_n536), .C1(new_n537), .C2(new_n534), .ZN(new_n538));
  AND2_X1   g352(.A1(new_n537), .A2(new_n536), .ZN(new_n539));
  XOR2_X1   g353(.A(KEYINPUT24), .B(G110), .Z(new_n540));
  AOI22_X1  g354(.A1(G110), .A2(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n434), .A2(new_n541), .ZN(new_n542));
  OAI22_X1  g356(.A1(new_n538), .A2(G110), .B1(new_n539), .B2(new_n540), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n543), .A2(new_n454), .A3(new_n448), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT77), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(KEYINPUT77), .B1(new_n542), .B2(new_n544), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n533), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n533), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n550), .B1(new_n545), .B2(new_n546), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n549), .A2(new_n322), .A3(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT25), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n549), .A2(KEYINPUT25), .A3(new_n322), .A4(new_n551), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n530), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  AND2_X1   g370(.A1(new_n549), .A2(new_n551), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n529), .A2(G902), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(G214), .B1(G237), .B2(G902), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(G210), .B1(G237), .B2(G902), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  XNOR2_X1  g377(.A(KEYINPUT90), .B(G224), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n565), .A2(G953), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n217), .A2(G125), .A3(new_n218), .ZN(new_n567));
  OAI211_X1 g381(.A(KEYINPUT89), .B(new_n567), .C1(new_n197), .C2(G125), .ZN(new_n568));
  OR2_X1    g382(.A1(new_n567), .A2(KEYINPUT89), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n566), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n568), .A2(new_n569), .A3(new_n566), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  AND3_X1   g388(.A1(new_n380), .A2(KEYINPUT4), .A3(new_n356), .ZN(new_n575));
  AND2_X1   g389(.A1(new_n245), .A2(new_n246), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n245), .A2(new_n246), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n383), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  OAI21_X1  g392(.A(KEYINPUT86), .B1(new_n575), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n245), .A2(KEYINPUT5), .ZN(new_n580));
  INV_X1    g394(.A(G113), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT5), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n581), .B1(new_n233), .B2(new_n582), .ZN(new_n583));
  AOI22_X1  g397(.A1(new_n580), .A2(new_n583), .B1(new_n246), .B2(new_n245), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n584), .B1(new_n386), .B2(new_n387), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT86), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n381), .A2(new_n271), .A3(new_n586), .A4(new_n383), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n579), .A2(new_n585), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(KEYINPUT87), .ZN(new_n589));
  XOR2_X1   g403(.A(G110), .B(G122), .Z(new_n590));
  INV_X1    g404(.A(KEYINPUT87), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n579), .A2(new_n591), .A3(new_n585), .A4(new_n587), .ZN(new_n592));
  AND3_X1   g406(.A1(new_n589), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n590), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n579), .A2(new_n594), .A3(new_n585), .A4(new_n587), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT88), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n595), .B(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(KEYINPUT6), .B1(new_n593), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n589), .A2(new_n590), .A3(new_n592), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT6), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n574), .B1(new_n598), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n568), .A2(new_n569), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n603), .A2(KEYINPUT7), .ZN(new_n604));
  AND2_X1   g418(.A1(new_n579), .A2(new_n587), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n605), .A2(new_n596), .A3(new_n594), .A4(new_n585), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n595), .A2(KEYINPUT88), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n604), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  AND3_X1   g422(.A1(new_n570), .A2(KEYINPUT93), .A3(KEYINPUT7), .ZN(new_n609));
  AOI21_X1  g423(.A(KEYINPUT93), .B1(new_n570), .B2(KEYINPUT7), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  XOR2_X1   g425(.A(new_n590), .B(KEYINPUT8), .Z(new_n612));
  NOR2_X1   g426(.A1(new_n360), .A2(new_n584), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(KEYINPUT92), .ZN(new_n614));
  OR2_X1    g428(.A1(new_n580), .A2(KEYINPUT91), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n580), .A2(KEYINPUT91), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n615), .A2(new_n583), .A3(new_n616), .ZN(new_n617));
  AND3_X1   g431(.A1(new_n617), .A2(new_n247), .A3(new_n360), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n612), .B1(new_n614), .B2(new_n618), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n608), .A2(new_n572), .A3(new_n611), .A4(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n322), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n563), .B1(new_n602), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n606), .A2(new_n607), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n600), .B1(new_n623), .B2(new_n599), .ZN(new_n624));
  INV_X1    g438(.A(new_n601), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n573), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n626), .A2(new_n322), .A3(new_n562), .A4(new_n620), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n561), .B1(new_n622), .B2(new_n627), .ZN(new_n628));
  AND4_X1   g442(.A1(new_n329), .A2(new_n528), .A3(new_n559), .A4(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(new_n354), .ZN(G3));
  INV_X1    g444(.A(new_n332), .ZN(new_n631));
  INV_X1    g445(.A(new_n420), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n398), .A2(new_n411), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n633), .A2(new_n413), .A3(new_n322), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n631), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n306), .A2(new_n322), .A3(new_n309), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(G472), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n635), .A2(new_n637), .A3(new_n310), .A4(new_n559), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT33), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n640), .A2(KEYINPUT102), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n640), .A2(KEYINPUT102), .ZN(new_n643));
  INV_X1    g457(.A(new_n521), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n518), .B1(new_n513), .B2(new_n515), .ZN(new_n645));
  OAI211_X1 g459(.A(new_n642), .B(new_n643), .C1(new_n644), .C2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT102), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n520), .A2(new_n521), .A3(new_n647), .A4(KEYINPUT33), .ZN(new_n648));
  AOI21_X1  g462(.A(G902), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n522), .A2(new_n523), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT103), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n522), .A2(KEYINPUT103), .A3(new_n523), .ZN(new_n653));
  AOI22_X1  g467(.A1(new_n649), .A2(G478), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n654), .A2(new_n473), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n656), .A2(new_n480), .ZN(new_n657));
  AND3_X1   g471(.A1(new_n622), .A2(KEYINPUT101), .A3(new_n627), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n560), .B1(new_n627), .B2(KEYINPUT101), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n639), .A2(new_n657), .A3(new_n660), .ZN(new_n661));
  XOR2_X1   g475(.A(new_n661), .B(KEYINPUT104), .Z(new_n662));
  XNOR2_X1  g476(.A(KEYINPUT34), .B(G104), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G6));
  NAND2_X1  g478(.A1(new_n473), .A2(new_n525), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n665), .A2(new_n480), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n639), .A2(new_n660), .A3(new_n666), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT35), .B(G107), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G9));
  NOR2_X1   g483(.A1(new_n550), .A2(KEYINPUT36), .ZN(new_n670));
  XOR2_X1   g484(.A(new_n545), .B(new_n670), .Z(new_n671));
  INV_X1    g485(.A(new_n558), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n554), .A2(new_n555), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n673), .B1(new_n674), .B2(new_n529), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT105), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g491(.A(KEYINPUT105), .B1(new_n556), .B2(new_n673), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n527), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n635), .A2(new_n679), .A3(new_n628), .A4(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n637), .A2(new_n310), .ZN(new_n682));
  OR2_X1    g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  XOR2_X1   g497(.A(KEYINPUT37), .B(G110), .Z(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G12));
  AND2_X1   g499(.A1(new_n329), .A2(new_n635), .ZN(new_n686));
  INV_X1    g500(.A(G900), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n476), .B1(new_n477), .B2(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n665), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n686), .A2(new_n660), .A3(new_n679), .A4(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G128), .ZN(G30));
  XNOR2_X1  g505(.A(new_n688), .B(KEYINPUT39), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n635), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n560), .B1(new_n694), .B2(KEYINPUT40), .ZN(new_n695));
  NOR3_X1   g509(.A1(new_n695), .A2(new_n526), .A3(new_n473), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n694), .A2(KEYINPUT40), .ZN(new_n697));
  INV_X1    g511(.A(new_n675), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n272), .A2(new_n303), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n322), .B1(new_n319), .B2(new_n285), .ZN(new_n700));
  OAI21_X1  g514(.A(G472), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n312), .A2(new_n328), .A3(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT106), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n312), .A2(KEYINPUT106), .A3(new_n328), .A4(new_n701), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n698), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n622), .A2(new_n627), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(KEYINPUT38), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n696), .A2(new_n697), .A3(new_n706), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G143), .ZN(G45));
  NAND4_X1  g524(.A1(new_n660), .A2(new_n329), .A3(new_n635), .A4(new_n679), .ZN(new_n711));
  NOR3_X1   g525(.A1(new_n654), .A2(new_n473), .A3(new_n688), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(new_n187), .ZN(G48));
  NOR2_X1   g529(.A1(new_n413), .A2(KEYINPUT107), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n717), .B1(new_n633), .B2(new_n322), .ZN(new_n718));
  AOI211_X1 g532(.A(G902), .B(new_n716), .C1(new_n398), .C2(new_n411), .ZN(new_n719));
  NOR3_X1   g533(.A1(new_n718), .A2(new_n719), .A3(new_n631), .ZN(new_n720));
  AND3_X1   g534(.A1(new_n660), .A2(new_n329), .A3(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n721), .A2(new_n559), .A3(new_n657), .ZN(new_n722));
  XNOR2_X1  g536(.A(KEYINPUT41), .B(G113), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(G15));
  NAND3_X1  g538(.A1(new_n721), .A2(new_n559), .A3(new_n666), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G116), .ZN(G18));
  NAND3_X1  g540(.A1(new_n721), .A2(new_n680), .A3(new_n679), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G119), .ZN(G21));
  INV_X1    g542(.A(new_n307), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n320), .B1(new_n313), .B2(new_n316), .ZN(new_n730));
  AOI22_X1  g544(.A1(new_n730), .A2(new_n303), .B1(new_n286), .B2(new_n292), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n291), .A2(KEYINPUT31), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n729), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n733), .B1(new_n636), .B2(G472), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n720), .A2(new_n734), .A3(new_n559), .A4(new_n481), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n622), .A2(KEYINPUT101), .A3(new_n627), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n602), .A2(new_n621), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT101), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n737), .A2(new_n738), .A3(new_n562), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n473), .A2(new_n526), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n736), .A2(new_n739), .A3(new_n560), .A4(new_n740), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n735), .A2(new_n741), .ZN(new_n742));
  XOR2_X1   g556(.A(new_n742), .B(G122), .Z(G24));
  AOI211_X1 g557(.A(new_n675), .B(new_n733), .C1(new_n636), .C2(G472), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n660), .A2(new_n744), .A3(new_n712), .A4(new_n720), .ZN(new_n745));
  XNOR2_X1  g559(.A(KEYINPUT108), .B(G125), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n745), .B(new_n746), .ZN(G27));
  NAND3_X1  g561(.A1(new_n622), .A2(new_n560), .A3(new_n627), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n421), .A2(new_n748), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n749), .A2(new_n329), .A3(new_n559), .A4(new_n712), .ZN(new_n750));
  NAND2_X1  g564(.A1(KEYINPUT109), .A2(KEYINPUT42), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  XOR2_X1   g566(.A(KEYINPUT109), .B(KEYINPUT42), .Z(new_n753));
  OAI21_X1  g567(.A(new_n752), .B1(new_n750), .B2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G131), .ZN(G33));
  NAND4_X1  g569(.A1(new_n749), .A2(new_n329), .A3(new_n559), .A4(new_n689), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT110), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n756), .B(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G134), .ZN(G36));
  INV_X1    g573(.A(new_n654), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(new_n473), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT111), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n762), .A2(KEYINPUT43), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  AOI22_X1  g578(.A1(new_n760), .A2(new_n473), .B1(new_n762), .B2(KEYINPUT43), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n764), .B1(new_n765), .B2(new_n763), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n766), .A2(new_n682), .A3(new_n698), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(KEYINPUT44), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n748), .B(KEYINPUT112), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(new_n770), .ZN(new_n771));
  OR2_X1    g585(.A1(new_n771), .A2(KEYINPUT113), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n419), .B(KEYINPUT45), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(G469), .ZN(new_n774));
  INV_X1    g588(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n413), .A2(new_n322), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(KEYINPUT46), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(new_n634), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n777), .A2(KEYINPUT46), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n332), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  OR2_X1    g595(.A1(new_n781), .A2(new_n692), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n771), .A2(KEYINPUT113), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n772), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G137), .ZN(G39));
  XNOR2_X1  g600(.A(new_n781), .B(KEYINPUT47), .ZN(new_n787));
  NOR3_X1   g601(.A1(new_n787), .A2(new_n713), .A3(new_n748), .ZN(new_n788));
  INV_X1    g602(.A(new_n329), .ZN(new_n789));
  INV_X1    g603(.A(new_n559), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n788), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G140), .ZN(G42));
  NAND2_X1  g606(.A1(new_n704), .A2(new_n705), .ZN(new_n793));
  NOR3_X1   g607(.A1(new_n793), .A2(new_n708), .A3(new_n761), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n718), .A2(new_n719), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n796), .A2(KEYINPUT49), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n796), .A2(KEYINPUT49), .ZN(new_n798));
  NOR4_X1   g612(.A1(new_n797), .A2(new_n798), .A3(new_n561), .A4(new_n631), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n794), .A2(new_n559), .A3(new_n799), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n787), .B1(new_n332), .B2(new_n796), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n766), .A2(new_n476), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n734), .A2(new_n559), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n805), .A2(new_n769), .ZN(new_n806));
  INV_X1    g620(.A(new_n720), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n559), .A2(new_n476), .ZN(new_n808));
  NOR4_X1   g622(.A1(new_n793), .A2(new_n807), .A3(new_n748), .A4(new_n808), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n654), .A2(new_n473), .ZN(new_n810));
  AOI22_X1  g624(.A1(new_n801), .A2(new_n806), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n807), .A2(new_n748), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n802), .A2(new_n744), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  NOR4_X1   g628(.A1(new_n804), .A2(new_n560), .A3(new_n708), .A4(new_n807), .ZN(new_n815));
  XOR2_X1   g629(.A(new_n815), .B(KEYINPUT50), .Z(new_n816));
  AOI21_X1  g630(.A(new_n814), .B1(KEYINPUT119), .B2(new_n816), .ZN(new_n817));
  OR2_X1    g631(.A1(new_n816), .A2(KEYINPUT119), .ZN(new_n818));
  AOI21_X1  g632(.A(KEYINPUT51), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(new_n689), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n745), .B1(new_n711), .B2(new_n820), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n821), .A2(new_n714), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT115), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n741), .A2(new_n421), .A3(new_n688), .ZN(new_n824));
  AND3_X1   g638(.A1(new_n706), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n823), .B1(new_n706), .B2(new_n824), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n822), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT52), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n822), .B(KEYINPUT52), .C1(new_n825), .C2(new_n826), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n665), .B1(new_n654), .B2(new_n473), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n832), .A2(new_n628), .A3(new_n481), .ZN(new_n833));
  OAI22_X1  g647(.A1(new_n681), .A2(new_n682), .B1(new_n638), .B2(new_n833), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n834), .A2(new_n629), .A3(new_n742), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT114), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n744), .A2(new_n712), .ZN(new_n837));
  INV_X1    g651(.A(new_n749), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n836), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n744), .A2(new_n749), .A3(KEYINPUT114), .A4(new_n712), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n721), .B(new_n559), .C1(new_n657), .C2(new_n666), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n835), .A2(new_n727), .A3(new_n841), .A4(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n679), .A2(new_n526), .A3(new_n473), .ZN(new_n844));
  OR4_X1    g658(.A1(new_n789), .A2(new_n838), .A3(new_n844), .A4(new_n688), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n758), .A2(new_n754), .A3(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n831), .A2(KEYINPUT53), .A3(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT116), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n849), .A2(new_n828), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n686), .A2(new_n660), .A3(new_n679), .A4(new_n712), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n690), .A2(new_n851), .A3(new_n745), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n793), .A2(new_n675), .A3(new_n824), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(KEYINPUT115), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n706), .A2(new_n823), .A3(new_n824), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n852), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT117), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n850), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  OAI211_X1 g672(.A(new_n827), .B(KEYINPUT117), .C1(new_n849), .C2(new_n828), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n830), .A2(new_n849), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n861), .A2(new_n847), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n848), .B1(new_n862), .B2(KEYINPUT53), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(KEYINPUT54), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT54), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n861), .A2(KEYINPUT53), .A3(new_n847), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT118), .ZN(new_n867));
  AOI211_X1 g681(.A(new_n867), .B(KEYINPUT53), .C1(new_n831), .C2(new_n847), .ZN(new_n868));
  INV_X1    g682(.A(new_n830), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n854), .A2(new_n855), .ZN(new_n870));
  AOI21_X1  g684(.A(KEYINPUT52), .B1(new_n870), .B2(new_n822), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n847), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT53), .ZN(new_n873));
  AOI21_X1  g687(.A(KEYINPUT118), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n865), .B(new_n866), .C1(new_n868), .C2(new_n874), .ZN(new_n875));
  NOR4_X1   g689(.A1(new_n804), .A2(new_n659), .A3(new_n658), .A4(new_n807), .ZN(new_n876));
  AOI211_X1 g690(.A(new_n475), .B(new_n876), .C1(new_n655), .C2(new_n809), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n864), .A2(new_n875), .A3(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT51), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n814), .A2(new_n879), .A3(new_n816), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n789), .A2(new_n790), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n802), .A2(new_n881), .A3(new_n812), .ZN(new_n882));
  XOR2_X1   g696(.A(new_n882), .B(KEYINPUT48), .Z(new_n883));
  NOR4_X1   g697(.A1(new_n819), .A2(new_n878), .A3(new_n880), .A4(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(G952), .A2(G953), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n800), .B1(new_n884), .B2(new_n885), .ZN(G75));
  NOR2_X1   g700(.A1(new_n624), .A2(new_n625), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(new_n574), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(new_n626), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n889), .B(KEYINPUT55), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT56), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n891), .B1(KEYINPUT120), .B2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n866), .B1(new_n868), .B2(new_n874), .ZN(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n896), .A2(new_n322), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(G210), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n894), .B1(new_n898), .B2(new_n892), .ZN(new_n899));
  AOI211_X1 g713(.A(KEYINPUT56), .B(new_n893), .C1(new_n897), .C2(G210), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n333), .A2(G952), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(G51));
  NAND2_X1  g716(.A1(new_n895), .A2(KEYINPUT54), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n903), .A2(KEYINPUT121), .A3(new_n875), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT121), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n895), .A2(new_n905), .A3(KEYINPUT54), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT57), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n776), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n904), .A2(new_n906), .A3(new_n908), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n776), .A2(new_n907), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n633), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n897), .A2(new_n775), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n901), .B1(new_n911), .B2(new_n912), .ZN(G54));
  NAND3_X1  g727(.A1(new_n897), .A2(KEYINPUT58), .A3(G475), .ZN(new_n914));
  INV_X1    g728(.A(new_n467), .ZN(new_n915));
  AND2_X1   g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n914), .A2(new_n915), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n916), .A2(new_n917), .A3(new_n901), .ZN(G60));
  NAND2_X1  g732(.A1(new_n646), .A2(new_n648), .ZN(new_n919));
  NAND2_X1  g733(.A1(G478), .A2(G902), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(KEYINPUT59), .ZN(new_n921));
  AND2_X1   g735(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n904), .A2(new_n906), .A3(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(new_n901), .ZN(new_n924));
  AND3_X1   g738(.A1(new_n923), .A2(KEYINPUT122), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(KEYINPUT122), .B1(new_n923), .B2(new_n924), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n864), .A2(new_n875), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n919), .B1(new_n927), .B2(new_n921), .ZN(new_n928));
  NOR3_X1   g742(.A1(new_n925), .A2(new_n926), .A3(new_n928), .ZN(G63));
  NAND2_X1  g743(.A1(G217), .A2(G902), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT60), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n671), .B(KEYINPUT123), .ZN(new_n932));
  OR3_X1    g746(.A1(new_n896), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(new_n557), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n934), .B1(new_n896), .B2(new_n931), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n933), .A2(new_n924), .A3(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT61), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n936), .B(new_n937), .ZN(G66));
  OAI21_X1  g752(.A(G953), .B1(new_n479), .B2(new_n565), .ZN(new_n939));
  AND3_X1   g753(.A1(new_n835), .A2(new_n727), .A3(new_n842), .ZN(new_n940));
  INV_X1    g754(.A(new_n333), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n939), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n887), .B1(G898), .B2(new_n333), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n942), .B(new_n943), .ZN(G69));
  OAI21_X1  g758(.A(new_n456), .B1(new_n457), .B2(new_n432), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n289), .B(new_n945), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(KEYINPUT124), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n881), .A2(new_n693), .A3(new_n749), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n949), .B1(new_n656), .B2(new_n665), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(KEYINPUT125), .ZN(new_n951));
  OR2_X1    g765(.A1(new_n950), .A2(KEYINPUT125), .ZN(new_n952));
  AND4_X1   g766(.A1(new_n785), .A2(new_n791), .A3(new_n951), .A4(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n709), .A2(new_n822), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT62), .Z(new_n955));
  NAND2_X1  g769(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n948), .B1(new_n956), .B2(new_n333), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n941), .A2(G900), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n758), .A2(new_n754), .ZN(new_n959));
  NOR3_X1   g773(.A1(new_n789), .A2(new_n790), .A3(new_n741), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n959), .B1(new_n783), .B2(new_n960), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n791), .A2(new_n785), .A3(new_n822), .A4(new_n961), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n946), .B(new_n958), .C1(new_n962), .C2(new_n941), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n963), .A2(KEYINPUT126), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n957), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n333), .B1(G227), .B2(G900), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(new_n966), .ZN(new_n968));
  NOR3_X1   g782(.A1(new_n957), .A2(new_n964), .A3(new_n968), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n967), .A2(new_n969), .ZN(G72));
  INV_X1    g784(.A(new_n699), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n953), .A2(new_n940), .A3(new_n955), .ZN(new_n972));
  XNOR2_X1  g786(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n973));
  NAND2_X1  g787(.A1(G472), .A2(G902), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n973), .B(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n971), .B1(new_n972), .B2(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(new_n940), .ZN(new_n977));
  OR2_X1    g791(.A1(new_n962), .A2(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n323), .B1(new_n978), .B2(new_n975), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n863), .A2(new_n323), .A3(new_n971), .A4(new_n975), .ZN(new_n980));
  INV_X1    g794(.A(new_n980), .ZN(new_n981));
  NOR4_X1   g795(.A1(new_n976), .A2(new_n979), .A3(new_n901), .A4(new_n981), .ZN(G57));
endmodule


