//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 0 1 1 1 1 1 0 0 1 0 0 0 0 0 1 0 0 0 1 0 0 0 1 1 0 1 0 1 1 1 0 0 0 0 1 1 0 1 1 0 0 0 1 1 1 0 0 1 1 0 1 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:50 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n447, new_n449, new_n451, new_n452, new_n454,
    new_n455, new_n457, new_n458, new_n459, new_n460, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n560, new_n562, new_n563, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n577, new_n578, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n619, new_n620, new_n623, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1182, new_n1183;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT64), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  NAND2_X1  g021(.A1(G94), .A2(G452), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT65), .Z(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  INV_X1    g025(.A(G567), .ZN(new_n451));
  NOR2_X1   g026(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT66), .ZN(G234));
  INV_X1    g028(.A(G2106), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n449), .A2(new_n454), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT67), .Z(G217));
  NAND4_X1  g031(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT2), .Z(new_n458));
  NOR4_X1   g033(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G325));
  XOR2_X1   g036(.A(new_n460), .B(KEYINPUT68), .Z(G261));
  OAI22_X1  g037(.A1(new_n458), .A2(new_n454), .B1(new_n451), .B2(new_n459), .ZN(new_n463));
  XNOR2_X1  g038(.A(new_n463), .B(KEYINPUT69), .ZN(G319));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n467), .A2(new_n469), .A3(G125), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n465), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n467), .A2(new_n469), .A3(G137), .ZN(new_n473));
  NAND2_X1  g048(.A1(G101), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(G2105), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n472), .A2(new_n475), .ZN(G160));
  NAND2_X1  g051(.A1(new_n467), .A2(new_n469), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n477), .A2(new_n465), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n477), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  NOR2_X1   g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI21_X1  g057(.A(G2104), .B1(new_n465), .B2(G112), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n479), .B(new_n481), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  XOR2_X1   g059(.A(new_n484), .B(KEYINPUT70), .Z(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  AND3_X1   g061(.A1(KEYINPUT71), .A2(KEYINPUT4), .A3(G138), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n487), .A2(new_n467), .A3(new_n469), .ZN(new_n488));
  NAND2_X1  g063(.A1(G102), .A2(G2104), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(new_n465), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n467), .A2(new_n469), .A3(G126), .ZN(new_n492));
  NAND2_X1  g067(.A1(G114), .A2(G2104), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G2105), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n467), .A2(new_n469), .A3(G138), .A4(new_n465), .ZN(new_n496));
  NAND2_X1  g071(.A1(KEYINPUT71), .A2(KEYINPUT4), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n491), .A2(new_n495), .A3(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  INV_X1    g075(.A(KEYINPUT6), .ZN(new_n501));
  INV_X1    g076(.A(G651), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT72), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT72), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G651), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n501), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n502), .A2(KEYINPUT6), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n508), .A2(G50), .A3(G543), .ZN(new_n509));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n510), .A2(KEYINPUT5), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT5), .ZN(new_n512));
  OAI21_X1  g087(.A(KEYINPUT73), .B1(new_n512), .B2(G543), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT73), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n514), .A2(new_n510), .A3(KEYINPUT5), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n511), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n508), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(G88), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n509), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n516), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n520));
  XNOR2_X1  g095(.A(KEYINPUT72), .B(G651), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n519), .A2(new_n523), .ZN(G166));
  OAI21_X1  g099(.A(KEYINPUT74), .B1(new_n506), .B2(new_n507), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT74), .ZN(new_n526));
  INV_X1    g101(.A(new_n507), .ZN(new_n527));
  OAI211_X1 g102(.A(new_n526), .B(new_n527), .C1(new_n521), .C2(new_n501), .ZN(new_n528));
  AND3_X1   g103(.A1(new_n525), .A2(G543), .A3(new_n528), .ZN(new_n529));
  XNOR2_X1  g104(.A(KEYINPUT75), .B(G51), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AND2_X1   g106(.A1(G76), .A2(G543), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n516), .A2(G63), .B1(KEYINPUT7), .B2(new_n532), .ZN(new_n533));
  OR2_X1    g108(.A1(new_n533), .A2(new_n502), .ZN(new_n534));
  AOI21_X1  g109(.A(KEYINPUT7), .B1(new_n532), .B2(G651), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n504), .A2(G651), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n502), .A2(KEYINPUT72), .ZN(new_n537));
  OAI21_X1  g112(.A(KEYINPUT6), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  AND3_X1   g113(.A1(new_n516), .A2(new_n538), .A3(new_n527), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n535), .B1(new_n539), .B2(G89), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n531), .A2(new_n534), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(KEYINPUT76), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT76), .ZN(new_n543));
  NAND4_X1  g118(.A1(new_n531), .A2(new_n543), .A3(new_n534), .A4(new_n540), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n542), .A2(new_n544), .ZN(G168));
  NAND2_X1  g120(.A1(new_n529), .A2(G52), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n516), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n547));
  OR2_X1    g122(.A1(new_n547), .A2(new_n522), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n539), .A2(G90), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n546), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(G171));
  NAND2_X1  g126(.A1(new_n529), .A2(G43), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n516), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n553));
  OR2_X1    g128(.A1(new_n553), .A2(new_n522), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n539), .A2(G81), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n552), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(new_n558));
  XOR2_X1   g133(.A(new_n558), .B(KEYINPUT77), .Z(G153));
  AND3_X1   g134(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G36), .ZN(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n560), .A2(new_n563), .ZN(G188));
  AND2_X1   g139(.A1(new_n525), .A2(new_n528), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT9), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n565), .A2(new_n566), .A3(G53), .A4(G543), .ZN(new_n567));
  NAND4_X1  g142(.A1(new_n525), .A2(G53), .A3(G543), .A4(new_n528), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(KEYINPUT9), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n516), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n571), .A2(new_n502), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n516), .A2(new_n538), .A3(G91), .A4(new_n527), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n570), .A2(new_n575), .ZN(G299));
  INV_X1    g151(.A(KEYINPUT78), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n550), .B(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(G301));
  INV_X1    g154(.A(G168), .ZN(G286));
  OR2_X1    g155(.A1(new_n519), .A2(new_n523), .ZN(G303));
  INV_X1    g156(.A(KEYINPUT79), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n529), .A2(new_n582), .A3(G49), .ZN(new_n583));
  OR2_X1    g158(.A1(new_n516), .A2(G74), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n539), .A2(G87), .B1(new_n584), .B2(G651), .ZN(new_n585));
  NAND4_X1  g160(.A1(new_n525), .A2(G49), .A3(G543), .A4(new_n528), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(KEYINPUT79), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n583), .A2(new_n585), .A3(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT80), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n586), .B(new_n582), .ZN(new_n591));
  AOI21_X1  g166(.A(KEYINPUT80), .B1(new_n591), .B2(new_n585), .ZN(new_n592));
  OR2_X1    g167(.A1(new_n590), .A2(new_n592), .ZN(G288));
  NAND3_X1  g168(.A1(new_n508), .A2(G48), .A3(G543), .ZN(new_n594));
  INV_X1    g169(.A(G86), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n517), .B2(new_n595), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n516), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n597), .A2(new_n522), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(G305));
  AND2_X1   g175(.A1(new_n529), .A2(G47), .ZN(new_n601));
  INV_X1    g176(.A(G85), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n516), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n603));
  OAI22_X1  g178(.A1(new_n517), .A2(new_n602), .B1(new_n603), .B2(new_n522), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(G290));
  NAND2_X1  g181(.A1(G301), .A2(G868), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n539), .A2(G92), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT10), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n608), .B(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n529), .A2(G54), .ZN(new_n611));
  AND2_X1   g186(.A1(new_n516), .A2(G66), .ZN(new_n612));
  AND2_X1   g187(.A1(G79), .A2(G543), .ZN(new_n613));
  OAI21_X1  g188(.A(G651), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n610), .A2(new_n611), .A3(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n607), .B1(G868), .B2(new_n616), .ZN(G284));
  OAI21_X1  g192(.A(new_n607), .B1(G868), .B2(new_n616), .ZN(G321));
  NAND2_X1  g193(.A1(G286), .A2(G868), .ZN(new_n619));
  INV_X1    g194(.A(G299), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(G868), .B2(new_n620), .ZN(G297));
  OAI21_X1  g196(.A(new_n619), .B1(G868), .B2(new_n620), .ZN(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n616), .B1(new_n623), .B2(G860), .ZN(G148));
  NAND2_X1  g199(.A1(new_n616), .A2(new_n623), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(G868), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(G868), .B2(new_n557), .ZN(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g203(.A1(new_n465), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(KEYINPUT12), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT13), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(G2100), .Z(new_n632));
  AOI22_X1  g207(.A1(G123), .A2(new_n478), .B1(new_n480), .B2(G135), .ZN(new_n633));
  OAI21_X1  g208(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n634));
  INV_X1    g209(.A(KEYINPUT81), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n634), .A2(new_n635), .ZN(new_n637));
  OAI211_X1 g212(.A(new_n636), .B(new_n637), .C1(G111), .C2(new_n465), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n633), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(G2096), .Z(new_n640));
  NAND2_X1  g215(.A1(new_n632), .A2(new_n640), .ZN(G156));
  XOR2_X1   g216(.A(KEYINPUT15), .B(G2435), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2438), .ZN(new_n643));
  XOR2_X1   g218(.A(G2427), .B(G2430), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT82), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n643), .B(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n646), .A2(KEYINPUT14), .ZN(new_n647));
  XOR2_X1   g222(.A(G2451), .B(G2454), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT16), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n647), .B(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(G1341), .B(G1348), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2443), .B(G2446), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n652), .B(new_n653), .Z(new_n654));
  AND2_X1   g229(.A1(new_n654), .A2(G14), .ZN(G401));
  XOR2_X1   g230(.A(G2084), .B(G2090), .Z(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G2067), .B(G2678), .Z(new_n658));
  OR2_X1    g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n657), .A2(new_n658), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n659), .A2(new_n660), .A3(KEYINPUT17), .ZN(new_n661));
  INV_X1    g236(.A(KEYINPUT18), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G2072), .B(G2078), .Z(new_n664));
  AOI21_X1  g239(.A(new_n664), .B1(new_n659), .B2(KEYINPUT18), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n663), .B(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G2096), .B(G2100), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT83), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n666), .B(new_n668), .ZN(G227));
  XOR2_X1   g244(.A(G1961), .B(G1966), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT84), .ZN(new_n671));
  XOR2_X1   g246(.A(G1956), .B(G2474), .Z(new_n672));
  NOR2_X1   g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1971), .B(G1976), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT19), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT85), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n671), .A2(new_n672), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n679), .A2(new_n676), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n680), .B(KEYINPUT20), .Z(new_n681));
  NAND3_X1  g256(.A1(new_n674), .A2(new_n679), .A3(new_n676), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n678), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1991), .B(G1996), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT86), .B(G1986), .ZN(new_n688));
  INV_X1    g263(.A(G1981), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n687), .B(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(G229));
  INV_X1    g267(.A(G29), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(G35), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n694), .B1(G162), .B2(new_n693), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT29), .Z(new_n696));
  INV_X1    g271(.A(G2090), .ZN(new_n697));
  OR2_X1    g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  OR2_X1    g273(.A1(G16), .A2(G22), .ZN(new_n699));
  INV_X1    g274(.A(G16), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n699), .B1(G303), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(KEYINPUT90), .ZN(new_n702));
  INV_X1    g277(.A(KEYINPUT90), .ZN(new_n703));
  OAI211_X1 g278(.A(new_n703), .B(new_n699), .C1(G303), .C2(new_n700), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(G1971), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n588), .A2(KEYINPUT89), .ZN(new_n708));
  INV_X1    g283(.A(KEYINPUT89), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n591), .A2(new_n709), .A3(new_n585), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G16), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(G16), .B2(G23), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT33), .B(G1976), .Z(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  OAI211_X1 g291(.A(new_n712), .B(new_n714), .C1(G16), .C2(G23), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n700), .A2(G6), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(new_n599), .B2(new_n700), .ZN(new_n719));
  XOR2_X1   g294(.A(KEYINPUT32), .B(G1981), .Z(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  NAND4_X1  g296(.A1(new_n707), .A2(new_n716), .A3(new_n717), .A4(new_n721), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n722), .A2(KEYINPUT34), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n722), .A2(KEYINPUT34), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT91), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n722), .A2(KEYINPUT91), .A3(KEYINPUT34), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n723), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(G24), .ZN(new_n729));
  OAI21_X1  g304(.A(KEYINPUT87), .B1(new_n729), .B2(G16), .ZN(new_n730));
  OR3_X1    g305(.A1(new_n729), .A2(KEYINPUT87), .A3(G16), .ZN(new_n731));
  OAI211_X1 g306(.A(new_n730), .B(new_n731), .C1(new_n605), .C2(new_n700), .ZN(new_n732));
  XOR2_X1   g307(.A(KEYINPUT88), .B(G1986), .Z(new_n733));
  XNOR2_X1  g308(.A(new_n732), .B(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n478), .A2(G119), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n480), .A2(G131), .ZN(new_n736));
  NOR2_X1   g311(.A1(G95), .A2(G2105), .ZN(new_n737));
  OAI21_X1  g312(.A(G2104), .B1(new_n465), .B2(G107), .ZN(new_n738));
  OAI211_X1 g313(.A(new_n735), .B(new_n736), .C1(new_n737), .C2(new_n738), .ZN(new_n739));
  MUX2_X1   g314(.A(G25), .B(new_n739), .S(G29), .Z(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT35), .B(G1991), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(new_n742), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n728), .A2(new_n734), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(KEYINPUT36), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT36), .ZN(new_n746));
  NAND4_X1  g321(.A1(new_n728), .A2(new_n746), .A3(new_n734), .A4(new_n743), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g323(.A1(G29), .A2(G33), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT94), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT25), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n480), .A2(G139), .ZN(new_n753));
  INV_X1    g328(.A(new_n477), .ZN(new_n754));
  AOI22_X1  g329(.A1(new_n754), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n755));
  OAI211_X1 g330(.A(new_n752), .B(new_n753), .C1(new_n465), .C2(new_n755), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT95), .Z(new_n757));
  AOI21_X1  g332(.A(new_n749), .B1(new_n757), .B2(G29), .ZN(new_n758));
  INV_X1    g333(.A(G2072), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n480), .A2(G141), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n478), .A2(G129), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n465), .A2(G105), .A3(G2104), .ZN(new_n763));
  NAND3_X1  g338(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT26), .Z(new_n765));
  NAND4_X1  g340(.A1(new_n761), .A2(new_n762), .A3(new_n763), .A4(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n767), .A2(G29), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G29), .B2(G32), .ZN(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT27), .B(G1996), .ZN(new_n770));
  INV_X1    g345(.A(G34), .ZN(new_n771));
  AND2_X1   g346(.A1(new_n771), .A2(KEYINPUT24), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n771), .A2(KEYINPUT24), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n693), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G160), .B2(new_n693), .ZN(new_n775));
  AOI22_X1  g350(.A1(new_n769), .A2(new_n770), .B1(G2084), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n760), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT96), .ZN(new_n778));
  AND2_X1   g353(.A1(new_n693), .A2(G26), .ZN(new_n779));
  OR2_X1    g354(.A1(G104), .A2(G2105), .ZN(new_n780));
  OAI211_X1 g355(.A(new_n780), .B(G2104), .C1(G116), .C2(new_n465), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT92), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n478), .A2(G128), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n480), .A2(G140), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n782), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT93), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n779), .B1(new_n786), .B2(G29), .ZN(new_n787));
  MUX2_X1   g362(.A(new_n779), .B(new_n787), .S(KEYINPUT28), .Z(new_n788));
  INV_X1    g363(.A(G2067), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n775), .A2(G2084), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(KEYINPUT97), .Z(new_n792));
  NOR2_X1   g367(.A1(G27), .A2(G29), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(G164), .B2(G29), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n794), .A2(G2078), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT30), .ZN(new_n796));
  OR2_X1    g371(.A1(new_n796), .A2(G28), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n796), .A2(G28), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n797), .A2(new_n798), .A3(new_n693), .ZN(new_n799));
  AND2_X1   g374(.A1(new_n795), .A2(new_n799), .ZN(new_n800));
  OAI221_X1 g375(.A(new_n800), .B1(new_n693), .B2(new_n639), .C1(new_n769), .C2(new_n770), .ZN(new_n801));
  NAND2_X1  g376(.A1(G171), .A2(G16), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(G5), .B2(G16), .ZN(new_n803));
  INV_X1    g378(.A(G1961), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(G2078), .B2(new_n794), .ZN(new_n806));
  AOI211_X1 g381(.A(new_n801), .B(new_n806), .C1(new_n696), .C2(new_n697), .ZN(new_n807));
  NAND4_X1  g382(.A1(new_n778), .A2(new_n790), .A3(new_n792), .A4(new_n807), .ZN(new_n808));
  XOR2_X1   g383(.A(KEYINPUT31), .B(G11), .Z(new_n809));
  NOR2_X1   g384(.A1(new_n788), .A2(new_n789), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n700), .A2(G4), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(new_n616), .B2(new_n700), .ZN(new_n812));
  INV_X1    g387(.A(G1348), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(G16), .A2(G21), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(G168), .B2(G16), .ZN(new_n816));
  INV_X1    g391(.A(G1966), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n700), .A2(KEYINPUT23), .A3(G20), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT23), .ZN(new_n820));
  INV_X1    g395(.A(G20), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n820), .B1(new_n821), .B2(G16), .ZN(new_n822));
  OAI211_X1 g397(.A(new_n819), .B(new_n822), .C1(new_n620), .C2(new_n700), .ZN(new_n823));
  INV_X1    g398(.A(G1956), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n823), .B(new_n824), .ZN(new_n825));
  OR2_X1    g400(.A1(new_n803), .A2(new_n804), .ZN(new_n826));
  NAND4_X1  g401(.A1(new_n814), .A2(new_n818), .A3(new_n825), .A4(new_n826), .ZN(new_n827));
  NOR4_X1   g402(.A1(new_n808), .A2(new_n809), .A3(new_n810), .A4(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n700), .A2(G19), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n829), .B1(new_n557), .B2(new_n700), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n830), .B(G1341), .Z(new_n831));
  AND4_X1   g406(.A1(new_n698), .A2(new_n748), .A3(new_n828), .A4(new_n831), .ZN(G311));
  NAND4_X1  g407(.A1(new_n748), .A2(new_n828), .A3(new_n698), .A4(new_n831), .ZN(G150));
  AOI22_X1  g408(.A1(new_n516), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n834), .A2(new_n522), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT98), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n529), .A2(G55), .ZN(new_n837));
  INV_X1    g412(.A(G93), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n837), .B1(new_n838), .B2(new_n517), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(G860), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n841), .B(KEYINPUT37), .Z(new_n842));
  NAND2_X1  g417(.A1(new_n616), .A2(G559), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT38), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT39), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n840), .A2(KEYINPUT99), .A3(new_n556), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n556), .A2(KEYINPUT99), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n556), .A2(KEYINPUT99), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n836), .A2(new_n839), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  AND2_X1   g425(.A1(new_n846), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n845), .B(new_n851), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n842), .B1(new_n852), .B2(G860), .ZN(G145));
  XOR2_X1   g428(.A(new_n639), .B(G160), .Z(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(new_n485), .ZN(new_n855));
  XNOR2_X1  g430(.A(G164), .B(new_n766), .ZN(new_n856));
  OR2_X1    g431(.A1(new_n786), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n786), .A2(new_n856), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n857), .A2(new_n756), .A3(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n756), .B(KEYINPUT95), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n861), .B1(new_n857), .B2(new_n858), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n630), .B1(new_n860), .B2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n862), .ZN(new_n864));
  INV_X1    g439(.A(new_n630), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n864), .A2(new_n865), .A3(new_n859), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n480), .A2(G142), .ZN(new_n868));
  OR2_X1    g443(.A1(new_n868), .A2(KEYINPUT100), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n478), .A2(G130), .ZN(new_n870));
  OR2_X1    g445(.A1(G106), .A2(G2105), .ZN(new_n871));
  OAI211_X1 g446(.A(new_n871), .B(G2104), .C1(G118), .C2(new_n465), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n868), .A2(KEYINPUT100), .ZN(new_n873));
  NAND4_X1  g448(.A1(new_n869), .A2(new_n870), .A3(new_n872), .A4(new_n873), .ZN(new_n874));
  XOR2_X1   g449(.A(KEYINPUT101), .B(KEYINPUT102), .Z(new_n875));
  XNOR2_X1  g450(.A(new_n874), .B(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(new_n739), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n867), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n863), .A2(new_n866), .A3(new_n877), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n855), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n881), .A2(G37), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n879), .A2(new_n855), .A3(new_n880), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(KEYINPUT103), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT103), .ZN(new_n885));
  NAND4_X1  g460(.A1(new_n879), .A2(new_n885), .A3(new_n855), .A4(new_n880), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n882), .A2(new_n884), .A3(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g463(.A1(G290), .A2(G166), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n605), .A2(G303), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(G305), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n599), .B1(new_n889), .B2(new_n890), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(new_n711), .ZN(new_n895));
  NAND4_X1  g470(.A1(new_n892), .A2(new_n708), .A3(new_n710), .A4(new_n893), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT42), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n897), .B1(KEYINPUT105), .B2(new_n898), .ZN(new_n899));
  AND2_X1   g474(.A1(new_n898), .A2(KEYINPUT105), .ZN(new_n900));
  OR2_X1    g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n851), .B(new_n625), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT104), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n615), .B1(new_n620), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(G299), .A2(KEYINPUT104), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n615), .A2(KEYINPUT104), .A3(G299), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT41), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n906), .A2(KEYINPUT41), .A3(new_n907), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n902), .A2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n908), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n913), .B1(new_n914), .B2(new_n902), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n899), .A2(new_n900), .ZN(new_n916));
  AND3_X1   g491(.A1(new_n901), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n915), .B1(new_n901), .B2(new_n916), .ZN(new_n918));
  OAI21_X1  g493(.A(G868), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n919), .B1(G868), .B2(new_n849), .ZN(G295));
  OAI21_X1  g495(.A(new_n919), .B1(G868), .B2(new_n849), .ZN(G331));
  INV_X1    g496(.A(KEYINPUT107), .ZN(new_n922));
  NAND2_X1  g497(.A1(G286), .A2(new_n550), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n578), .A2(G168), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n851), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n846), .A2(new_n850), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n927), .A2(new_n923), .A3(new_n924), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(new_n914), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n910), .A2(new_n911), .A3(new_n926), .A4(new_n928), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(new_n897), .ZN(new_n933));
  INV_X1    g508(.A(G37), .ZN(new_n934));
  AND2_X1   g509(.A1(new_n895), .A2(new_n896), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n935), .A2(new_n931), .A3(new_n930), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n933), .A2(new_n934), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n922), .B1(new_n937), .B2(KEYINPUT43), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n931), .A2(KEYINPUT106), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n932), .A2(new_n939), .A3(new_n897), .ZN(new_n940));
  OAI211_X1 g515(.A(new_n931), .B(new_n930), .C1(new_n935), .C2(KEYINPUT106), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n940), .A2(new_n941), .A3(new_n934), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n938), .B1(KEYINPUT43), .B2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT44), .ZN(new_n944));
  OR3_X1    g519(.A1(new_n942), .A2(KEYINPUT107), .A3(KEYINPUT43), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n944), .B1(new_n942), .B2(KEYINPUT43), .ZN(new_n947));
  OR2_X1    g522(.A1(new_n937), .A2(KEYINPUT43), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT108), .ZN(new_n949));
  AND3_X1   g524(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n949), .B1(new_n947), .B2(new_n948), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n946), .B1(new_n950), .B2(new_n951), .ZN(G397));
  NOR2_X1   g527(.A1(G290), .A2(G1986), .ZN(new_n953));
  XOR2_X1   g528(.A(new_n953), .B(KEYINPUT110), .Z(new_n954));
  INV_X1    g529(.A(G1384), .ZN(new_n955));
  AOI21_X1  g530(.A(KEYINPUT45), .B1(new_n499), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  XNOR2_X1  g532(.A(KEYINPUT109), .B(G40), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(G160), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n957), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n954), .A2(new_n961), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n962), .B(KEYINPUT48), .ZN(new_n963));
  XNOR2_X1  g538(.A(new_n786), .B(new_n789), .ZN(new_n964));
  INV_X1    g539(.A(G1996), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n766), .B(new_n965), .ZN(new_n966));
  AND2_X1   g541(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  OR2_X1    g542(.A1(new_n739), .A2(new_n741), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n969), .B1(new_n741), .B2(new_n739), .ZN(new_n970));
  INV_X1    g545(.A(new_n961), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n963), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n971), .B1(new_n964), .B2(new_n767), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT46), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n973), .B1(KEYINPUT127), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n961), .A2(new_n965), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n974), .A2(KEYINPUT127), .ZN(new_n977));
  XNOR2_X1  g552(.A(new_n976), .B(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n975), .A2(new_n978), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n979), .B(KEYINPUT47), .ZN(new_n980));
  INV_X1    g555(.A(new_n967), .ZN(new_n981));
  OAI22_X1  g556(.A1(new_n981), .A2(new_n968), .B1(G2067), .B2(new_n786), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n961), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n972), .A2(new_n980), .A3(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT126), .ZN(new_n986));
  NAND2_X1  g561(.A1(G290), .A2(G1986), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n987), .B(KEYINPUT111), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n954), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n971), .B1(new_n970), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n711), .A2(G1976), .ZN(new_n991));
  INV_X1    g566(.A(G1976), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n992), .B1(new_n590), .B2(new_n592), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT52), .ZN(new_n994));
  AOI21_X1  g569(.A(G2105), .B1(new_n488), .B2(new_n489), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n465), .B1(new_n492), .B2(new_n493), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(G1384), .B1(new_n997), .B2(new_n498), .ZN(new_n998));
  NOR3_X1   g573(.A1(new_n472), .A2(new_n475), .A3(new_n958), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(G8), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n991), .A2(new_n993), .A3(new_n994), .A4(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT49), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n599), .A2(new_n689), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n599), .A2(new_n689), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1004), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1007), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1009), .A2(KEYINPUT49), .A3(new_n1005), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1008), .A2(new_n1010), .A3(new_n1002), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n992), .B1(new_n708), .B2(new_n710), .ZN(new_n1012));
  OAI21_X1  g587(.A(KEYINPUT52), .B1(new_n1012), .B2(new_n1001), .ZN(new_n1013));
  AND3_X1   g588(.A1(new_n1003), .A2(new_n1011), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT55), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1015), .B1(G303), .B2(G8), .ZN(new_n1016));
  INV_X1    g591(.A(G8), .ZN(new_n1017));
  NOR3_X1   g592(.A1(G166), .A2(KEYINPUT55), .A3(new_n1017), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n499), .A2(new_n955), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT113), .B1(new_n1020), .B2(KEYINPUT50), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT50), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n960), .B1(new_n998), .B2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1020), .A2(KEYINPUT113), .A3(KEYINPUT50), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1022), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1026), .A2(G2090), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT112), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1028), .B1(new_n998), .B2(KEYINPUT45), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n960), .B1(new_n998), .B2(KEYINPUT45), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT45), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1020), .A2(KEYINPUT112), .A3(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1029), .A2(new_n1030), .A3(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(new_n706), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  OAI211_X1 g610(.A(G8), .B(new_n1019), .C1(new_n1027), .C2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1014), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(new_n992), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1005), .B1(new_n1040), .B2(G288), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(new_n1002), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1038), .A2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n999), .B1(new_n1020), .B2(KEYINPUT50), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n998), .A2(new_n1023), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(new_n697), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1017), .B1(new_n1034), .B2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(KEYINPUT114), .B1(new_n1048), .B2(new_n1019), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1019), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT114), .ZN(new_n1051));
  AOI22_X1  g626(.A1(new_n1033), .A2(new_n706), .B1(new_n1046), .B2(new_n697), .ZN(new_n1052));
  OAI211_X1 g627(.A(new_n1050), .B(new_n1051), .C1(new_n1052), .C2(new_n1017), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1049), .A2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n499), .A2(KEYINPUT45), .A3(new_n955), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n957), .A2(new_n999), .A3(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(new_n817), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1057), .B1(new_n1026), .B2(G2084), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(G8), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1059), .A2(G286), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1014), .A2(new_n1054), .A3(new_n1036), .A4(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT115), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT63), .ZN(new_n1063));
  AND3_X1   g638(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1062), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  AND2_X1   g641(.A1(new_n1014), .A2(new_n1036), .ZN(new_n1067));
  OAI21_X1  g642(.A(G8), .B1(new_n1027), .B2(new_n1035), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1063), .B1(new_n1068), .B2(new_n1050), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1067), .A2(new_n1060), .A3(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1043), .B1(new_n1066), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT122), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1072), .B1(G168), .B2(new_n1017), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n542), .A2(KEYINPUT122), .A3(G8), .A4(new_n544), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(new_n1058), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT123), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1075), .A2(KEYINPUT123), .A3(new_n1058), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  AND2_X1   g655(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(new_n1059), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT51), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT124), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1084), .B1(new_n1058), .B2(G8), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1082), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1081), .A2(new_n1084), .A3(KEYINPUT51), .A4(new_n1059), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1080), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(G2078), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1029), .A2(new_n1030), .A3(new_n1089), .A4(new_n1032), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT53), .ZN(new_n1091));
  AOI22_X1  g666(.A1(new_n1026), .A2(new_n804), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  AND2_X1   g667(.A1(new_n957), .A2(new_n1055), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1091), .A2(G2078), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1093), .A2(new_n999), .A3(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1092), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(new_n578), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT62), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  OR2_X1    g674(.A1(new_n1088), .A2(new_n1099), .ZN(new_n1100));
  AND2_X1   g675(.A1(new_n1067), .A2(new_n1054), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT120), .ZN(new_n1102));
  OAI211_X1 g677(.A(KEYINPUT116), .B(new_n573), .C1(new_n571), .C2(new_n502), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT57), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(new_n569), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n568), .A2(KEYINPUT9), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1105), .B(new_n575), .C1(new_n1106), .C2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1105), .B1(new_n570), .B2(new_n575), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  XNOR2_X1  g686(.A(KEYINPUT56), .B(G2072), .ZN(new_n1112));
  XNOR2_X1  g687(.A(new_n1112), .B(KEYINPUT117), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1029), .A2(new_n1030), .A3(new_n1032), .A4(new_n1113), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n824), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1111), .A2(new_n1116), .ZN(new_n1117));
  OAI211_X1 g692(.A(new_n1115), .B(new_n1114), .C1(new_n1109), .C2(new_n1110), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1102), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT61), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1000), .A2(G2067), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1121), .B1(new_n1026), .B2(new_n813), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n615), .A2(KEYINPUT60), .ZN(new_n1123));
  AOI22_X1  g698(.A1(new_n1119), .A2(new_n1120), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  AND3_X1   g699(.A1(new_n1020), .A2(KEYINPUT113), .A3(KEYINPUT50), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1125), .A2(new_n1021), .ZN(new_n1126));
  AOI21_X1  g701(.A(G1348), .B1(new_n1126), .B2(new_n1024), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n616), .B1(new_n1127), .B2(new_n1121), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1122), .A2(new_n615), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  XNOR2_X1  g705(.A(KEYINPUT118), .B(G1996), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1033), .A2(new_n1131), .ZN(new_n1132));
  XOR2_X1   g707(.A(KEYINPUT58), .B(G1341), .Z(new_n1133));
  NAND2_X1  g708(.A1(new_n1000), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(KEYINPUT119), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT119), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1000), .A2(new_n1136), .A3(new_n1133), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n557), .B1(new_n1132), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(KEYINPUT59), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT59), .ZN(new_n1141));
  OAI211_X1 g716(.A(new_n1141), .B(new_n557), .C1(new_n1132), .C2(new_n1138), .ZN(new_n1142));
  AOI22_X1  g717(.A1(new_n1130), .A2(KEYINPUT60), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(KEYINPUT120), .ZN(new_n1145));
  AOI21_X1  g720(.A(KEYINPUT121), .B1(new_n1145), .B2(KEYINPUT61), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT121), .ZN(new_n1147));
  NOR3_X1   g722(.A1(new_n1144), .A2(new_n1147), .A3(new_n1120), .ZN(new_n1148));
  OAI211_X1 g723(.A(new_n1124), .B(new_n1143), .C1(new_n1146), .C2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1117), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1128), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1150), .B1(new_n1151), .B2(new_n1118), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1096), .A2(new_n578), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1093), .A2(G40), .A3(G160), .A4(new_n1094), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n550), .B1(new_n1092), .B2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g730(.A(KEYINPUT54), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1092), .A2(G301), .A3(new_n1154), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1157), .A2(KEYINPUT125), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT54), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT125), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1092), .A2(new_n1160), .A3(G301), .A4(new_n1154), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n1158), .A2(new_n1097), .A3(new_n1159), .A4(new_n1161), .ZN(new_n1162));
  AOI22_X1  g737(.A1(new_n1149), .A2(new_n1152), .B1(new_n1156), .B2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1096), .A2(new_n1098), .A3(new_n578), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1088), .A2(new_n1164), .ZN(new_n1165));
  OAI211_X1 g740(.A(new_n1100), .B(new_n1101), .C1(new_n1163), .C2(new_n1165), .ZN(new_n1166));
  AOI211_X1 g741(.A(new_n986), .B(new_n990), .C1(new_n1071), .C2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(new_n1043), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1169), .A2(KEYINPUT115), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1170), .A2(new_n1171), .A3(new_n1070), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1149), .A2(new_n1152), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1162), .A2(new_n1156), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1165), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1101), .B1(new_n1088), .B2(new_n1099), .ZN(new_n1176));
  OAI211_X1 g751(.A(new_n1168), .B(new_n1172), .C1(new_n1175), .C2(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(new_n990), .ZN(new_n1178));
  AOI21_X1  g753(.A(KEYINPUT126), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n985), .B1(new_n1167), .B2(new_n1179), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g755(.A1(G401), .A2(G227), .ZN(new_n1182));
  AND3_X1   g756(.A1(new_n887), .A2(G319), .A3(new_n1182), .ZN(new_n1183));
  NAND4_X1  g757(.A1(new_n1183), .A2(new_n691), .A3(new_n943), .A4(new_n945), .ZN(G225));
  INV_X1    g758(.A(G225), .ZN(G308));
endmodule


