//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1 1 1 0 0 1 1 1 1 1 0 0 0 0 0 1 1 0 1 1 1 0 1 1 1 1 0 0 1 1 0 0 1 1 0 1 1 1 0 0 1 0 1 0 0 1 1 1 1 0 1 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:40 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n565, new_n567, new_n568, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n583, new_n584, new_n586, new_n587, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n620, new_n622, new_n623, new_n624, new_n625, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n848, new_n849, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1193, new_n1194, new_n1195;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  XNOR2_X1  g016(.A(KEYINPUT64), .B(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT65), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G125), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n463), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AND2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  OAI211_X1 g044(.A(G137), .B(new_n463), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G101), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n463), .A2(G2104), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n467), .A2(new_n473), .ZN(G160));
  INV_X1    g049(.A(KEYINPUT3), .ZN(new_n475));
  INV_X1    g050(.A(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n463), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n463), .A2(G112), .ZN(new_n481));
  OR3_X1    g056(.A1(KEYINPUT67), .A2(G100), .A3(G2105), .ZN(new_n482));
  OAI21_X1  g057(.A(KEYINPUT67), .B1(G100), .B2(G2105), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n482), .A2(G2104), .A3(new_n483), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n480), .B1(new_n481), .B2(new_n484), .ZN(new_n485));
  AOI21_X1  g060(.A(G2105), .B1(new_n477), .B2(new_n478), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT66), .ZN(new_n487));
  XNOR2_X1  g062(.A(new_n486), .B(new_n487), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n485), .B1(new_n488), .B2(G136), .ZN(G162));
  OAI211_X1 g064(.A(G138), .B(new_n463), .C1(new_n468), .C2(new_n469), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT70), .ZN(new_n491));
  OAI21_X1  g066(.A(KEYINPUT69), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT69), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n486), .A2(new_n493), .A3(G138), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n492), .A2(KEYINPUT4), .A3(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  OAI211_X1 g071(.A(KEYINPUT69), .B(new_n496), .C1(new_n490), .C2(new_n491), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT68), .ZN(new_n498));
  OAI21_X1  g073(.A(G2104), .B1(new_n463), .B2(G114), .ZN(new_n499));
  NOR2_X1   g074(.A1(G102), .A2(G2105), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  OR2_X1    g076(.A1(G102), .A2(G2105), .ZN(new_n502));
  INV_X1    g077(.A(G114), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G2105), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n502), .A2(new_n504), .A3(KEYINPUT68), .A4(G2104), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n501), .A2(new_n505), .B1(new_n479), .B2(G126), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n495), .A2(new_n497), .A3(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(G164));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  OAI21_X1  g084(.A(KEYINPUT71), .B1(new_n509), .B2(KEYINPUT6), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT71), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT6), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n511), .A2(new_n512), .A3(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n509), .A2(KEYINPUT6), .ZN(new_n515));
  AND2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n516), .A2(G50), .A3(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(KEYINPUT72), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n514), .A2(new_n515), .ZN(new_n519));
  INV_X1    g094(.A(G543), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT72), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n521), .A2(new_n522), .A3(G50), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n518), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n520), .A2(KEYINPUT5), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT5), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G543), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n528), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n529), .A2(new_n509), .ZN(new_n530));
  AND3_X1   g105(.A1(new_n516), .A2(G88), .A3(new_n528), .ZN(new_n531));
  INV_X1    g106(.A(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n524), .A2(new_n530), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(KEYINPUT73), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n531), .B1(new_n518), .B2(new_n523), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT73), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n535), .A2(new_n536), .A3(new_n530), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n534), .A2(new_n537), .ZN(G166));
  NAND3_X1  g113(.A1(new_n516), .A2(G51), .A3(G543), .ZN(new_n539));
  NAND3_X1  g114(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT7), .ZN(new_n541));
  NAND4_X1  g116(.A1(new_n528), .A2(new_n514), .A3(G89), .A4(new_n515), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n528), .A2(G63), .A3(G651), .ZN(new_n543));
  NAND4_X1  g118(.A1(new_n539), .A2(new_n541), .A3(new_n542), .A4(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(G168));
  NAND2_X1  g120(.A1(G77), .A2(G543), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n525), .A2(new_n527), .ZN(new_n547));
  INV_X1    g122(.A(G64), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n521), .A2(G52), .B1(G651), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n519), .A2(new_n547), .ZN(new_n551));
  XOR2_X1   g126(.A(KEYINPUT74), .B(G90), .Z(new_n552));
  NAND2_X1  g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n550), .A2(new_n553), .ZN(G301));
  INV_X1    g129(.A(G301), .ZN(G171));
  AOI22_X1  g130(.A1(new_n528), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n556));
  OR2_X1    g131(.A1(new_n556), .A2(new_n509), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n516), .A2(G43), .A3(G543), .ZN(new_n558));
  NAND4_X1  g133(.A1(new_n528), .A2(new_n514), .A3(G81), .A4(new_n515), .ZN(new_n559));
  AND3_X1   g134(.A1(new_n558), .A2(KEYINPUT75), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g135(.A(KEYINPUT75), .B1(new_n558), .B2(new_n559), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n557), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(G153));
  AND3_X1   g139(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G36), .ZN(G176));
  NAND2_X1  g141(.A1(G1), .A2(G3), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT8), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n565), .A2(new_n568), .ZN(G188));
  NAND4_X1  g144(.A1(new_n514), .A2(G53), .A3(G543), .A4(new_n515), .ZN(new_n570));
  OR2_X1    g145(.A1(new_n570), .A2(KEYINPUT9), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(KEYINPUT9), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n571), .A2(new_n572), .B1(G91), .B2(new_n551), .ZN(new_n573));
  NAND2_X1  g148(.A1(G78), .A2(G543), .ZN(new_n574));
  XOR2_X1   g149(.A(new_n574), .B(KEYINPUT76), .Z(new_n575));
  AND3_X1   g150(.A1(new_n525), .A2(new_n527), .A3(G65), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(KEYINPUT77), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT77), .ZN(new_n579));
  OAI211_X1 g154(.A(new_n579), .B(G651), .C1(new_n575), .C2(new_n576), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n573), .A2(new_n581), .ZN(G299));
  AND2_X1   g157(.A1(new_n544), .A2(KEYINPUT78), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n544), .A2(KEYINPUT78), .ZN(new_n584));
  OR2_X1    g159(.A1(new_n583), .A2(new_n584), .ZN(G286));
  AND4_X1   g160(.A1(new_n536), .A2(new_n524), .A3(new_n530), .A4(new_n532), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n536), .B1(new_n535), .B2(new_n530), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n586), .A2(new_n587), .ZN(G303));
  NAND4_X1  g163(.A1(new_n528), .A2(new_n514), .A3(G87), .A4(new_n515), .ZN(new_n589));
  OAI21_X1  g164(.A(G651), .B1(new_n528), .B2(G74), .ZN(new_n590));
  NAND4_X1  g165(.A1(new_n514), .A2(G49), .A3(G543), .A4(new_n515), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(G288));
  NAND2_X1  g167(.A1(G73), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G61), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n547), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n595), .A2(G651), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT79), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND4_X1  g173(.A1(new_n528), .A2(new_n514), .A3(G86), .A4(new_n515), .ZN(new_n599));
  NAND4_X1  g174(.A1(new_n514), .A2(G48), .A3(G543), .A4(new_n515), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n595), .A2(KEYINPUT79), .A3(G651), .ZN(new_n601));
  NAND4_X1  g176(.A1(new_n598), .A2(new_n599), .A3(new_n600), .A4(new_n601), .ZN(G305));
  AOI22_X1  g177(.A1(new_n528), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n603));
  OR2_X1    g178(.A1(new_n603), .A2(new_n509), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n551), .A2(G85), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n521), .A2(G47), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(G290));
  NAND2_X1  g182(.A1(G301), .A2(G868), .ZN(new_n608));
  NAND4_X1  g183(.A1(new_n528), .A2(new_n514), .A3(G92), .A4(new_n515), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT10), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n609), .B(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n521), .A2(G54), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n528), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n613));
  OR2_X1    g188(.A1(new_n613), .A2(new_n509), .ZN(new_n614));
  AND3_X1   g189(.A1(new_n611), .A2(new_n612), .A3(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n608), .B1(new_n615), .B2(G868), .ZN(G321));
  XOR2_X1   g191(.A(G321), .B(KEYINPUT80), .Z(G284));
  MUX2_X1   g192(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g193(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n615), .B1(new_n620), .B2(G860), .ZN(G148));
  NAND3_X1  g196(.A1(new_n611), .A2(new_n612), .A3(new_n614), .ZN(new_n622));
  NOR2_X1   g197(.A1(new_n622), .A2(G559), .ZN(new_n623));
  INV_X1    g198(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(G868), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(G868), .B2(new_n563), .ZN(G323));
  XNOR2_X1  g201(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g202(.A1(new_n479), .A2(G123), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(KEYINPUT82), .Z(new_n629));
  INV_X1    g204(.A(G111), .ZN(new_n630));
  AND3_X1   g205(.A1(new_n630), .A2(KEYINPUT83), .A3(G2105), .ZN(new_n631));
  AOI21_X1  g206(.A(KEYINPUT83), .B1(new_n630), .B2(G2105), .ZN(new_n632));
  OAI221_X1 g207(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n631), .C2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n488), .A2(G135), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n629), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  INV_X1    g210(.A(G2096), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT81), .B(KEYINPUT12), .ZN(new_n638));
  NOR3_X1   g213(.A1(new_n475), .A2(new_n476), .A3(G2105), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT13), .B(G2100), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n637), .A2(new_n642), .ZN(G156));
  XNOR2_X1  g218(.A(G2451), .B(G2454), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT84), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT16), .ZN(new_n646));
  XNOR2_X1  g221(.A(G1341), .B(G1348), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT85), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n646), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2443), .B(G2446), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(KEYINPUT15), .B(G2430), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2435), .ZN(new_n653));
  XOR2_X1   g228(.A(G2427), .B(G2438), .Z(new_n654));
  XOR2_X1   g229(.A(new_n653), .B(new_n654), .Z(new_n655));
  NAND2_X1  g230(.A1(new_n655), .A2(KEYINPUT14), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n651), .B(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n657), .A2(G14), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(G401));
  XNOR2_X1  g234(.A(G2067), .B(G2678), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT86), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2072), .B(G2078), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2084), .B(G2090), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n661), .A2(new_n662), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT87), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT18), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n662), .B(KEYINPUT17), .ZN(new_n668));
  NOR3_X1   g243(.A1(new_n668), .A2(new_n661), .A3(new_n663), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT89), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n668), .A2(new_n661), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n663), .B1(new_n661), .B2(new_n662), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(KEYINPUT88), .Z(new_n673));
  AOI21_X1  g248(.A(new_n670), .B1(new_n671), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n667), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n675), .A2(G2100), .ZN(new_n676));
  INV_X1    g251(.A(G2100), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n667), .A2(new_n674), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n679), .A2(KEYINPUT90), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n679), .A2(KEYINPUT90), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n636), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(new_n682), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n684), .A2(G2096), .A3(new_n680), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n683), .A2(new_n685), .ZN(G227));
  XNOR2_X1  g261(.A(G1971), .B(G1976), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT19), .ZN(new_n688));
  XOR2_X1   g263(.A(G1956), .B(G2474), .Z(new_n689));
  XOR2_X1   g264(.A(G1961), .B(G1966), .Z(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(new_n688), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n689), .A2(new_n690), .ZN(new_n694));
  AOI22_X1  g269(.A1(new_n692), .A2(KEYINPUT20), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(new_n694), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n696), .A2(new_n688), .A3(new_n691), .ZN(new_n697));
  OAI211_X1 g272(.A(new_n695), .B(new_n697), .C1(KEYINPUT20), .C2(new_n692), .ZN(new_n698));
  XOR2_X1   g273(.A(G1991), .B(G1996), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1981), .B(G1986), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XOR2_X1   g277(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(G229));
  NOR2_X1   g279(.A1(G16), .A2(G22), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(G166), .B2(G16), .ZN(new_n706));
  INV_X1    g281(.A(G1971), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(G16), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G6), .ZN(new_n710));
  INV_X1    g285(.A(G305), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n710), .B1(new_n711), .B2(new_n709), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT94), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT32), .B(G1981), .Z(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  NOR2_X1   g290(.A1(G16), .A2(G23), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT95), .ZN(new_n717));
  XNOR2_X1  g292(.A(G288), .B(new_n717), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n716), .B1(new_n718), .B2(G16), .ZN(new_n719));
  XOR2_X1   g294(.A(KEYINPUT33), .B(G1976), .Z(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT96), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n719), .B(new_n721), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n708), .A2(new_n715), .A3(new_n722), .ZN(new_n723));
  XNOR2_X1  g298(.A(KEYINPUT93), .B(KEYINPUT34), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  AND2_X1   g300(.A1(KEYINPUT91), .A2(G29), .ZN(new_n726));
  NOR2_X1   g301(.A1(KEYINPUT91), .A2(G29), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(G25), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n479), .A2(G119), .ZN(new_n730));
  NOR2_X1   g305(.A1(G95), .A2(G2105), .ZN(new_n731));
  OAI21_X1  g306(.A(G2104), .B1(new_n463), .B2(G107), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n730), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(new_n488), .B2(G131), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n729), .B1(new_n734), .B2(new_n728), .ZN(new_n735));
  XNOR2_X1  g310(.A(KEYINPUT35), .B(G1991), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  AND2_X1   g312(.A1(new_n709), .A2(G24), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(G290), .B2(G16), .ZN(new_n739));
  MUX2_X1   g314(.A(new_n738), .B(new_n739), .S(KEYINPUT92), .Z(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n737), .B1(new_n741), .B2(G1986), .ZN(new_n742));
  AND2_X1   g317(.A1(new_n725), .A2(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(G1986), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n740), .A2(new_n744), .ZN(new_n745));
  OR2_X1    g320(.A1(new_n723), .A2(new_n724), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n743), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n747), .A2(KEYINPUT36), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT36), .ZN(new_n749));
  NAND4_X1  g324(.A1(new_n743), .A2(new_n749), .A3(new_n745), .A4(new_n746), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n709), .A2(G5), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G171), .B2(new_n709), .ZN(new_n752));
  INV_X1    g327(.A(G1961), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(G29), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n755), .A2(G33), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT25), .ZN(new_n758));
  AOI22_X1  g333(.A1(new_n464), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n759), .A2(new_n463), .ZN(new_n760));
  AOI211_X1 g335(.A(new_n758), .B(new_n760), .C1(G139), .C2(new_n488), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n756), .B1(new_n761), .B2(new_n755), .ZN(new_n762));
  NOR2_X1   g337(.A1(G16), .A2(G21), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(G168), .B2(G16), .ZN(new_n764));
  AOI22_X1  g339(.A1(new_n762), .A2(G2072), .B1(new_n764), .B2(G1966), .ZN(new_n765));
  OAI211_X1 g340(.A(new_n754), .B(new_n765), .C1(G2072), .C2(new_n762), .ZN(new_n766));
  NOR2_X1   g341(.A1(G164), .A2(new_n728), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(G27), .B2(new_n728), .ZN(new_n768));
  INV_X1    g343(.A(G2078), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n615), .A2(G16), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G4), .B2(G16), .ZN(new_n772));
  INV_X1    g347(.A(G1348), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n728), .A2(G35), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G162), .B2(new_n728), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT29), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n777), .A2(G2090), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n768), .A2(new_n769), .ZN(new_n779));
  NAND4_X1  g354(.A1(new_n770), .A2(new_n774), .A3(new_n778), .A4(new_n779), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT24), .B(G34), .ZN(new_n781));
  AOI22_X1  g356(.A1(G160), .A2(G29), .B1(new_n728), .B2(new_n781), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n782), .A2(G2084), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT103), .Z(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT102), .B(KEYINPUT30), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(G28), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n786), .A2(new_n755), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(new_n635), .B2(new_n728), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(G2084), .B2(new_n782), .ZN(new_n789));
  OAI211_X1 g364(.A(new_n784), .B(new_n789), .C1(new_n773), .C2(new_n772), .ZN(new_n790));
  NOR3_X1   g365(.A1(new_n766), .A2(new_n780), .A3(new_n790), .ZN(new_n791));
  XNOR2_X1  g366(.A(KEYINPUT31), .B(G11), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT23), .ZN(new_n793));
  AND2_X1   g368(.A1(new_n709), .A2(G20), .ZN(new_n794));
  AOI211_X1 g369(.A(new_n793), .B(new_n794), .C1(G299), .C2(G16), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(new_n793), .B2(new_n794), .ZN(new_n796));
  INV_X1    g371(.A(G1956), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  AND3_X1   g373(.A1(new_n791), .A2(new_n792), .A3(new_n798), .ZN(new_n799));
  NOR2_X1   g374(.A1(G29), .A2(G32), .ZN(new_n800));
  NAND3_X1  g375(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT100), .ZN(new_n802));
  INV_X1    g377(.A(KEYINPUT26), .ZN(new_n803));
  INV_X1    g378(.A(G105), .ZN(new_n804));
  OAI22_X1  g379(.A1(new_n802), .A2(new_n803), .B1(new_n804), .B2(new_n472), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(new_n803), .B2(new_n802), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n479), .A2(G129), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  AND2_X1   g383(.A1(new_n488), .A2(G141), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  AOI211_X1 g385(.A(KEYINPUT101), .B(new_n800), .C1(new_n810), .C2(G29), .ZN(new_n811));
  INV_X1    g386(.A(new_n810), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n812), .A2(new_n755), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n811), .B1(KEYINPUT101), .B2(new_n813), .ZN(new_n814));
  XOR2_X1   g389(.A(KEYINPUT27), .B(G1996), .Z(new_n815));
  INV_X1    g390(.A(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  OR2_X1    g392(.A1(new_n777), .A2(G2090), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n818), .A2(KEYINPUT104), .ZN(new_n819));
  INV_X1    g394(.A(G1341), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n563), .A2(new_n709), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n821), .B1(new_n709), .B2(G19), .ZN(new_n822));
  OAI211_X1 g397(.A(new_n817), .B(new_n819), .C1(new_n820), .C2(new_n822), .ZN(new_n823));
  OAI22_X1  g398(.A1(new_n814), .A2(new_n816), .B1(new_n818), .B2(KEYINPUT104), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n822), .A2(new_n820), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(G1966), .B2(new_n764), .ZN(new_n826));
  NOR3_X1   g401(.A1(new_n823), .A2(new_n824), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n479), .A2(G128), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT97), .Z(new_n829));
  OAI21_X1  g404(.A(KEYINPUT98), .B1(G104), .B2(G2105), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  NOR3_X1   g406(.A1(KEYINPUT98), .A2(G104), .A3(G2105), .ZN(new_n832));
  OAI221_X1 g407(.A(G2104), .B1(G116), .B2(new_n463), .C1(new_n831), .C2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n488), .A2(G140), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n829), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n835), .A2(G29), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n728), .A2(KEYINPUT28), .A3(G26), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g413(.A(KEYINPUT28), .B1(new_n728), .B2(G26), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(KEYINPUT99), .B(G2067), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n799), .A2(new_n827), .A3(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT105), .ZN(new_n844));
  OR2_X1    g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n843), .A2(new_n844), .ZN(new_n846));
  AOI22_X1  g421(.A1(new_n748), .A2(new_n750), .B1(new_n845), .B2(new_n846), .ZN(G311));
  NAND2_X1  g422(.A1(new_n748), .A2(new_n750), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n845), .A2(new_n846), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(G150));
  INV_X1    g425(.A(KEYINPUT107), .ZN(new_n851));
  OAI211_X1 g426(.A(new_n851), .B(new_n557), .C1(new_n560), .C2(new_n561), .ZN(new_n852));
  AOI22_X1  g427(.A1(new_n528), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n853));
  OR2_X1    g428(.A1(new_n853), .A2(new_n509), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n551), .A2(G93), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n521), .A2(G55), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n852), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n558), .A2(new_n559), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT75), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n558), .A2(KEYINPUT75), .A3(new_n559), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n851), .B1(new_n864), .B2(new_n557), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n859), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n562), .A2(KEYINPUT107), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n867), .A2(new_n858), .A3(new_n852), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(KEYINPUT106), .B(KEYINPUT38), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n869), .B(new_n870), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n622), .A2(new_n620), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT39), .ZN(new_n873));
  AND2_X1   g448(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n871), .A2(new_n873), .ZN(new_n875));
  NOR3_X1   g450(.A1(new_n874), .A2(new_n875), .A3(G860), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(KEYINPUT108), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n857), .A2(G860), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT109), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(KEYINPUT37), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n877), .A2(new_n880), .ZN(G145));
  XNOR2_X1  g456(.A(G162), .B(KEYINPUT110), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n810), .B(new_n640), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n835), .B(G164), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n884), .B(new_n885), .ZN(new_n886));
  XOR2_X1   g461(.A(new_n635), .B(G160), .Z(new_n887));
  NAND2_X1  g462(.A1(new_n479), .A2(G130), .ZN(new_n888));
  NOR2_X1   g463(.A1(G106), .A2(G2105), .ZN(new_n889));
  OAI21_X1  g464(.A(G2104), .B1(new_n463), .B2(G118), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n891), .B1(new_n488), .B2(G142), .ZN(new_n892));
  XOR2_X1   g467(.A(new_n734), .B(new_n892), .Z(new_n893));
  AND2_X1   g468(.A1(new_n893), .A2(new_n761), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n893), .A2(new_n761), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n887), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n894), .A2(new_n895), .ZN(new_n897));
  INV_X1    g472(.A(new_n887), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n886), .B1(new_n896), .B2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n886), .A2(new_n899), .A3(new_n896), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n883), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n902), .ZN(new_n904));
  NOR3_X1   g479(.A1(new_n904), .A2(new_n900), .A3(new_n882), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(KEYINPUT111), .B(G37), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g484(.A1(new_n857), .A2(G868), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n869), .B(new_n624), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n615), .A2(G299), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n622), .A2(new_n573), .A3(new_n581), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n912), .A2(KEYINPUT112), .A3(new_n913), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n914), .B1(KEYINPUT112), .B2(new_n912), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n911), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(KEYINPUT41), .B1(new_n912), .B2(new_n913), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n918), .B1(new_n915), .B2(KEYINPUT41), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n917), .B1(new_n911), .B2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT113), .ZN(new_n921));
  OR2_X1    g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n718), .A2(new_n711), .ZN(new_n923));
  XNOR2_X1  g498(.A(G288), .B(KEYINPUT95), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(G305), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n926), .A2(new_n537), .A3(new_n534), .ZN(new_n927));
  OAI211_X1 g502(.A(new_n925), .B(new_n923), .C1(new_n586), .C2(new_n587), .ZN(new_n928));
  INV_X1    g503(.A(G290), .ZN(new_n929));
  AND3_X1   g504(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n929), .B1(new_n927), .B2(new_n928), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  XOR2_X1   g507(.A(new_n932), .B(KEYINPUT42), .Z(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n920), .A2(new_n921), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n922), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n933), .A2(new_n921), .A3(new_n920), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n910), .B1(new_n938), .B2(G868), .ZN(G295));
  AOI21_X1  g514(.A(new_n910), .B1(new_n938), .B2(G868), .ZN(G331));
  OAI21_X1  g515(.A(G171), .B1(new_n583), .B2(new_n584), .ZN(new_n941));
  NAND2_X1  g516(.A1(G168), .A2(G301), .ZN(new_n942));
  AND2_X1   g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n859), .A2(new_n865), .ZN(new_n944));
  NOR3_X1   g519(.A1(new_n563), .A2(new_n851), .A3(new_n858), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n943), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n941), .A2(new_n942), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n866), .A2(new_n868), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(new_n919), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n946), .A2(new_n915), .A3(new_n948), .ZN(new_n951));
  AND3_X1   g526(.A1(new_n950), .A2(new_n932), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n932), .B1(new_n950), .B2(new_n951), .ZN(new_n953));
  NOR3_X1   g528(.A1(new_n952), .A2(new_n953), .A3(G37), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT43), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT114), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n912), .A2(new_n913), .ZN(new_n957));
  AND3_X1   g532(.A1(new_n866), .A2(new_n868), .A3(new_n947), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n947), .B1(new_n866), .B2(new_n868), .ZN(new_n959));
  OAI211_X1 g534(.A(KEYINPUT41), .B(new_n957), .C1(new_n958), .C2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(new_n932), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n916), .B1(new_n949), .B2(KEYINPUT41), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n907), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  OR3_X1    g538(.A1(new_n963), .A2(KEYINPUT43), .A3(new_n953), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n950), .A2(new_n951), .ZN(new_n965));
  INV_X1    g540(.A(new_n932), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(G37), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n950), .A2(new_n932), .A3(new_n951), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n967), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT114), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n970), .A2(new_n971), .A3(KEYINPUT43), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n956), .A2(new_n964), .A3(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT44), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(KEYINPUT43), .B1(new_n963), .B2(new_n953), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n967), .A2(new_n955), .A3(new_n968), .A4(new_n969), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n976), .A2(KEYINPUT44), .A3(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(KEYINPUT115), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT115), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n976), .A2(new_n977), .A3(new_n980), .A4(KEYINPUT44), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n975), .A2(new_n982), .ZN(G397));
  XOR2_X1   g558(.A(KEYINPUT116), .B(G1384), .Z(new_n984));
  AOI21_X1  g559(.A(KEYINPUT45), .B1(new_n507), .B2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(G40), .ZN(new_n986));
  NOR3_X1   g561(.A1(new_n467), .A2(new_n986), .A3(new_n473), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n810), .B(G1996), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n835), .B(G2067), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(new_n736), .ZN(new_n992));
  AND2_X1   g567(.A1(new_n734), .A2(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n989), .A2(new_n991), .A3(new_n993), .ZN(new_n994));
  OR2_X1    g569(.A1(new_n835), .A2(G2067), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n988), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(new_n988), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n997), .B1(new_n990), .B2(new_n812), .ZN(new_n998));
  INV_X1    g573(.A(G1996), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n997), .A2(KEYINPUT46), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT46), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n1001), .B1(new_n988), .B2(G1996), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n998), .A2(new_n1000), .A3(new_n1002), .ZN(new_n1003));
  XOR2_X1   g578(.A(new_n1003), .B(KEYINPUT47), .Z(new_n1004));
  NAND2_X1  g579(.A1(new_n989), .A2(new_n991), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n734), .A2(new_n992), .ZN(new_n1006));
  NOR3_X1   g581(.A1(new_n1005), .A2(new_n993), .A3(new_n1006), .ZN(new_n1007));
  OR2_X1    g582(.A1(new_n1007), .A2(new_n988), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n997), .A2(new_n744), .A3(new_n929), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n1009), .B(KEYINPUT48), .ZN(new_n1010));
  AOI211_X1 g585(.A(new_n996), .B(new_n1004), .C1(new_n1008), .C2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(new_n987), .ZN(new_n1012));
  INV_X1    g587(.A(G1384), .ZN(new_n1013));
  AND3_X1   g588(.A1(new_n492), .A2(KEYINPUT4), .A3(new_n494), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n506), .A2(new_n497), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1013), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT45), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1012), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  AND2_X1   g593(.A1(new_n506), .A2(new_n497), .ZN(new_n1019));
  AOI21_X1  g594(.A(G1384), .B1(new_n1019), .B2(new_n495), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(KEYINPUT45), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1018), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(G1966), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g599(.A(KEYINPUT117), .B(KEYINPUT50), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  OAI211_X1 g601(.A(new_n1013), .B(new_n1026), .C1(new_n1014), .C2(new_n1015), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(new_n987), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT50), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1029), .B1(new_n507), .B2(new_n1013), .ZN(new_n1030));
  OR3_X1    g605(.A1(new_n1028), .A2(G2084), .A3(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1024), .A2(new_n1031), .ZN(new_n1032));
  OAI211_X1 g607(.A(KEYINPUT51), .B(G8), .C1(new_n1032), .C2(new_n544), .ZN(new_n1033));
  AOI21_X1  g608(.A(G1966), .B1(new_n1018), .B2(new_n1021), .ZN(new_n1034));
  NOR3_X1   g609(.A1(new_n1028), .A2(G2084), .A3(new_n1030), .ZN(new_n1035));
  OAI21_X1  g610(.A(G8), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT51), .ZN(new_n1037));
  INV_X1    g612(.A(G8), .ZN(new_n1038));
  NOR2_X1   g613(.A1(G168), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1036), .A2(new_n1037), .A3(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1033), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1032), .A2(new_n1039), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(KEYINPUT62), .ZN(new_n1045));
  XNOR2_X1  g620(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1046), .B1(G166), .B2(new_n1038), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1046), .ZN(new_n1048));
  NAND3_X1  g623(.A1(G303), .A2(G8), .A3(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT119), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1026), .B1(new_n507), .B2(new_n1013), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1051), .B1(new_n1052), .B2(new_n1012), .ZN(new_n1053));
  OAI211_X1 g628(.A(KEYINPUT119), .B(new_n987), .C1(new_n1020), .C2(new_n1026), .ZN(new_n1054));
  INV_X1    g629(.A(G2090), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1020), .A2(new_n1029), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1053), .A2(new_n1054), .A3(new_n1055), .A4(new_n1056), .ZN(new_n1057));
  OAI211_X1 g632(.A(KEYINPUT45), .B(new_n984), .C1(new_n1014), .C2(new_n1015), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n987), .B(new_n1058), .C1(new_n1020), .C2(KEYINPUT45), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(new_n707), .ZN(new_n1060));
  AND2_X1   g635(.A1(new_n1057), .A2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1050), .B1(new_n1061), .B2(new_n1038), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n596), .A2(new_n599), .A3(new_n600), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(G1981), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1064), .B1(G305), .B2(G1981), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT49), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n987), .B(new_n1013), .C1(new_n1014), .C2(new_n1015), .ZN(new_n1068));
  OAI211_X1 g643(.A(KEYINPUT49), .B(new_n1064), .C1(G305), .C2(G1981), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1067), .A2(G8), .A3(new_n1068), .A4(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(G1976), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n924), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1068), .A2(G8), .ZN(new_n1073));
  OAI21_X1  g648(.A(KEYINPUT52), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n718), .A2(G1976), .ZN(new_n1075));
  AOI21_X1  g650(.A(KEYINPUT52), .B1(G288), .B2(new_n1071), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1075), .A2(G8), .A3(new_n1068), .A4(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1070), .A2(new_n1074), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT120), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1070), .A2(new_n1074), .A3(new_n1077), .A4(KEYINPUT120), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1016), .A2(KEYINPUT50), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1083), .A2(new_n1055), .A3(new_n987), .A4(new_n1027), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1038), .B1(new_n1060), .B2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1047), .A2(new_n1049), .A3(new_n1085), .ZN(new_n1086));
  AND3_X1   g661(.A1(new_n1062), .A2(new_n1082), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1059), .ZN(new_n1088));
  AOI21_X1  g663(.A(KEYINPUT53), .B1(new_n1088), .B2(new_n769), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT122), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1091), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1083), .A2(KEYINPUT122), .A3(new_n987), .A4(new_n1027), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(new_n753), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n769), .A2(KEYINPUT53), .ZN(new_n1096));
  OAI211_X1 g671(.A(new_n1090), .B(new_n1095), .C1(new_n1022), .C2(new_n1096), .ZN(new_n1097));
  AND2_X1   g672(.A1(new_n1097), .A2(G171), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT62), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1042), .A2(new_n1099), .A3(new_n1043), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1045), .A2(new_n1087), .A3(new_n1098), .A4(new_n1100), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1036), .A2(G286), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1062), .A2(new_n1082), .A3(new_n1086), .A4(new_n1102), .ZN(new_n1103));
  XNOR2_X1  g678(.A(KEYINPUT121), .B(KEYINPUT63), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1078), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1050), .ZN(new_n1107));
  OAI211_X1 g682(.A(KEYINPUT63), .B(new_n1106), .C1(new_n1107), .C2(new_n1085), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1105), .A2(new_n1108), .ZN(new_n1109));
  OR2_X1    g684(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1086), .A2(new_n1078), .ZN(new_n1111));
  INV_X1    g686(.A(G288), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1070), .A2(new_n1071), .A3(new_n1112), .ZN(new_n1113));
  OR2_X1    g688(.A1(G305), .A2(G1981), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1073), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1111), .A2(new_n1115), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1101), .A2(new_n1109), .A3(new_n1110), .A4(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1053), .A2(new_n1056), .A3(new_n1054), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(new_n797), .ZN(new_n1119));
  XNOR2_X1  g694(.A(KEYINPUT56), .B(G2072), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1088), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  AND3_X1   g697(.A1(new_n573), .A2(new_n581), .A3(KEYINPUT57), .ZN(new_n1123));
  AOI21_X1  g698(.A(KEYINPUT57), .B1(new_n573), .B2(new_n581), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1122), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1125), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1119), .A2(new_n1127), .A3(new_n1121), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1126), .A2(KEYINPUT61), .A3(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT61), .ZN(new_n1130));
  AOI221_X4 g705(.A(new_n1125), .B1(new_n1088), .B2(new_n1120), .C1(new_n1118), .C2(new_n797), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1127), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1130), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT59), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT125), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1136), .A2(new_n999), .A3(new_n987), .A4(new_n1058), .ZN(new_n1137));
  XOR2_X1   g712(.A(KEYINPUT58), .B(G1341), .Z(new_n1138));
  NAND2_X1  g713(.A1(new_n1068), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(KEYINPUT124), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT124), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1068), .A2(new_n1141), .A3(new_n1138), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1137), .A2(new_n1140), .A3(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1135), .B1(new_n1143), .B2(new_n563), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1143), .A2(new_n1135), .A3(new_n563), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1134), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  AND3_X1   g722(.A1(new_n1143), .A2(new_n1135), .A3(new_n563), .ZN(new_n1148));
  NOR3_X1   g723(.A1(new_n1148), .A2(new_n1144), .A3(KEYINPUT59), .ZN(new_n1149));
  OAI211_X1 g724(.A(new_n1129), .B(new_n1133), .C1(new_n1147), .C2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT126), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1145), .A2(new_n1134), .A3(new_n1146), .ZN(new_n1153));
  OAI21_X1  g728(.A(KEYINPUT59), .B1(new_n1148), .B2(new_n1144), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1155), .A2(KEYINPUT126), .A3(new_n1129), .A4(new_n1133), .ZN(new_n1156));
  AOI21_X1  g731(.A(G1348), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1068), .A2(G2067), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1159), .A2(KEYINPUT60), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT60), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1162), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT127), .ZN(new_n1164));
  AND3_X1   g739(.A1(new_n1163), .A2(new_n1164), .A3(new_n615), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1164), .B1(new_n1163), .B2(new_n615), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1161), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1163), .A2(new_n615), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1168), .A2(KEYINPUT127), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1163), .A2(new_n1164), .A3(new_n615), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1169), .A2(new_n1160), .A3(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1167), .A2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1152), .A2(new_n1156), .A3(new_n1172), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n1159), .A2(new_n622), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1128), .B1(new_n1174), .B2(new_n1132), .ZN(new_n1175));
  XNOR2_X1  g750(.A(new_n1175), .B(KEYINPUT123), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1173), .A2(new_n1176), .ZN(new_n1177));
  OR2_X1    g752(.A1(new_n1097), .A2(G171), .ZN(new_n1178));
  INV_X1    g753(.A(new_n1095), .ZN(new_n1179));
  INV_X1    g754(.A(new_n1058), .ZN(new_n1180));
  NOR4_X1   g755(.A1(new_n1180), .A2(new_n985), .A3(new_n1012), .A4(new_n1096), .ZN(new_n1181));
  NOR3_X1   g756(.A1(new_n1179), .A2(new_n1089), .A3(new_n1181), .ZN(new_n1182));
  OAI211_X1 g757(.A(new_n1178), .B(KEYINPUT54), .C1(G301), .C2(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT54), .ZN(new_n1184));
  NOR4_X1   g759(.A1(new_n1179), .A2(G171), .A3(new_n1089), .A4(new_n1181), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1184), .B1(new_n1098), .B2(new_n1185), .ZN(new_n1186));
  AND4_X1   g761(.A1(new_n1044), .A2(new_n1183), .A3(new_n1087), .A4(new_n1186), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1117), .B1(new_n1177), .B2(new_n1187), .ZN(new_n1188));
  XNOR2_X1  g763(.A(G290), .B(new_n744), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n988), .B1(new_n1007), .B2(new_n1189), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1011), .B1(new_n1188), .B2(new_n1190), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g766(.A1(new_n683), .A2(new_n685), .A3(new_n658), .ZN(new_n1193));
  AOI21_X1  g767(.A(new_n1193), .B1(new_n906), .B2(new_n907), .ZN(new_n1194));
  NOR2_X1   g768(.A1(G229), .A2(new_n461), .ZN(new_n1195));
  AND3_X1   g769(.A1(new_n973), .A2(new_n1194), .A3(new_n1195), .ZN(G308));
  NAND3_X1  g770(.A1(new_n973), .A2(new_n1194), .A3(new_n1195), .ZN(G225));
endmodule


