//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 1 0 1 1 0 1 1 1 1 1 1 0 0 0 0 0 0 1 0 1 0 0 1 1 0 0 0 1 0 0 0 1 1 1 1 1 1 0 0 0 0 1 0 0 0 0 1 0 0 1 0 0 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:25 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n804, new_n805, new_n806, new_n807, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n982,
    new_n984, new_n985, new_n986, new_n987, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n996, new_n997, new_n998, new_n999,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  NOR2_X1   g001(.A1(G237), .A2(G953), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G210), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n189), .B(KEYINPUT27), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT26), .B(G101), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n190), .B(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(KEYINPUT0), .A2(G128), .ZN(new_n194));
  OR2_X1    g008(.A1(KEYINPUT0), .A2(G128), .ZN(new_n195));
  INV_X1    g009(.A(G143), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n196), .A2(G146), .ZN(new_n197));
  INV_X1    g011(.A(G146), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n198), .A2(G143), .ZN(new_n199));
  OAI211_X1 g013(.A(new_n194), .B(new_n195), .C1(new_n197), .C2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(G143), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n196), .A2(G146), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT0), .A4(G128), .ZN(new_n203));
  AND2_X1   g017(.A1(new_n200), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT11), .ZN(new_n205));
  INV_X1    g019(.A(G134), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n205), .B1(new_n206), .B2(G137), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(G137), .ZN(new_n208));
  INV_X1    g022(.A(G137), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n209), .A2(KEYINPUT11), .A3(G134), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n207), .A2(new_n208), .A3(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G131), .ZN(new_n212));
  INV_X1    g026(.A(G131), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n207), .A2(new_n210), .A3(new_n213), .A4(new_n208), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n204), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(KEYINPUT2), .B(G113), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  XNOR2_X1  g032(.A(G116), .B(G119), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n219), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(new_n217), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(G128), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n225), .A2(KEYINPUT1), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n226), .A2(new_n201), .A3(new_n202), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(G128), .B1(new_n201), .B2(new_n202), .ZN(new_n229));
  AND3_X1   g043(.A1(new_n196), .A2(KEYINPUT1), .A3(G146), .ZN(new_n230));
  OAI21_X1  g044(.A(KEYINPUT64), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n199), .A2(KEYINPUT1), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT64), .ZN(new_n233));
  XNOR2_X1  g047(.A(G143), .B(G146), .ZN(new_n234));
  OAI211_X1 g048(.A(new_n232), .B(new_n233), .C1(new_n234), .C2(G128), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n228), .B1(new_n231), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n208), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n206), .A2(G137), .ZN(new_n238));
  OAI21_X1  g052(.A(G131), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(new_n214), .ZN(new_n240));
  OAI211_X1 g054(.A(new_n216), .B(new_n224), .C1(new_n236), .C2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n242), .A2(KEYINPUT28), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n225), .B1(new_n197), .B2(new_n199), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n233), .B1(new_n244), .B2(new_n232), .ZN(new_n245));
  NOR3_X1   g059(.A1(new_n229), .A2(KEYINPUT64), .A3(new_n230), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n227), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n240), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n249), .A2(KEYINPUT65), .A3(new_n224), .A4(new_n216), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT65), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n241), .A2(new_n251), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n216), .B1(new_n236), .B2(new_n240), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(new_n223), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n250), .A2(new_n252), .A3(new_n254), .ZN(new_n255));
  AOI211_X1 g069(.A(new_n193), .B(new_n243), .C1(new_n255), .C2(KEYINPUT28), .ZN(new_n256));
  AOI21_X1  g070(.A(G902), .B1(new_n256), .B2(KEYINPUT29), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n243), .B1(new_n255), .B2(KEYINPUT28), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(new_n192), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT29), .ZN(new_n260));
  AND2_X1   g074(.A1(new_n250), .A2(new_n252), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT30), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n262), .B1(new_n249), .B2(new_n216), .ZN(new_n263));
  OAI211_X1 g077(.A(new_n216), .B(new_n262), .C1(new_n236), .C2(new_n240), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n223), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n261), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(new_n193), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n259), .A2(new_n260), .A3(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n187), .B1(new_n257), .B2(new_n269), .ZN(new_n270));
  NOR2_X1   g084(.A1(G472), .A2(G902), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n253), .A2(KEYINPUT30), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n224), .B1(new_n272), .B2(new_n264), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n250), .A2(new_n252), .ZN(new_n274));
  NOR3_X1   g088(.A1(new_n273), .A2(new_n274), .A3(new_n193), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT31), .ZN(new_n276));
  OAI22_X1  g090(.A1(new_n275), .A2(new_n276), .B1(new_n258), .B2(new_n192), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n261), .A2(new_n266), .A3(new_n276), .A4(new_n192), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n271), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(KEYINPUT32), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT32), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n282), .B(new_n271), .C1(new_n277), .C2(new_n279), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n270), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G234), .ZN(new_n285));
  OAI21_X1  g099(.A(G217), .B1(new_n285), .B2(G902), .ZN(new_n286));
  XNOR2_X1  g100(.A(new_n286), .B(KEYINPUT66), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT25), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT16), .ZN(new_n289));
  INV_X1    g103(.A(G140), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n289), .A2(new_n290), .A3(G125), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(G125), .ZN(new_n292));
  INV_X1    g106(.A(G125), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(G140), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  OAI211_X1 g109(.A(G146), .B(new_n291), .C1(new_n295), .C2(new_n289), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(KEYINPUT70), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n291), .B1(new_n295), .B2(new_n289), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(new_n198), .ZN(new_n299));
  XNOR2_X1  g113(.A(G125), .B(G140), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(KEYINPUT16), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT70), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n301), .A2(new_n302), .A3(G146), .A4(new_n291), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n297), .A2(new_n299), .A3(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G119), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(G128), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n306), .B(KEYINPUT67), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n225), .A2(G119), .ZN(new_n308));
  XOR2_X1   g122(.A(KEYINPUT24), .B(G110), .Z(new_n309));
  NAND3_X1  g123(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  AND3_X1   g124(.A1(new_n306), .A2(KEYINPUT68), .A3(KEYINPUT23), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT69), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n308), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT23), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n308), .A2(new_n312), .ZN(new_n315));
  AOI21_X1  g129(.A(KEYINPUT68), .B1(new_n305), .B2(G128), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n314), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n313), .A2(G110), .A3(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n304), .A2(new_n310), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n300), .A2(new_n198), .ZN(new_n320));
  AND2_X1   g134(.A1(new_n296), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(G110), .B1(new_n313), .B2(new_n317), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n309), .B1(new_n307), .B2(new_n308), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n321), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n319), .A2(new_n324), .ZN(new_n325));
  XNOR2_X1  g139(.A(KEYINPUT22), .B(G137), .ZN(new_n326));
  INV_X1    g140(.A(G953), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n327), .A2(G221), .A3(G234), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n326), .B(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n325), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT71), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n325), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n319), .A2(new_n324), .A3(KEYINPUT71), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n329), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n331), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n288), .B1(new_n337), .B2(G902), .ZN(new_n338));
  INV_X1    g152(.A(new_n334), .ZN(new_n339));
  AOI21_X1  g153(.A(KEYINPUT71), .B1(new_n319), .B2(new_n324), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n336), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(new_n330), .ZN(new_n342));
  INV_X1    g156(.A(G902), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n342), .A2(KEYINPUT25), .A3(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n287), .B1(new_n338), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n286), .A2(new_n343), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n337), .A2(new_n346), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n284), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(G478), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n351), .A2(KEYINPUT15), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT82), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n353), .B1(new_n225), .B2(G143), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n196), .A2(KEYINPUT82), .A3(G128), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n225), .A2(G143), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(KEYINPUT83), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT83), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n356), .A2(new_n360), .A3(new_n357), .ZN(new_n361));
  AOI21_X1  g175(.A(G134), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT13), .ZN(new_n363));
  AOI22_X1  g177(.A1(new_n356), .A2(new_n363), .B1(new_n225), .B2(G143), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n354), .A2(KEYINPUT13), .A3(new_n355), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n206), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(G107), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(KEYINPUT73), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT73), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(G107), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(G122), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(G116), .ZN(new_n373));
  INV_X1    g187(.A(G116), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(G122), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  XOR2_X1   g190(.A(new_n371), .B(new_n376), .Z(new_n377));
  NOR3_X1   g191(.A1(new_n362), .A2(new_n366), .A3(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  AND3_X1   g193(.A1(new_n356), .A2(new_n360), .A3(new_n357), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n360), .B1(new_n356), .B2(new_n357), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n206), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n359), .A2(G134), .A3(new_n361), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n371), .A2(new_n376), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n374), .A2(KEYINPUT14), .A3(G122), .ZN(new_n386));
  OAI211_X1 g200(.A(G107), .B(new_n386), .C1(new_n376), .C2(KEYINPUT14), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT84), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  AND2_X1   g203(.A1(new_n386), .A2(G107), .ZN(new_n390));
  OAI211_X1 g204(.A(new_n390), .B(KEYINPUT84), .C1(KEYINPUT14), .C2(new_n376), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n385), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  AND3_X1   g206(.A1(new_n384), .A2(KEYINPUT85), .A3(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(KEYINPUT85), .B1(new_n384), .B2(new_n392), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n379), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  XNOR2_X1  g209(.A(KEYINPUT9), .B(G234), .ZN(new_n396));
  INV_X1    g210(.A(G217), .ZN(new_n397));
  NOR3_X1   g211(.A1(new_n396), .A2(new_n397), .A3(G953), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n395), .A2(new_n399), .ZN(new_n400));
  NOR3_X1   g214(.A1(new_n380), .A2(new_n381), .A3(new_n206), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n392), .B1(new_n401), .B2(new_n362), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT85), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n384), .A2(KEYINPUT85), .A3(new_n392), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n406), .A2(new_n379), .A3(new_n398), .ZN(new_n407));
  AOI21_X1  g221(.A(G902), .B1(new_n400), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT86), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AOI211_X1 g224(.A(KEYINPUT86), .B(G902), .C1(new_n400), .C2(new_n407), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n352), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n398), .B1(new_n406), .B2(new_n379), .ZN(new_n413));
  AOI211_X1 g227(.A(new_n378), .B(new_n399), .C1(new_n404), .C2(new_n405), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n343), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(KEYINPUT86), .ZN(new_n416));
  INV_X1    g230(.A(new_n352), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(G952), .ZN(new_n419));
  AOI211_X1 g233(.A(G953), .B(new_n419), .C1(G234), .C2(G237), .ZN(new_n420));
  AOI211_X1 g234(.A(new_n343), .B(new_n327), .C1(G234), .C2(G237), .ZN(new_n421));
  XNOR2_X1  g235(.A(KEYINPUT21), .B(G898), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n420), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n412), .A2(new_n418), .A3(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(G475), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT78), .ZN(new_n427));
  INV_X1    g241(.A(G237), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n428), .A2(new_n327), .A3(G214), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT77), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n430), .A2(G143), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n188), .B(G214), .C1(new_n430), .C2(G143), .ZN(new_n433));
  AND2_X1   g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n427), .B1(new_n434), .B2(new_n213), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n432), .A2(new_n433), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n436), .A2(KEYINPUT78), .A3(G131), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n304), .B1(new_n438), .B2(KEYINPUT17), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT17), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n434), .A2(new_n213), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n435), .A2(new_n440), .A3(new_n437), .A4(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(KEYINPUT80), .ZN(new_n443));
  AOI21_X1  g257(.A(KEYINPUT78), .B1(new_n436), .B2(G131), .ZN(new_n444));
  AOI211_X1 g258(.A(new_n427), .B(new_n213), .C1(new_n432), .C2(new_n433), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT80), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n446), .A2(new_n447), .A3(new_n440), .A4(new_n441), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n439), .A2(new_n443), .A3(new_n448), .ZN(new_n449));
  XNOR2_X1  g263(.A(G113), .B(G122), .ZN(new_n450));
  INV_X1    g264(.A(G104), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n450), .B(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT18), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n434), .B1(new_n453), .B2(new_n213), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n436), .A2(KEYINPUT18), .A3(G131), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n295), .A2(G146), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(new_n320), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n454), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  AND3_X1   g272(.A1(new_n449), .A2(new_n452), .A3(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n452), .B1(new_n449), .B2(new_n458), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n343), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n426), .B1(new_n461), .B2(KEYINPUT81), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT81), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n463), .B(new_n343), .C1(new_n459), .C2(new_n460), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n449), .A2(new_n452), .A3(new_n458), .ZN(new_n466));
  AND2_X1   g280(.A1(new_n446), .A2(new_n441), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT79), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n295), .B(KEYINPUT19), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n468), .B1(new_n469), .B2(G146), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n300), .B(KEYINPUT19), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n471), .A2(KEYINPUT79), .A3(new_n198), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n470), .A2(new_n296), .A3(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n458), .B1(new_n467), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n452), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n466), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g291(.A1(G475), .A2(G902), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(KEYINPUT20), .ZN(new_n480));
  INV_X1    g294(.A(new_n478), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n481), .B1(new_n466), .B2(new_n476), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT20), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n480), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n465), .A2(new_n485), .ZN(new_n486));
  OAI21_X1  g300(.A(G210), .B1(G237), .B2(G902), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(G104), .B1(new_n368), .B2(new_n370), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT74), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n490), .B1(new_n451), .B2(G107), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n367), .A2(KEYINPUT74), .A3(G104), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(G101), .B1(new_n489), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n219), .A2(KEYINPUT5), .ZN(new_n495));
  NOR3_X1   g309(.A1(new_n374), .A2(KEYINPUT5), .A3(G119), .ZN(new_n496));
  INV_X1    g310(.A(G113), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n495), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT3), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n500), .B1(new_n367), .B2(G104), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n367), .A2(G104), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n451), .A2(KEYINPUT3), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n504), .A2(new_n368), .A3(new_n370), .ZN(new_n505));
  INV_X1    g319(.A(G101), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n503), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n494), .A2(new_n499), .A3(new_n507), .A4(new_n220), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(KEYINPUT4), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n506), .B1(new_n503), .B2(new_n505), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n503), .A2(new_n505), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT4), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n512), .A2(new_n513), .A3(G101), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n223), .A2(new_n514), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n508), .B1(new_n511), .B2(new_n515), .ZN(new_n516));
  XNOR2_X1  g330(.A(G110), .B(G122), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  OAI211_X1 g333(.A(new_n517), .B(new_n508), .C1(new_n511), .C2(new_n515), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n519), .A2(KEYINPUT6), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n236), .A2(new_n293), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n200), .A2(new_n203), .ZN(new_n523));
  AOI21_X1  g337(.A(KEYINPUT75), .B1(new_n523), .B2(G125), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n523), .A2(KEYINPUT75), .A3(G125), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n522), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(G224), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n528), .A2(G953), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  AND3_X1   g344(.A1(new_n523), .A2(KEYINPUT75), .A3(G125), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n531), .A2(new_n524), .ZN(new_n532));
  INV_X1    g346(.A(new_n529), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n532), .A2(new_n533), .A3(new_n522), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n530), .A2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT6), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n516), .A2(new_n536), .A3(new_n518), .ZN(new_n537));
  AND3_X1   g351(.A1(new_n521), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT7), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n527), .B1(new_n539), .B2(new_n529), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n532), .A2(KEYINPUT7), .A3(new_n533), .A4(new_n522), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n494), .A2(new_n507), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n499), .A2(new_n220), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT76), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n517), .B(KEYINPUT8), .ZN(new_n546));
  AND2_X1   g360(.A1(new_n542), .A2(new_n543), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n508), .A2(KEYINPUT76), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n545), .B(new_n546), .C1(new_n547), .C2(new_n548), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n540), .A2(new_n520), .A3(new_n541), .A4(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(new_n343), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n488), .B1(new_n538), .B2(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n521), .A2(new_n535), .A3(new_n537), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n553), .A2(new_n343), .A3(new_n487), .A4(new_n550), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(G469), .ZN(new_n556));
  AND3_X1   g370(.A1(new_n494), .A2(KEYINPUT10), .A3(new_n507), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n247), .A2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n215), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n244), .A2(new_n227), .A3(new_n232), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n494), .A2(new_n560), .A3(new_n507), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT10), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n204), .B(new_n514), .C1(new_n509), .C2(new_n510), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n558), .A2(new_n559), .A3(new_n563), .A4(new_n564), .ZN(new_n565));
  XNOR2_X1  g379(.A(G110), .B(G140), .ZN(new_n566));
  INV_X1    g380(.A(G227), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n567), .A2(G953), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n566), .B(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n565), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n236), .A2(new_n542), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(new_n561), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n573), .A2(KEYINPUT12), .A3(new_n215), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n215), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT12), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n571), .B1(new_n574), .B2(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n523), .B1(new_n513), .B2(new_n510), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n512), .A2(G101), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n580), .A2(KEYINPUT4), .A3(new_n507), .ZN(new_n581));
  AOI22_X1  g395(.A1(new_n579), .A2(new_n581), .B1(new_n561), .B2(new_n562), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(new_n558), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(new_n215), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n570), .B1(new_n584), .B2(new_n565), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n556), .B(new_n343), .C1(new_n578), .C2(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n584), .A2(new_n570), .A3(new_n565), .ZN(new_n587));
  INV_X1    g401(.A(new_n565), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n588), .B1(new_n577), .B2(new_n574), .ZN(new_n589));
  OAI211_X1 g403(.A(new_n587), .B(G469), .C1(new_n589), .C2(new_n570), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n556), .A2(new_n343), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n586), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  OAI21_X1  g407(.A(G214), .B1(G237), .B2(G902), .ZN(new_n594));
  OAI21_X1  g408(.A(G221), .B1(new_n396), .B2(G902), .ZN(new_n595));
  XOR2_X1   g409(.A(new_n595), .B(KEYINPUT72), .Z(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n555), .A2(new_n593), .A3(new_n594), .A4(new_n597), .ZN(new_n598));
  NOR3_X1   g412(.A1(new_n425), .A2(new_n486), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n350), .A2(new_n599), .ZN(new_n600));
  XOR2_X1   g414(.A(KEYINPUT87), .B(G101), .Z(new_n601));
  XNOR2_X1  g415(.A(new_n600), .B(new_n601), .ZN(G3));
  INV_X1    g416(.A(new_n594), .ZN(new_n603));
  AND2_X1   g417(.A1(new_n550), .A2(new_n343), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n487), .B1(new_n604), .B2(new_n553), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT88), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n603), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n552), .A2(KEYINPUT88), .A3(new_n554), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  AOI22_X1  g423(.A1(new_n462), .A2(new_n464), .B1(new_n480), .B2(new_n484), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n351), .A2(new_n343), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n611), .B1(new_n408), .B2(new_n351), .ZN(new_n612));
  OAI21_X1  g426(.A(KEYINPUT33), .B1(new_n413), .B2(new_n414), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT33), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n400), .A2(new_n407), .A3(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n613), .A2(G478), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  NOR4_X1   g431(.A1(new_n609), .A2(new_n610), .A3(new_n423), .A4(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n261), .A2(new_n266), .A3(new_n192), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(KEYINPUT31), .ZN(new_n620));
  OAI211_X1 g434(.A(new_n620), .B(new_n278), .C1(new_n192), .C2(new_n258), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(new_n343), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(G472), .ZN(new_n623));
  AOI21_X1  g437(.A(KEYINPUT12), .B1(new_n573), .B2(new_n215), .ZN(new_n624));
  AOI211_X1 g438(.A(new_n576), .B(new_n559), .C1(new_n572), .C2(new_n561), .ZN(new_n625));
  OAI211_X1 g439(.A(new_n570), .B(new_n565), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n559), .B1(new_n582), .B2(new_n558), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n569), .B1(new_n588), .B2(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(G902), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n591), .B1(new_n629), .B2(new_n556), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n596), .B1(new_n630), .B2(new_n590), .ZN(new_n631));
  AND4_X1   g445(.A1(new_n280), .A2(new_n348), .A3(new_n623), .A4(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n618), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(KEYINPUT89), .ZN(new_n634));
  XNOR2_X1  g448(.A(KEYINPUT34), .B(G104), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G6));
  NAND2_X1  g450(.A1(new_n408), .A2(new_n409), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n417), .B1(new_n416), .B2(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n410), .A2(new_n352), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n465), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT90), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n641), .B1(new_n479), .B2(KEYINPUT20), .ZN(new_n642));
  NOR3_X1   g456(.A1(new_n482), .A2(KEYINPUT90), .A3(new_n483), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT92), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n484), .A2(KEYINPUT91), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT91), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n482), .A2(new_n647), .A3(new_n483), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n644), .A2(new_n645), .A3(new_n649), .ZN(new_n650));
  OAI21_X1  g464(.A(KEYINPUT90), .B1(new_n482), .B2(new_n483), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n479), .A2(new_n641), .A3(KEYINPUT20), .ZN(new_n652));
  AND3_X1   g466(.A1(new_n482), .A2(new_n647), .A3(new_n483), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n647), .B1(new_n482), .B2(new_n483), .ZN(new_n654));
  OAI211_X1 g468(.A(new_n651), .B(new_n652), .C1(new_n653), .C2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(KEYINPUT92), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n640), .B1(new_n650), .B2(new_n656), .ZN(new_n657));
  AND3_X1   g471(.A1(new_n607), .A2(new_n424), .A3(new_n608), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n657), .A2(new_n632), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(KEYINPUT93), .ZN(new_n660));
  XNOR2_X1  g474(.A(KEYINPUT35), .B(G107), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G9));
  INV_X1    g476(.A(KEYINPUT95), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n623), .A2(new_n280), .ZN(new_n664));
  INV_X1    g478(.A(new_n346), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n336), .A2(KEYINPUT36), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(KEYINPUT94), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n335), .B(new_n667), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n345), .B1(new_n665), .B2(new_n668), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n663), .B1(new_n664), .B2(new_n669), .ZN(new_n670));
  AOI22_X1  g484(.A1(new_n622), .A2(G472), .B1(new_n271), .B2(new_n621), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n338), .A2(new_n344), .ZN(new_n672));
  INV_X1    g486(.A(new_n287), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n668), .A2(new_n665), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n671), .A2(KEYINPUT95), .A3(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n670), .A2(new_n599), .A3(new_n677), .ZN(new_n678));
  XOR2_X1   g492(.A(KEYINPUT37), .B(G110), .Z(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(KEYINPUT96), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n678), .B(new_n680), .ZN(G12));
  NAND2_X1  g495(.A1(new_n656), .A2(new_n650), .ZN(new_n682));
  AOI22_X1  g496(.A1(new_n412), .A2(new_n418), .B1(new_n464), .B2(new_n462), .ZN(new_n683));
  INV_X1    g497(.A(G900), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n420), .B1(new_n421), .B2(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n682), .A2(new_n683), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n257), .A2(new_n269), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(G472), .ZN(new_n689));
  INV_X1    g503(.A(new_n283), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n282), .B1(new_n621), .B2(new_n271), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n689), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n609), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n692), .A2(new_n631), .A3(new_n693), .A4(new_n676), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n687), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(new_n225), .ZN(G30));
  XOR2_X1   g510(.A(new_n555), .B(KEYINPUT38), .Z(new_n697));
  NOR3_X1   g511(.A1(new_n697), .A2(new_n603), .A3(new_n676), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n412), .A2(new_n418), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(new_n486), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT40), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n593), .A2(new_n597), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n685), .B(KEYINPUT39), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n700), .B1(new_n701), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n281), .A2(new_n283), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n193), .B1(new_n261), .B2(new_n266), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n343), .B1(new_n255), .B2(new_n192), .ZN(new_n708));
  OAI21_X1  g522(.A(G472), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  OAI21_X1  g524(.A(KEYINPUT40), .B1(new_n702), .B2(new_n703), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n698), .A2(new_n705), .A3(new_n710), .A4(new_n711), .ZN(new_n712));
  XOR2_X1   g526(.A(KEYINPUT97), .B(G143), .Z(new_n713));
  XNOR2_X1  g527(.A(new_n712), .B(new_n713), .ZN(G45));
  NOR3_X1   g528(.A1(new_n284), .A2(new_n702), .A3(new_n669), .ZN(new_n715));
  INV_X1    g529(.A(new_n617), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n486), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n717), .A2(new_n685), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n715), .A2(KEYINPUT98), .A3(new_n693), .A4(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT98), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n610), .A2(new_n617), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(new_n686), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n720), .B1(new_n694), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n719), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G146), .ZN(G48));
  NOR2_X1   g539(.A1(new_n629), .A2(new_n556), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n727), .A2(new_n597), .A3(new_n586), .ZN(new_n728));
  INV_X1    g542(.A(new_n728), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n350), .A2(new_n618), .A3(KEYINPUT99), .A4(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT99), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n692), .A2(new_n348), .A3(new_n729), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n658), .A2(new_n721), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n731), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n730), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(KEYINPUT41), .B(G113), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n735), .B(new_n736), .ZN(G15));
  NOR3_X1   g551(.A1(new_n284), .A2(new_n349), .A3(new_n728), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT100), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n738), .A2(new_n739), .A3(new_n658), .A4(new_n657), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n655), .A2(KEYINPUT92), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n645), .B1(new_n644), .B2(new_n649), .ZN(new_n742));
  OAI211_X1 g556(.A(new_n658), .B(new_n683), .C1(new_n741), .C2(new_n742), .ZN(new_n743));
  OAI21_X1  g557(.A(KEYINPUT100), .B1(new_n743), .B2(new_n732), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n740), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G116), .ZN(G18));
  NOR4_X1   g560(.A1(new_n425), .A2(new_n609), .A3(new_n486), .A4(new_n728), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n284), .A2(new_n669), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G119), .ZN(G21));
  NOR2_X1   g564(.A1(new_n728), .A2(new_n423), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n751), .A2(new_n693), .A3(new_n486), .A4(new_n699), .ZN(new_n752));
  INV_X1    g566(.A(new_n347), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n674), .A2(KEYINPUT102), .A3(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT102), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n755), .B1(new_n345), .B2(new_n347), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n277), .A2(KEYINPUT101), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT101), .ZN(new_n759));
  OAI211_X1 g573(.A(new_n620), .B(new_n759), .C1(new_n192), .C2(new_n258), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n758), .A2(new_n278), .A3(new_n760), .ZN(new_n761));
  AOI22_X1  g575(.A1(new_n761), .A2(new_n271), .B1(new_n622), .B2(G472), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n757), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n752), .A2(new_n763), .ZN(new_n764));
  XOR2_X1   g578(.A(KEYINPUT103), .B(G122), .Z(new_n765));
  XNOR2_X1  g579(.A(new_n764), .B(new_n765), .ZN(G24));
  NAND2_X1  g580(.A1(new_n761), .A2(new_n271), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n767), .A2(new_n676), .A3(new_n623), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT104), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n762), .A2(KEYINPUT104), .A3(new_n676), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n722), .A2(new_n609), .A3(new_n728), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(new_n293), .ZN(G27));
  AOI22_X1  g589(.A1(new_n706), .A2(new_n689), .B1(new_n754), .B2(new_n756), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n552), .A2(new_n594), .A3(new_n554), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT105), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n778), .B1(new_n631), .B2(new_n779), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n702), .A2(KEYINPUT105), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n780), .A2(new_n781), .A3(KEYINPUT106), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT106), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n777), .B1(new_n702), .B2(KEYINPUT105), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n631), .A2(new_n779), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n783), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  OAI211_X1 g600(.A(new_n776), .B(new_n718), .C1(new_n782), .C2(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n692), .A2(new_n348), .ZN(new_n788));
  OAI21_X1  g602(.A(KEYINPUT106), .B1(new_n780), .B2(new_n781), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n784), .A2(new_n783), .A3(new_n785), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n788), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n717), .A2(KEYINPUT42), .A3(new_n685), .ZN(new_n792));
  AOI22_X1  g606(.A1(new_n787), .A2(KEYINPUT42), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(KEYINPUT107), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT107), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT42), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n722), .B1(new_n789), .B2(new_n790), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n796), .B1(new_n797), .B2(new_n776), .ZN(new_n798));
  OAI211_X1 g612(.A(new_n792), .B(new_n350), .C1(new_n782), .C2(new_n786), .ZN(new_n799));
  INV_X1    g613(.A(new_n799), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n795), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n794), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(G131), .ZN(G33));
  INV_X1    g617(.A(KEYINPUT108), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n687), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n657), .A2(KEYINPUT108), .A3(new_n686), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n791), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(G134), .ZN(G36));
  NOR2_X1   g622(.A1(new_n589), .A2(new_n570), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n571), .A2(new_n627), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n811), .A2(KEYINPUT45), .ZN(new_n812));
  OAI21_X1  g626(.A(G469), .B1(new_n811), .B2(KEYINPUT45), .ZN(new_n813));
  OR2_X1    g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(new_n814), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n815), .A2(new_n591), .ZN(new_n816));
  OR2_X1    g630(.A1(new_n816), .A2(KEYINPUT46), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(KEYINPUT109), .ZN(new_n818));
  INV_X1    g632(.A(new_n586), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n819), .B1(new_n816), .B2(KEYINPUT46), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n817), .A2(KEYINPUT109), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n597), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n823), .A2(new_n703), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n486), .A2(new_n617), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n825), .B(KEYINPUT43), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n826), .A2(new_n664), .A3(new_n676), .ZN(new_n827));
  INV_X1    g641(.A(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n777), .B1(new_n828), .B2(KEYINPUT44), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n824), .B(new_n829), .C1(KEYINPUT44), .C2(new_n828), .ZN(new_n830));
  XNOR2_X1  g644(.A(KEYINPUT110), .B(G137), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n830), .B(new_n831), .ZN(G39));
  INV_X1    g646(.A(KEYINPUT47), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n833), .A2(KEYINPUT111), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n833), .A2(KEYINPUT111), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n823), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  OR2_X1    g650(.A1(new_n823), .A2(new_n835), .ZN(new_n837));
  NOR4_X1   g651(.A1(new_n722), .A2(new_n692), .A3(new_n348), .A4(new_n777), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n839), .B(G140), .ZN(G42));
  INV_X1    g654(.A(KEYINPUT116), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT115), .ZN(new_n842));
  INV_X1    g656(.A(new_n752), .ZN(new_n843));
  INV_X1    g657(.A(new_n763), .ZN(new_n844));
  AOI22_X1  g658(.A1(new_n843), .A2(new_n844), .B1(new_n747), .B2(new_n748), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n745), .A2(new_n735), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n787), .A2(KEYINPUT42), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(new_n799), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n842), .B1(new_n846), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n692), .A2(new_n676), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n609), .A2(new_n728), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n638), .A2(new_n639), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n851), .A2(new_n610), .A3(new_n852), .A4(new_n424), .ZN(new_n853));
  OAI22_X1  g667(.A1(new_n850), .A2(new_n853), .B1(new_n752), .B2(new_n763), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n854), .B1(new_n734), .B2(new_n730), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n855), .A2(new_n793), .A3(KEYINPUT115), .A4(new_n745), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n849), .A2(new_n856), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n682), .A2(new_n683), .A3(new_n686), .ZN(new_n858));
  NOR4_X1   g672(.A1(new_n284), .A2(new_n669), .A3(new_n702), .A4(new_n609), .ZN(new_n859));
  AOI22_X1  g673(.A1(new_n772), .A2(new_n773), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n700), .A2(new_n609), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n676), .A2(new_n702), .A3(new_n685), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n861), .A2(new_n710), .A3(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n860), .A2(new_n724), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(KEYINPUT52), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n702), .A2(new_n345), .A3(new_n347), .ZN(new_n866));
  AOI211_X1 g680(.A(new_n423), .B(new_n603), .C1(new_n552), .C2(new_n554), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n866), .A2(new_n721), .A3(new_n671), .A4(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(new_n598), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n869), .A2(new_n852), .A3(new_n610), .A4(new_n424), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n868), .B1(new_n788), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(KEYINPUT112), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT112), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n600), .A2(new_n873), .A3(new_n868), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  OAI211_X1 g689(.A(new_n485), .B(new_n465), .C1(new_n638), .C2(new_n639), .ZN(new_n876));
  INV_X1    g690(.A(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n632), .A2(new_n867), .A3(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n678), .A2(new_n878), .A3(KEYINPUT113), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n678), .A2(new_n878), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT113), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n875), .A2(new_n879), .A3(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT52), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n860), .A2(new_n724), .A3(new_n884), .A4(new_n863), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n699), .A2(new_n685), .A3(new_n777), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n715), .A2(new_n465), .A3(new_n682), .A4(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n797), .A2(new_n772), .ZN(new_n888));
  AND4_X1   g702(.A1(KEYINPUT53), .A2(new_n807), .A3(new_n887), .A4(new_n888), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n865), .A2(new_n883), .A3(new_n885), .A4(new_n889), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n841), .B1(new_n857), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n865), .A2(new_n885), .ZN(new_n892));
  INV_X1    g706(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n849), .A2(new_n856), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n875), .A2(new_n882), .A3(new_n879), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT53), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n807), .A2(new_n887), .A3(new_n888), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n893), .A2(new_n894), .A3(KEYINPUT116), .A4(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n891), .A2(new_n899), .ZN(new_n900));
  AND3_X1   g714(.A1(new_n807), .A2(new_n887), .A3(new_n888), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n901), .A2(new_n794), .A3(new_n801), .ZN(new_n902));
  AOI22_X1  g716(.A1(new_n872), .A2(new_n874), .B1(new_n880), .B2(new_n881), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n903), .A2(new_n745), .A3(new_n855), .A4(new_n879), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n892), .A2(new_n902), .A3(new_n904), .ZN(new_n905));
  OAI21_X1  g719(.A(KEYINPUT114), .B1(new_n905), .B2(KEYINPUT53), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT114), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n895), .A2(new_n846), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n802), .A2(new_n908), .A3(new_n901), .ZN(new_n909));
  OAI211_X1 g723(.A(new_n907), .B(new_n896), .C1(new_n909), .C2(new_n892), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n900), .A2(new_n906), .A3(new_n910), .ZN(new_n911));
  OR2_X1    g725(.A1(new_n911), .A2(KEYINPUT54), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n905), .B(KEYINPUT53), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(KEYINPUT54), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n729), .A2(new_n420), .A3(new_n778), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n826), .A2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  XNOR2_X1  g732(.A(KEYINPUT118), .B(KEYINPUT48), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n918), .A2(new_n776), .A3(new_n919), .ZN(new_n920));
  AND4_X1   g734(.A1(new_n706), .A2(new_n916), .A3(new_n348), .A4(new_n709), .ZN(new_n921));
  AOI211_X1 g735(.A(new_n419), .B(G953), .C1(new_n921), .C2(new_n721), .ZN(new_n922));
  AND3_X1   g736(.A1(new_n826), .A2(new_n420), .A3(new_n844), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(new_n851), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT48), .ZN(new_n925));
  INV_X1    g739(.A(new_n776), .ZN(new_n926));
  OAI211_X1 g740(.A(KEYINPUT118), .B(new_n925), .C1(new_n917), .C2(new_n926), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n920), .A2(new_n922), .A3(new_n924), .A4(new_n927), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n923), .A2(new_n603), .A3(new_n697), .A4(new_n729), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n929), .B(KEYINPUT50), .Z(new_n930));
  NOR2_X1   g744(.A1(new_n486), .A2(new_n716), .ZN(new_n931));
  AOI22_X1  g745(.A1(new_n918), .A2(new_n772), .B1(new_n921), .B2(new_n931), .ZN(new_n932));
  AND2_X1   g746(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n819), .A2(new_n726), .ZN(new_n934));
  AOI22_X1  g748(.A1(new_n837), .A2(new_n836), .B1(new_n596), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n923), .A2(new_n778), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n933), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT51), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n928), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  OAI221_X1 g753(.A(KEYINPUT51), .B1(new_n935), .B2(new_n936), .C1(new_n933), .C2(KEYINPUT117), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n933), .A2(KEYINPUT117), .ZN(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n939), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  OAI22_X1  g757(.A1(new_n915), .A2(new_n943), .B1(G952), .B2(G953), .ZN(new_n944));
  INV_X1    g758(.A(new_n934), .ZN(new_n945));
  OR2_X1    g759(.A1(new_n945), .A2(KEYINPUT49), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(KEYINPUT49), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n596), .A2(new_n603), .ZN(new_n948));
  AND3_X1   g762(.A1(new_n946), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n949), .A2(new_n697), .A3(new_n757), .A4(new_n825), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n944), .B1(new_n710), .B2(new_n950), .ZN(G75));
  NOR2_X1   g765(.A1(new_n327), .A2(G952), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT120), .ZN(new_n953));
  INV_X1    g767(.A(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n521), .A2(new_n537), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n955), .B(new_n535), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(KEYINPUT55), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n911), .A2(G210), .A3(G902), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT56), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n957), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  AND3_X1   g774(.A1(new_n911), .A2(KEYINPUT119), .A3(G902), .ZN(new_n961));
  AOI21_X1  g775(.A(KEYINPUT119), .B1(new_n911), .B2(G902), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n963), .A2(new_n488), .ZN(new_n964));
  AND2_X1   g778(.A1(new_n957), .A2(new_n959), .ZN(new_n965));
  AOI211_X1 g779(.A(new_n954), .B(new_n960), .C1(new_n964), .C2(new_n965), .ZN(G51));
  INV_X1    g780(.A(KEYINPUT122), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n967), .B1(new_n963), .B2(new_n815), .ZN(new_n968));
  NOR4_X1   g782(.A1(new_n961), .A2(new_n962), .A3(KEYINPUT122), .A4(new_n814), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n911), .A2(KEYINPUT54), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n912), .A2(KEYINPUT121), .A3(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT121), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n911), .A2(new_n973), .A3(KEYINPUT54), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n591), .B(KEYINPUT57), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n972), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n626), .A2(new_n628), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n952), .B1(new_n970), .B2(new_n978), .ZN(G54));
  AND2_X1   g793(.A1(KEYINPUT58), .A2(G475), .ZN(new_n980));
  AND3_X1   g794(.A1(new_n963), .A2(new_n477), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n477), .B1(new_n963), .B2(new_n980), .ZN(new_n982));
  NOR3_X1   g796(.A1(new_n981), .A2(new_n982), .A3(new_n952), .ZN(G60));
  NAND2_X1  g797(.A1(new_n613), .A2(new_n615), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n611), .B(KEYINPUT59), .Z(new_n985));
  AND4_X1   g799(.A1(new_n984), .A2(new_n972), .A3(new_n974), .A4(new_n985), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n984), .B1(new_n915), .B2(new_n985), .ZN(new_n987));
  NOR3_X1   g801(.A1(new_n986), .A2(new_n954), .A3(new_n987), .ZN(G63));
  XNOR2_X1  g802(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n397), .A2(new_n343), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n989), .B(new_n990), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n911), .A2(new_n668), .A3(new_n991), .ZN(new_n992));
  AND2_X1   g806(.A1(new_n911), .A2(new_n991), .ZN(new_n993));
  OAI211_X1 g807(.A(new_n953), .B(new_n992), .C1(new_n993), .C2(new_n342), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n994), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g809(.A(G953), .B1(new_n422), .B2(new_n528), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n996), .B1(new_n908), .B2(G953), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n955), .B1(G898), .B2(new_n327), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n998), .B(KEYINPUT124), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n997), .B(new_n999), .ZN(G69));
  NOR2_X1   g814(.A1(new_n263), .A2(new_n265), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n1001), .B(new_n471), .ZN(new_n1002));
  INV_X1    g816(.A(new_n1002), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n1003), .B1(new_n684), .B2(new_n327), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n824), .A2(new_n861), .A3(new_n776), .ZN(new_n1005));
  NAND4_X1  g819(.A1(new_n839), .A2(new_n830), .A3(new_n1005), .A4(new_n807), .ZN(new_n1006));
  AND2_X1   g820(.A1(new_n860), .A2(new_n724), .ZN(new_n1007));
  INV_X1    g821(.A(new_n1007), .ZN(new_n1008));
  NOR2_X1   g822(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  AND2_X1   g823(.A1(new_n1009), .A2(new_n802), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n1004), .B1(new_n1010), .B2(new_n327), .ZN(new_n1011));
  XOR2_X1   g825(.A(new_n1002), .B(KEYINPUT125), .Z(new_n1012));
  NAND2_X1  g826(.A1(new_n717), .A2(new_n876), .ZN(new_n1013));
  NAND4_X1  g827(.A1(new_n350), .A2(new_n1013), .A3(new_n704), .A4(new_n778), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n839), .A2(new_n830), .A3(new_n1014), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1007), .A2(new_n712), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1015), .B1(KEYINPUT62), .B2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g831(.A1(new_n1016), .A2(KEYINPUT62), .ZN(new_n1018));
  XOR2_X1   g832(.A(new_n1018), .B(KEYINPUT126), .Z(new_n1019));
  NAND2_X1  g833(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n1012), .B1(new_n1020), .B2(new_n327), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n327), .B1(G227), .B2(G900), .ZN(new_n1022));
  OR3_X1    g836(.A1(new_n1011), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n1022), .B1(new_n1011), .B2(new_n1021), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1023), .A2(new_n1024), .ZN(G72));
  NAND3_X1  g839(.A1(new_n1009), .A2(new_n802), .A3(new_n908), .ZN(new_n1026));
  XNOR2_X1  g840(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n1027));
  NOR2_X1   g841(.A1(new_n187), .A2(new_n343), .ZN(new_n1028));
  XOR2_X1   g842(.A(new_n1027), .B(new_n1028), .Z(new_n1029));
  INV_X1    g843(.A(new_n1029), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1026), .A2(new_n1030), .ZN(new_n1031));
  NOR2_X1   g845(.A1(new_n267), .A2(new_n192), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n952), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n1029), .B1(new_n268), .B2(new_n619), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n913), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g850(.A(new_n1030), .B1(new_n1020), .B2(new_n904), .ZN(new_n1037));
  AOI21_X1  g851(.A(new_n1036), .B1(new_n707), .B2(new_n1037), .ZN(G57));
endmodule


