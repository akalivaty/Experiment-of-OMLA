

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756;

  XNOR2_X1 U361 ( .A(n479), .B(n434), .ZN(n746) );
  XNOR2_X1 U362 ( .A(n741), .B(n460), .ZN(n689) );
  XNOR2_X2 U363 ( .A(G137), .B(KEYINPUT4), .ZN(n381) );
  XNOR2_X2 U364 ( .A(G101), .B(KEYINPUT3), .ZN(n448) );
  XNOR2_X2 U365 ( .A(n430), .B(n449), .ZN(n502) );
  XNOR2_X2 U366 ( .A(G110), .B(G107), .ZN(n430) );
  XNOR2_X2 U367 ( .A(G146), .B(G125), .ZN(n479) );
  XNOR2_X2 U368 ( .A(n527), .B(KEYINPUT33), .ZN(n571) );
  XNOR2_X2 U369 ( .A(n348), .B(n343), .ZN(n657) );
  INV_X2 U370 ( .A(G953), .ZN(n752) );
  XNOR2_X1 U371 ( .A(n592), .B(KEYINPUT102), .ZN(n371) );
  AND2_X1 U372 ( .A1(n439), .A2(n615), .ZN(n723) );
  BUF_X1 U373 ( .A(n700), .Z(n704) );
  NOR2_X1 U374 ( .A1(n661), .A2(n660), .ZN(n665) );
  NAND2_X1 U375 ( .A1(n371), .A2(n582), .ZN(n685) );
  XNOR2_X1 U376 ( .A(n587), .B(KEYINPUT32), .ZN(n682) );
  XNOR2_X1 U377 ( .A(n361), .B(n626), .ZN(n691) );
  XNOR2_X1 U378 ( .A(n359), .B(n617), .ZN(n756) );
  XNOR2_X1 U379 ( .A(n491), .B(n405), .ZN(n616) );
  AND2_X1 U380 ( .A1(n419), .A2(n417), .ZN(n416) );
  BUF_X1 U381 ( .A(n545), .Z(n618) );
  XNOR2_X1 U382 ( .A(n432), .B(n431), .ZN(n376) );
  XNOR2_X1 U383 ( .A(n448), .B(G119), .ZN(n432) );
  XNOR2_X1 U384 ( .A(n433), .B(G131), .ZN(n492) );
  NAND2_X1 U385 ( .A1(n416), .A2(n413), .ZN(n633) );
  NOR2_X1 U386 ( .A1(n365), .A2(n364), .ZN(n354) );
  NAND2_X1 U387 ( .A1(n643), .A2(n734), .ZN(n364) );
  NOR2_X1 U388 ( .A1(n625), .A2(n447), .ZN(n435) );
  AND2_X1 U389 ( .A1(n546), .A2(n598), .ZN(n399) );
  OR2_X1 U390 ( .A1(n689), .A2(n424), .ZN(n423) );
  NAND2_X1 U391 ( .A1(n426), .A2(n425), .ZN(n424) );
  INV_X1 U392 ( .A(n671), .ZN(n425) );
  INV_X1 U393 ( .A(n464), .ZN(n426) );
  XNOR2_X1 U394 ( .A(n367), .B(n620), .ZN(n624) );
  XNOR2_X1 U395 ( .A(G116), .B(G113), .ZN(n431) );
  NAND2_X1 U396 ( .A1(n618), .A2(n441), .ZN(n440) );
  NOR2_X1 U397 ( .A1(n614), .A2(n442), .ZN(n441) );
  INV_X1 U398 ( .A(n628), .ZN(n442) );
  NOR2_X1 U399 ( .A1(n588), .A2(n377), .ZN(n589) );
  XNOR2_X1 U400 ( .A(n350), .B(KEYINPUT70), .ZN(n349) );
  NAND2_X1 U401 ( .A1(n368), .A2(n370), .ZN(n350) );
  AND2_X1 U402 ( .A1(n685), .A2(n682), .ZN(n370) );
  XNOR2_X1 U403 ( .A(n369), .B(KEYINPUT65), .ZN(n368) );
  XNOR2_X1 U404 ( .A(KEYINPUT15), .B(G902), .ZN(n506) );
  XOR2_X1 U405 ( .A(KEYINPUT68), .B(KEYINPUT48), .Z(n446) );
  XNOR2_X1 U406 ( .A(KEYINPUT10), .B(G140), .ZN(n434) );
  XNOR2_X1 U407 ( .A(n380), .B(n492), .ZN(n375) );
  XNOR2_X1 U408 ( .A(n381), .B(n406), .ZN(n380) );
  INV_X1 U409 ( .A(KEYINPUT67), .ZN(n406) );
  INV_X1 U410 ( .A(n506), .ZN(n671) );
  XNOR2_X1 U411 ( .A(n495), .B(KEYINPUT93), .ZN(n496) );
  XNOR2_X1 U412 ( .A(G128), .B(KEYINPUT78), .ZN(n519) );
  XNOR2_X1 U413 ( .A(G110), .B(KEYINPUT24), .ZN(n520) );
  XNOR2_X1 U414 ( .A(KEYINPUT87), .B(KEYINPUT23), .ZN(n514) );
  XNOR2_X1 U415 ( .A(G119), .B(KEYINPUT73), .ZN(n363) );
  INV_X1 U416 ( .A(KEYINPUT8), .ZN(n473) );
  XNOR2_X1 U417 ( .A(n407), .B(G101), .ZN(n374) );
  INV_X1 U418 ( .A(G140), .ZN(n407) );
  INV_X1 U419 ( .A(G104), .ZN(n449) );
  AND2_X1 U420 ( .A1(n534), .A2(n575), .ZN(n627) );
  NAND2_X1 U421 ( .A1(n387), .A2(n382), .ZN(n655) );
  NOR2_X1 U422 ( .A1(n385), .A2(n384), .ZN(n383) );
  AND2_X1 U423 ( .A1(n624), .A2(n436), .ZN(n366) );
  AND2_X1 U424 ( .A1(n692), .A2(n523), .ZN(n362) );
  NAND2_X1 U425 ( .A1(n616), .A2(n723), .ZN(n359) );
  NAND2_X1 U426 ( .A1(n756), .A2(KEYINPUT46), .ZN(n358) );
  XOR2_X1 U427 ( .A(KEYINPUT89), .B(KEYINPUT20), .Z(n508) );
  AND2_X1 U428 ( .A1(n356), .A2(n606), .ZN(n351) );
  INV_X1 U429 ( .A(KEYINPUT66), .ZN(n433) );
  XNOR2_X1 U430 ( .A(G113), .B(G143), .ZN(n483) );
  XOR2_X1 U431 ( .A(G122), .B(G104), .Z(n484) );
  XNOR2_X1 U432 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n455) );
  XNOR2_X1 U433 ( .A(KEYINPUT18), .B(KEYINPUT84), .ZN(n453) );
  XNOR2_X1 U434 ( .A(KEYINPUT75), .B(KEYINPUT76), .ZN(n452) );
  NAND2_X1 U435 ( .A1(n389), .A2(KEYINPUT39), .ZN(n388) );
  NOR2_X1 U436 ( .A1(n422), .A2(n562), .ZN(n421) );
  INV_X1 U437 ( .A(n427), .ZN(n422) );
  NOR2_X1 U438 ( .A1(n428), .A2(n563), .ZN(n418) );
  XNOR2_X1 U439 ( .A(n615), .B(KEYINPUT1), .ZN(n546) );
  INV_X1 U440 ( .A(G902), .ZN(n523) );
  BUF_X1 U441 ( .A(n657), .Z(n735) );
  XNOR2_X1 U442 ( .A(G116), .B(G107), .ZN(n470) );
  XNOR2_X1 U443 ( .A(n472), .B(G134), .ZN(n493) );
  BUF_X1 U444 ( .A(n662), .Z(n394) );
  INV_X1 U445 ( .A(KEYINPUT41), .ZN(n405) );
  XNOR2_X1 U446 ( .A(n633), .B(n564), .ZN(n724) );
  XNOR2_X1 U447 ( .A(n599), .B(KEYINPUT92), .ZN(n622) );
  INV_X1 U448 ( .A(n594), .ZN(n602) );
  BUF_X1 U449 ( .A(n618), .Z(n600) );
  XNOR2_X1 U450 ( .A(n496), .B(n497), .ZN(n444) );
  XNOR2_X1 U451 ( .A(n429), .B(n376), .ZN(n741) );
  XNOR2_X1 U452 ( .A(n502), .B(n451), .ZN(n429) );
  XNOR2_X1 U453 ( .A(KEYINPUT72), .B(KEYINPUT16), .ZN(n450) );
  XNOR2_X1 U454 ( .A(n438), .B(n437), .ZN(n692) );
  XNOR2_X1 U455 ( .A(n522), .B(n521), .ZN(n437) );
  XNOR2_X1 U456 ( .A(n516), .B(n517), .ZN(n438) );
  XNOR2_X1 U457 ( .A(n379), .B(n372), .ZN(n707) );
  XNOR2_X1 U458 ( .A(n373), .B(n503), .ZN(n372) );
  XNOR2_X1 U459 ( .A(n502), .B(n374), .ZN(n373) );
  XNOR2_X1 U460 ( .A(KEYINPUT111), .B(KEYINPUT40), .ZN(n626) );
  INV_X1 U461 ( .A(KEYINPUT35), .ZN(n378) );
  XNOR2_X1 U462 ( .A(n440), .B(n342), .ZN(n439) );
  NAND2_X1 U463 ( .A1(n386), .A2(n366), .ZN(n641) );
  BUF_X1 U464 ( .A(n724), .Z(n357) );
  INV_X1 U465 ( .A(n696), .ZN(n697) );
  INV_X1 U466 ( .A(KEYINPUT60), .ZN(n397) );
  INV_X1 U467 ( .A(n625), .ZN(n537) );
  XNOR2_X1 U468 ( .A(n622), .B(n621), .ZN(n623) );
  XOR2_X1 U469 ( .A(KEYINPUT79), .B(n735), .Z(n339) );
  AND2_X2 U470 ( .A1(n576), .A2(n614), .ZN(n598) );
  AND2_X1 U471 ( .A1(n423), .A2(n427), .ZN(n340) );
  NOR2_X1 U472 ( .A1(n575), .A2(n574), .ZN(n341) );
  XOR2_X1 U473 ( .A(KEYINPUT28), .B(KEYINPUT110), .Z(n342) );
  INV_X1 U474 ( .A(KEYINPUT39), .ZN(n391) );
  XNOR2_X1 U475 ( .A(KEYINPUT81), .B(KEYINPUT45), .ZN(n343) );
  XOR2_X1 U476 ( .A(n702), .B(n701), .Z(n344) );
  XOR2_X1 U477 ( .A(n689), .B(n688), .Z(n345) );
  XOR2_X1 U478 ( .A(n676), .B(n678), .Z(n346) );
  NOR2_X1 U479 ( .A1(n752), .A2(G952), .ZN(n710) );
  INV_X1 U480 ( .A(n710), .ZN(n400) );
  XOR2_X1 U481 ( .A(KEYINPUT122), .B(KEYINPUT56), .Z(n347) );
  NAND2_X1 U482 ( .A1(n351), .A2(n349), .ZN(n348) );
  XNOR2_X1 U483 ( .A(n352), .B(n446), .ZN(n355) );
  NAND2_X1 U484 ( .A1(n354), .A2(n353), .ZN(n352) );
  NAND2_X1 U485 ( .A1(n393), .A2(n392), .ZN(n353) );
  NAND2_X1 U486 ( .A1(n355), .A2(n652), .ZN(n654) );
  NAND2_X1 U487 ( .A1(n691), .A2(KEYINPUT46), .ZN(n360) );
  NAND2_X1 U488 ( .A1(n590), .A2(KEYINPUT44), .ZN(n356) );
  NAND2_X1 U489 ( .A1(n420), .A2(KEYINPUT83), .ZN(n419) );
  NAND2_X1 U490 ( .A1(n423), .A2(n421), .ZN(n420) );
  AND2_X1 U491 ( .A1(n390), .A2(n388), .ZN(n387) );
  NAND2_X1 U492 ( .A1(n360), .A2(n358), .ZN(n365) );
  NAND2_X1 U493 ( .A1(n624), .A2(n435), .ZN(n389) );
  NAND2_X1 U494 ( .A1(n618), .A2(n644), .ZN(n367) );
  NAND2_X1 U495 ( .A1(n415), .A2(n414), .ZN(n413) );
  AND2_X2 U496 ( .A1(n586), .A2(n525), .ZN(n592) );
  NAND2_X1 U497 ( .A1(n655), .A2(n627), .ZN(n361) );
  XNOR2_X2 U498 ( .A(n362), .B(n524), .ZN(n614) );
  XNOR2_X1 U499 ( .A(n363), .B(G137), .ZN(n515) );
  NAND2_X1 U500 ( .A1(n409), .A2(n408), .ZN(n369) );
  XNOR2_X2 U501 ( .A(n581), .B(n580), .ZN(n586) );
  XNOR2_X2 U502 ( .A(n747), .B(G146), .ZN(n379) );
  XNOR2_X2 U503 ( .A(n375), .B(n493), .ZN(n747) );
  XNOR2_X1 U504 ( .A(n444), .B(n376), .ZN(n443) );
  INV_X1 U505 ( .A(n409), .ZN(n377) );
  XNOR2_X1 U506 ( .A(n409), .B(G122), .ZN(G24) );
  XNOR2_X2 U507 ( .A(n410), .B(n378), .ZN(n409) );
  XNOR2_X1 U508 ( .A(n379), .B(n443), .ZN(n676) );
  NAND2_X1 U509 ( .A1(n623), .A2(KEYINPUT39), .ZN(n390) );
  NAND2_X1 U510 ( .A1(n386), .A2(n383), .ZN(n382) );
  NAND2_X1 U511 ( .A1(n435), .A2(n391), .ZN(n384) );
  INV_X1 U512 ( .A(n624), .ZN(n385) );
  INV_X1 U513 ( .A(n623), .ZN(n386) );
  NOR2_X1 U514 ( .A1(n756), .A2(KEYINPUT46), .ZN(n392) );
  INV_X1 U515 ( .A(n691), .ZN(n393) );
  NAND2_X1 U516 ( .A1(n656), .A2(n684), .ZN(n662) );
  NOR2_X2 U517 ( .A1(n662), .A2(n657), .ZN(n673) );
  NOR2_X2 U518 ( .A1(n673), .A2(KEYINPUT80), .ZN(n672) );
  XNOR2_X1 U519 ( .A(n395), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U520 ( .A1(n402), .A2(n400), .ZN(n395) );
  XNOR2_X1 U521 ( .A(n396), .B(n347), .ZN(G51) );
  NAND2_X1 U522 ( .A1(n403), .A2(n400), .ZN(n396) );
  XNOR2_X1 U523 ( .A(n398), .B(n397), .ZN(G60) );
  NAND2_X1 U524 ( .A1(n401), .A2(n400), .ZN(n398) );
  NAND2_X1 U525 ( .A1(n399), .A2(n526), .ZN(n527) );
  XNOR2_X1 U526 ( .A(n703), .B(n344), .ZN(n401) );
  XNOR2_X1 U527 ( .A(n679), .B(n346), .ZN(n402) );
  XNOR2_X1 U528 ( .A(n690), .B(n345), .ZN(n403) );
  NAND2_X1 U529 ( .A1(n615), .A2(n598), .ZN(n599) );
  XNOR2_X2 U530 ( .A(n505), .B(n504), .ZN(n615) );
  XNOR2_X2 U531 ( .A(n404), .B(KEYINPUT0), .ZN(n594) );
  NOR2_X2 U532 ( .A1(n724), .A2(n570), .ZN(n404) );
  XNOR2_X2 U533 ( .A(n672), .B(n671), .ZN(n675) );
  INV_X1 U534 ( .A(KEYINPUT44), .ZN(n408) );
  NAND2_X1 U535 ( .A1(n411), .A2(n341), .ZN(n410) );
  XNOR2_X1 U536 ( .A(n572), .B(n412), .ZN(n411) );
  INV_X1 U537 ( .A(KEYINPUT34), .ZN(n412) );
  AND2_X1 U538 ( .A1(n428), .A2(n563), .ZN(n414) );
  INV_X1 U539 ( .A(n420), .ZN(n415) );
  INV_X1 U540 ( .A(n418), .ZN(n417) );
  NAND2_X1 U541 ( .A1(n428), .A2(n340), .ZN(n651) );
  NAND2_X1 U542 ( .A1(n464), .A2(n671), .ZN(n427) );
  NAND2_X1 U543 ( .A1(n689), .A2(n464), .ZN(n428) );
  INV_X1 U544 ( .A(n647), .ZN(n525) );
  NOR2_X2 U545 ( .A1(G902), .A2(n707), .ZN(n505) );
  INV_X1 U546 ( .A(n447), .ZN(n436) );
  XOR2_X1 U547 ( .A(KEYINPUT53), .B(n670), .Z(G75) );
  NOR2_X1 U548 ( .A1(n612), .A2(n611), .ZN(n447) );
  XNOR2_X1 U549 ( .A(KEYINPUT69), .B(G469), .ZN(n504) );
  INV_X1 U550 ( .A(KEYINPUT83), .ZN(n563) );
  INV_X1 U551 ( .A(n692), .ZN(n693) );
  XNOR2_X1 U552 ( .A(n450), .B(G122), .ZN(n451) );
  XNOR2_X1 U553 ( .A(n453), .B(n452), .ZN(n457) );
  NAND2_X1 U554 ( .A1(n752), .A2(G224), .ZN(n454) );
  XNOR2_X1 U555 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U556 ( .A(n457), .B(n456), .ZN(n459) );
  XNOR2_X1 U557 ( .A(G128), .B(G143), .ZN(n472) );
  XNOR2_X1 U558 ( .A(n479), .B(n472), .ZN(n458) );
  XNOR2_X1 U559 ( .A(n459), .B(n458), .ZN(n460) );
  INV_X1 U560 ( .A(G237), .ZN(n461) );
  NAND2_X1 U561 ( .A1(n523), .A2(n461), .ZN(n466) );
  NAND2_X1 U562 ( .A1(n466), .A2(G210), .ZN(n463) );
  INV_X1 U563 ( .A(KEYINPUT77), .ZN(n462) );
  XNOR2_X1 U564 ( .A(n463), .B(n462), .ZN(n464) );
  INV_X1 U565 ( .A(KEYINPUT38), .ZN(n465) );
  XNOR2_X1 U566 ( .A(n651), .B(n465), .ZN(n625) );
  NAND2_X1 U567 ( .A1(n466), .A2(G214), .ZN(n644) );
  NAND2_X1 U568 ( .A1(n537), .A2(n644), .ZN(n535) );
  XOR2_X1 U569 ( .A(KEYINPUT100), .B(KEYINPUT9), .Z(n468) );
  XNOR2_X1 U570 ( .A(G122), .B(KEYINPUT99), .ZN(n467) );
  XNOR2_X1 U571 ( .A(n468), .B(n467), .ZN(n469) );
  XOR2_X1 U572 ( .A(n469), .B(KEYINPUT7), .Z(n471) );
  XNOR2_X1 U573 ( .A(n471), .B(n470), .ZN(n477) );
  NAND2_X1 U574 ( .A1(G234), .A2(n752), .ZN(n474) );
  XNOR2_X1 U575 ( .A(n474), .B(n473), .ZN(n518) );
  NAND2_X1 U576 ( .A1(n518), .A2(G217), .ZN(n475) );
  XNOR2_X1 U577 ( .A(n493), .B(n475), .ZN(n476) );
  XNOR2_X1 U578 ( .A(n477), .B(n476), .ZN(n696) );
  NAND2_X1 U579 ( .A1(n696), .A2(n523), .ZN(n478) );
  XNOR2_X1 U580 ( .A(n478), .B(G478), .ZN(n533) );
  XNOR2_X1 U581 ( .A(n492), .B(KEYINPUT97), .ZN(n480) );
  XNOR2_X1 U582 ( .A(n480), .B(n746), .ZN(n488) );
  XOR2_X1 U583 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n482) );
  NOR2_X1 U584 ( .A1(G953), .A2(G237), .ZN(n494) );
  NAND2_X1 U585 ( .A1(G214), .A2(n494), .ZN(n481) );
  XNOR2_X1 U586 ( .A(n482), .B(n481), .ZN(n486) );
  XNOR2_X1 U587 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U588 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U589 ( .A(n488), .B(n487), .ZN(n702) );
  NAND2_X1 U590 ( .A1(n702), .A2(n523), .ZN(n490) );
  XOR2_X1 U591 ( .A(KEYINPUT13), .B(G475), .Z(n489) );
  XNOR2_X1 U592 ( .A(n490), .B(n489), .ZN(n573) );
  OR2_X1 U593 ( .A1(n533), .A2(n573), .ZN(n578) );
  NOR2_X1 U594 ( .A1(n535), .A2(n578), .ZN(n491) );
  NAND2_X1 U595 ( .A1(n494), .A2(G210), .ZN(n495) );
  XOR2_X1 U596 ( .A(KEYINPUT5), .B(KEYINPUT94), .Z(n497) );
  NAND2_X1 U597 ( .A1(n676), .A2(n523), .ZN(n500) );
  INV_X1 U598 ( .A(KEYINPUT95), .ZN(n498) );
  XNOR2_X1 U599 ( .A(n498), .B(G472), .ZN(n499) );
  XNOR2_X2 U600 ( .A(n500), .B(n499), .ZN(n545) );
  XNOR2_X1 U601 ( .A(n545), .B(KEYINPUT6), .ZN(n583) );
  INV_X1 U602 ( .A(n583), .ZN(n526) );
  NAND2_X1 U603 ( .A1(G227), .A2(n752), .ZN(n501) );
  XNOR2_X1 U604 ( .A(KEYINPUT74), .B(n501), .ZN(n503) );
  NAND2_X1 U605 ( .A1(G234), .A2(n506), .ZN(n507) );
  XNOR2_X1 U606 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U607 ( .A(n509), .B(KEYINPUT88), .ZN(n511) );
  NAND2_X1 U608 ( .A1(n511), .A2(G221), .ZN(n510) );
  XNOR2_X1 U609 ( .A(n510), .B(KEYINPUT21), .ZN(n613) );
  XNOR2_X1 U610 ( .A(n613), .B(KEYINPUT91), .ZN(n576) );
  NAND2_X1 U611 ( .A1(n511), .A2(G217), .ZN(n513) );
  XNOR2_X1 U612 ( .A(KEYINPUT90), .B(KEYINPUT25), .ZN(n512) );
  XNOR2_X1 U613 ( .A(n513), .B(n512), .ZN(n524) );
  INV_X1 U614 ( .A(n746), .ZN(n517) );
  XNOR2_X1 U615 ( .A(n515), .B(n514), .ZN(n516) );
  NAND2_X1 U616 ( .A1(n518), .A2(G221), .ZN(n522) );
  XNOR2_X1 U617 ( .A(n520), .B(n519), .ZN(n521) );
  BUF_X1 U618 ( .A(n571), .Z(n528) );
  NAND2_X1 U619 ( .A1(n616), .A2(n528), .ZN(n529) );
  AND2_X1 U620 ( .A1(n529), .A2(n752), .ZN(n669) );
  NAND2_X1 U621 ( .A1(G234), .A2(G237), .ZN(n530) );
  XNOR2_X1 U622 ( .A(n530), .B(KEYINPUT14), .ZN(n566) );
  NAND2_X1 U623 ( .A1(G952), .A2(n566), .ZN(n567) );
  INV_X1 U624 ( .A(KEYINPUT98), .ZN(n531) );
  XNOR2_X1 U625 ( .A(n573), .B(n531), .ZN(n532) );
  AND2_X1 U626 ( .A1(n532), .A2(n533), .ZN(n729) );
  INV_X1 U627 ( .A(n532), .ZN(n534) );
  INV_X1 U628 ( .A(n533), .ZN(n575) );
  OR2_X1 U629 ( .A1(n729), .A2(n627), .ZN(n636) );
  INV_X1 U630 ( .A(n636), .ZN(n603) );
  NOR2_X1 U631 ( .A1(n603), .A2(n535), .ZN(n536) );
  XOR2_X1 U632 ( .A(KEYINPUT119), .B(n536), .Z(n541) );
  NOR2_X1 U633 ( .A1(n537), .A2(n644), .ZN(n538) );
  NOR2_X1 U634 ( .A1(n578), .A2(n538), .ZN(n539) );
  XNOR2_X1 U635 ( .A(KEYINPUT118), .B(n539), .ZN(n540) );
  NOR2_X1 U636 ( .A1(n541), .A2(n540), .ZN(n543) );
  INV_X1 U637 ( .A(n528), .ZN(n542) );
  NOR2_X1 U638 ( .A1(n543), .A2(n542), .ZN(n557) );
  INV_X1 U639 ( .A(n614), .ZN(n629) );
  NAND2_X1 U640 ( .A1(n629), .A2(n613), .ZN(n544) );
  XOR2_X1 U641 ( .A(KEYINPUT49), .B(n544), .Z(n550) );
  BUF_X1 U642 ( .A(n546), .Z(n647) );
  NOR2_X1 U643 ( .A1(n598), .A2(n647), .ZN(n547) );
  XNOR2_X1 U644 ( .A(KEYINPUT50), .B(n547), .ZN(n548) );
  NOR2_X1 U645 ( .A1(n600), .A2(n548), .ZN(n549) );
  NAND2_X1 U646 ( .A1(n550), .A2(n549), .ZN(n552) );
  AND2_X1 U647 ( .A1(n600), .A2(n647), .ZN(n551) );
  NAND2_X1 U648 ( .A1(n598), .A2(n551), .ZN(n595) );
  NAND2_X1 U649 ( .A1(n552), .A2(n595), .ZN(n553) );
  XNOR2_X1 U650 ( .A(KEYINPUT51), .B(n553), .ZN(n555) );
  INV_X1 U651 ( .A(n616), .ZN(n554) );
  NOR2_X1 U652 ( .A1(n555), .A2(n554), .ZN(n556) );
  NOR2_X1 U653 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U654 ( .A(n558), .B(KEYINPUT120), .Z(n559) );
  XOR2_X1 U655 ( .A(KEYINPUT52), .B(n559), .Z(n560) );
  NOR2_X1 U656 ( .A1(n567), .A2(n560), .ZN(n561) );
  XOR2_X1 U657 ( .A(KEYINPUT121), .B(n561), .Z(n667) );
  INV_X1 U658 ( .A(n644), .ZN(n562) );
  XNOR2_X1 U659 ( .A(KEYINPUT64), .B(KEYINPUT19), .ZN(n564) );
  NOR2_X1 U660 ( .A1(G898), .A2(n752), .ZN(n565) );
  XOR2_X1 U661 ( .A(KEYINPUT86), .B(n565), .Z(n742) );
  NAND2_X1 U662 ( .A1(G902), .A2(n566), .ZN(n607) );
  OR2_X1 U663 ( .A1(n742), .A2(n607), .ZN(n569) );
  NOR2_X1 U664 ( .A1(G953), .A2(n567), .ZN(n568) );
  XNOR2_X1 U665 ( .A(n568), .B(KEYINPUT85), .ZN(n610) );
  AND2_X1 U666 ( .A1(n569), .A2(n610), .ZN(n570) );
  NAND2_X1 U667 ( .A1(n571), .A2(n594), .ZN(n572) );
  INV_X1 U668 ( .A(n573), .ZN(n574) );
  INV_X1 U669 ( .A(n576), .ZN(n577) );
  NOR2_X1 U670 ( .A1(n578), .A2(n577), .ZN(n579) );
  NAND2_X1 U671 ( .A1(n594), .A2(n579), .ZN(n581) );
  XNOR2_X1 U672 ( .A(KEYINPUT71), .B(KEYINPUT22), .ZN(n580) );
  NOR2_X1 U673 ( .A1(n614), .A2(n600), .ZN(n582) );
  NAND2_X1 U674 ( .A1(n629), .A2(n647), .ZN(n584) );
  NOR2_X1 U675 ( .A1(n526), .A2(n584), .ZN(n585) );
  NAND2_X1 U676 ( .A1(n586), .A2(n585), .ZN(n587) );
  INV_X1 U677 ( .A(n682), .ZN(n588) );
  NAND2_X1 U678 ( .A1(n589), .A2(n685), .ZN(n590) );
  NOR2_X1 U679 ( .A1(n526), .A2(n629), .ZN(n591) );
  NAND2_X1 U680 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U681 ( .A(n593), .B(KEYINPUT101), .ZN(n686) );
  NOR2_X1 U682 ( .A1(n602), .A2(n595), .ZN(n597) );
  XOR2_X1 U683 ( .A(KEYINPUT96), .B(KEYINPUT31), .Z(n596) );
  XNOR2_X1 U684 ( .A(n597), .B(n596), .ZN(n730) );
  OR2_X1 U685 ( .A1(n622), .A2(n600), .ZN(n601) );
  NOR2_X1 U686 ( .A1(n602), .A2(n601), .ZN(n715) );
  NOR2_X1 U687 ( .A1(n730), .A2(n715), .ZN(n604) );
  NOR2_X1 U688 ( .A1(n604), .A2(n603), .ZN(n605) );
  NOR2_X1 U689 ( .A1(n686), .A2(n605), .ZN(n606) );
  NOR2_X1 U690 ( .A1(n339), .A2(KEYINPUT2), .ZN(n661) );
  OR2_X1 U691 ( .A1(n752), .A2(n607), .ZN(n608) );
  XNOR2_X1 U692 ( .A(KEYINPUT104), .B(n608), .ZN(n609) );
  NOR2_X1 U693 ( .A1(G900), .A2(n609), .ZN(n612) );
  INV_X1 U694 ( .A(n610), .ZN(n611) );
  NOR2_X1 U695 ( .A1(n613), .A2(n447), .ZN(n628) );
  INV_X1 U696 ( .A(KEYINPUT42), .ZN(n617) );
  XNOR2_X1 U697 ( .A(KEYINPUT108), .B(KEYINPUT109), .ZN(n619) );
  XNOR2_X1 U698 ( .A(n619), .B(KEYINPUT30), .ZN(n620) );
  INV_X1 U699 ( .A(KEYINPUT107), .ZN(n621) );
  XNOR2_X1 U700 ( .A(n627), .B(KEYINPUT103), .ZN(n712) );
  NAND2_X1 U701 ( .A1(n629), .A2(n628), .ZN(n630) );
  NOR2_X1 U702 ( .A1(n630), .A2(n583), .ZN(n631) );
  XNOR2_X1 U703 ( .A(n631), .B(KEYINPUT105), .ZN(n632) );
  NOR2_X1 U704 ( .A1(n712), .A2(n632), .ZN(n645) );
  AND2_X1 U705 ( .A1(n645), .A2(n633), .ZN(n634) );
  XNOR2_X1 U706 ( .A(n634), .B(KEYINPUT36), .ZN(n635) );
  NAND2_X1 U707 ( .A1(n635), .A2(n647), .ZN(n734) );
  NAND2_X1 U708 ( .A1(n723), .A2(n636), .ZN(n637) );
  NOR2_X1 U709 ( .A1(n637), .A2(n357), .ZN(n638) );
  XNOR2_X1 U710 ( .A(n638), .B(KEYINPUT47), .ZN(n642) );
  INV_X1 U711 ( .A(n651), .ZN(n639) );
  NAND2_X1 U712 ( .A1(n341), .A2(n639), .ZN(n640) );
  OR2_X1 U713 ( .A1(n641), .A2(n640), .ZN(n680) );
  AND2_X1 U714 ( .A1(n642), .A2(n680), .ZN(n643) );
  NAND2_X1 U715 ( .A1(n645), .A2(n644), .ZN(n646) );
  OR2_X1 U716 ( .A1(n647), .A2(n646), .ZN(n649) );
  XNOR2_X1 U717 ( .A(KEYINPUT43), .B(KEYINPUT106), .ZN(n648) );
  XNOR2_X1 U718 ( .A(n649), .B(n648), .ZN(n650) );
  AND2_X1 U719 ( .A1(n651), .A2(n650), .ZN(n687) );
  INV_X1 U720 ( .A(n687), .ZN(n652) );
  INV_X1 U721 ( .A(KEYINPUT82), .ZN(n653) );
  XNOR2_X1 U722 ( .A(n654), .B(n653), .ZN(n656) );
  NAND2_X1 U723 ( .A1(n655), .A2(n729), .ZN(n684) );
  INV_X1 U724 ( .A(KEYINPUT79), .ZN(n658) );
  NAND2_X1 U725 ( .A1(n658), .A2(KEYINPUT2), .ZN(n659) );
  NOR2_X1 U726 ( .A1(n673), .A2(n659), .ZN(n660) );
  INV_X1 U727 ( .A(n394), .ZN(n663) );
  NOR2_X1 U728 ( .A1(n663), .A2(KEYINPUT2), .ZN(n664) );
  NOR2_X1 U729 ( .A1(n665), .A2(n664), .ZN(n666) );
  NOR2_X1 U730 ( .A1(n667), .A2(n666), .ZN(n668) );
  NAND2_X1 U731 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U732 ( .A(n673), .B(KEYINPUT2), .ZN(n674) );
  NOR2_X4 U733 ( .A1(n675), .A2(n674), .ZN(n700) );
  NAND2_X1 U734 ( .A1(n700), .A2(G472), .ZN(n679) );
  XNOR2_X1 U735 ( .A(KEYINPUT112), .B(KEYINPUT113), .ZN(n677) );
  XNOR2_X1 U736 ( .A(n677), .B(KEYINPUT62), .ZN(n678) );
  XNOR2_X1 U737 ( .A(n680), .B(G143), .ZN(G45) );
  XOR2_X1 U738 ( .A(G119), .B(KEYINPUT127), .Z(n681) );
  XNOR2_X1 U739 ( .A(n682), .B(n681), .ZN(G21) );
  XOR2_X1 U740 ( .A(G134), .B(KEYINPUT117), .Z(n683) );
  XNOR2_X1 U741 ( .A(n684), .B(n683), .ZN(G36) );
  XNOR2_X1 U742 ( .A(n685), .B(G110), .ZN(G12) );
  XOR2_X1 U743 ( .A(G101), .B(n686), .Z(G3) );
  XOR2_X1 U744 ( .A(G140), .B(n687), .Z(G42) );
  NAND2_X1 U745 ( .A1(n700), .A2(G210), .ZN(n690) );
  XOR2_X1 U746 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n688) );
  XOR2_X1 U747 ( .A(n691), .B(G131), .Z(G33) );
  NAND2_X1 U748 ( .A1(n704), .A2(G217), .ZN(n694) );
  XNOR2_X1 U749 ( .A(n694), .B(n693), .ZN(n695) );
  NOR2_X1 U750 ( .A1(n695), .A2(n710), .ZN(G66) );
  NAND2_X1 U751 ( .A1(n704), .A2(G478), .ZN(n698) );
  XNOR2_X1 U752 ( .A(n698), .B(n697), .ZN(n699) );
  NOR2_X1 U753 ( .A1(n699), .A2(n710), .ZN(G63) );
  NAND2_X1 U754 ( .A1(n700), .A2(G475), .ZN(n703) );
  XNOR2_X1 U755 ( .A(KEYINPUT124), .B(KEYINPUT59), .ZN(n701) );
  NAND2_X1 U756 ( .A1(n704), .A2(G469), .ZN(n709) );
  XNOR2_X1 U757 ( .A(KEYINPUT123), .B(KEYINPUT57), .ZN(n705) );
  XNOR2_X1 U758 ( .A(n705), .B(KEYINPUT58), .ZN(n706) );
  XNOR2_X1 U759 ( .A(n707), .B(n706), .ZN(n708) );
  XNOR2_X1 U760 ( .A(n709), .B(n708), .ZN(n711) );
  NOR2_X1 U761 ( .A1(n711), .A2(n710), .ZN(G54) );
  INV_X1 U762 ( .A(n712), .ZN(n727) );
  NAND2_X1 U763 ( .A1(n715), .A2(n727), .ZN(n713) );
  XNOR2_X1 U764 ( .A(n713), .B(KEYINPUT114), .ZN(n714) );
  XNOR2_X1 U765 ( .A(G104), .B(n714), .ZN(G6) );
  XOR2_X1 U766 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n717) );
  NAND2_X1 U767 ( .A1(n715), .A2(n729), .ZN(n716) );
  XNOR2_X1 U768 ( .A(n717), .B(n716), .ZN(n718) );
  XNOR2_X1 U769 ( .A(G107), .B(n718), .ZN(G9) );
  NAND2_X1 U770 ( .A1(n723), .A2(n729), .ZN(n719) );
  NOR2_X1 U771 ( .A1(n719), .A2(n357), .ZN(n721) );
  XNOR2_X1 U772 ( .A(KEYINPUT115), .B(KEYINPUT29), .ZN(n720) );
  XNOR2_X1 U773 ( .A(n721), .B(n720), .ZN(n722) );
  XOR2_X1 U774 ( .A(G128), .B(n722), .Z(G30) );
  NAND2_X1 U775 ( .A1(n723), .A2(n727), .ZN(n725) );
  NOR2_X1 U776 ( .A1(n725), .A2(n357), .ZN(n726) );
  XOR2_X1 U777 ( .A(G146), .B(n726), .Z(G48) );
  NAND2_X1 U778 ( .A1(n730), .A2(n727), .ZN(n728) );
  XNOR2_X1 U779 ( .A(n728), .B(G113), .ZN(G15) );
  NAND2_X1 U780 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U781 ( .A(n731), .B(KEYINPUT116), .ZN(n732) );
  XNOR2_X1 U782 ( .A(G116), .B(n732), .ZN(G18) );
  XOR2_X1 U783 ( .A(G125), .B(KEYINPUT37), .Z(n733) );
  XNOR2_X1 U784 ( .A(n734), .B(n733), .ZN(G27) );
  INV_X1 U785 ( .A(n735), .ZN(n736) );
  NAND2_X1 U786 ( .A1(n736), .A2(n752), .ZN(n740) );
  NAND2_X1 U787 ( .A1(G953), .A2(G224), .ZN(n737) );
  XNOR2_X1 U788 ( .A(KEYINPUT61), .B(n737), .ZN(n738) );
  NAND2_X1 U789 ( .A1(n738), .A2(G898), .ZN(n739) );
  NAND2_X1 U790 ( .A1(n740), .A2(n739), .ZN(n745) );
  XOR2_X1 U791 ( .A(KEYINPUT125), .B(n741), .Z(n743) );
  NAND2_X1 U792 ( .A1(n743), .A2(n742), .ZN(n744) );
  XOR2_X1 U793 ( .A(n745), .B(n744), .Z(G69) );
  XNOR2_X1 U794 ( .A(n747), .B(n746), .ZN(n751) );
  XNOR2_X1 U795 ( .A(n751), .B(G227), .ZN(n748) );
  NAND2_X1 U796 ( .A1(n748), .A2(G900), .ZN(n749) );
  NAND2_X1 U797 ( .A1(G953), .A2(n749), .ZN(n750) );
  XNOR2_X1 U798 ( .A(n750), .B(KEYINPUT126), .ZN(n755) );
  XNOR2_X1 U799 ( .A(n394), .B(n751), .ZN(n753) );
  NAND2_X1 U800 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U801 ( .A1(n755), .A2(n754), .ZN(G72) );
  XOR2_X1 U802 ( .A(G137), .B(n756), .Z(G39) );
endmodule

