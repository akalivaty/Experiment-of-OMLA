

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594;

  XNOR2_X1 U324 ( .A(n356), .B(KEYINPUT45), .ZN(n357) );
  AND2_X1 U325 ( .A1(n576), .A2(n442), .ZN(n443) );
  XNOR2_X1 U326 ( .A(n350), .B(n349), .ZN(n353) );
  XNOR2_X1 U327 ( .A(KEYINPUT46), .B(KEYINPUT110), .ZN(n394) );
  XNOR2_X1 U328 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U329 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U330 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U331 ( .A(KEYINPUT76), .B(G36GAT), .Z(n337) );
  XNOR2_X1 U332 ( .A(n319), .B(n318), .ZN(n321) );
  XOR2_X1 U333 ( .A(n370), .B(n369), .Z(n582) );
  XOR2_X1 U334 ( .A(n329), .B(n328), .Z(n587) );
  INV_X1 U335 ( .A(G190GAT), .ZN(n463) );
  XNOR2_X1 U336 ( .A(n463), .B(KEYINPUT58), .ZN(n464) );
  XNOR2_X1 U337 ( .A(n465), .B(n464), .ZN(G1351GAT) );
  XOR2_X1 U338 ( .A(G64GAT), .B(KEYINPUT94), .Z(n293) );
  XNOR2_X1 U339 ( .A(G204GAT), .B(G92GAT), .ZN(n292) );
  XNOR2_X1 U340 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U341 ( .A(n337), .B(n294), .Z(n296) );
  NAND2_X1 U342 ( .A1(G226GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U343 ( .A(n296), .B(n295), .ZN(n298) );
  XNOR2_X1 U344 ( .A(G8GAT), .B(G211GAT), .ZN(n297) );
  XNOR2_X1 U345 ( .A(n297), .B(KEYINPUT78), .ZN(n327) );
  XOR2_X1 U346 ( .A(n298), .B(n327), .Z(n309) );
  XOR2_X1 U347 ( .A(KEYINPUT17), .B(KEYINPUT19), .Z(n300) );
  XNOR2_X1 U348 ( .A(KEYINPUT18), .B(KEYINPUT85), .ZN(n299) );
  XNOR2_X1 U349 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U350 ( .A(n301), .B(KEYINPUT86), .Z(n303) );
  XNOR2_X1 U351 ( .A(G190GAT), .B(G183GAT), .ZN(n302) );
  XNOR2_X1 U352 ( .A(n303), .B(n302), .ZN(n305) );
  XOR2_X1 U353 ( .A(G169GAT), .B(G176GAT), .Z(n304) );
  XOR2_X1 U354 ( .A(n305), .B(n304), .Z(n459) );
  XOR2_X1 U355 ( .A(KEYINPUT21), .B(KEYINPUT91), .Z(n307) );
  XNOR2_X1 U356 ( .A(G197GAT), .B(G218GAT), .ZN(n306) );
  XNOR2_X1 U357 ( .A(n307), .B(n306), .ZN(n427) );
  XNOR2_X1 U358 ( .A(n459), .B(n427), .ZN(n308) );
  XNOR2_X1 U359 ( .A(n309), .B(n308), .ZN(n526) );
  XNOR2_X1 U360 ( .A(G71GAT), .B(G57GAT), .ZN(n315) );
  INV_X1 U361 ( .A(KEYINPUT13), .ZN(n310) );
  NAND2_X1 U362 ( .A1(G64GAT), .A2(n310), .ZN(n313) );
  INV_X1 U363 ( .A(G64GAT), .ZN(n311) );
  NAND2_X1 U364 ( .A1(n311), .A2(KEYINPUT13), .ZN(n312) );
  NAND2_X1 U365 ( .A1(n313), .A2(n312), .ZN(n314) );
  XNOR2_X1 U366 ( .A(n315), .B(n314), .ZN(n366) );
  XOR2_X1 U367 ( .A(G15GAT), .B(G127GAT), .Z(n448) );
  XNOR2_X1 U368 ( .A(n366), .B(n448), .ZN(n319) );
  AND2_X1 U369 ( .A1(G231GAT), .A2(G233GAT), .ZN(n317) );
  INV_X1 U370 ( .A(KEYINPUT80), .ZN(n316) );
  XOR2_X1 U371 ( .A(KEYINPUT72), .B(G1GAT), .Z(n376) );
  XNOR2_X1 U372 ( .A(n376), .B(G183GAT), .ZN(n320) );
  XNOR2_X1 U373 ( .A(n321), .B(n320), .ZN(n325) );
  XOR2_X1 U374 ( .A(KEYINPUT79), .B(KEYINPUT12), .Z(n323) );
  XNOR2_X1 U375 ( .A(KEYINPUT15), .B(KEYINPUT14), .ZN(n322) );
  XNOR2_X1 U376 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U377 ( .A(n325), .B(n324), .Z(n329) );
  XOR2_X1 U378 ( .A(G22GAT), .B(G155GAT), .Z(n326) );
  XOR2_X1 U379 ( .A(G78GAT), .B(n326), .Z(n426) );
  XNOR2_X1 U380 ( .A(n426), .B(n327), .ZN(n328) );
  INV_X1 U381 ( .A(n587), .ZN(n563) );
  XNOR2_X1 U382 ( .A(KEYINPUT36), .B(KEYINPUT102), .ZN(n355) );
  XOR2_X1 U383 ( .A(KEYINPUT74), .B(KEYINPUT73), .Z(n331) );
  XNOR2_X1 U384 ( .A(G99GAT), .B(G92GAT), .ZN(n330) );
  XNOR2_X1 U385 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U386 ( .A(G85GAT), .B(n332), .Z(n370) );
  INV_X1 U387 ( .A(G162GAT), .ZN(n333) );
  NAND2_X1 U388 ( .A1(G50GAT), .A2(n333), .ZN(n336) );
  INV_X1 U389 ( .A(G50GAT), .ZN(n334) );
  NAND2_X1 U390 ( .A1(n334), .A2(G162GAT), .ZN(n335) );
  NAND2_X1 U391 ( .A1(n336), .A2(n335), .ZN(n436) );
  XNOR2_X1 U392 ( .A(n337), .B(n436), .ZN(n339) );
  AND2_X1 U393 ( .A1(G232GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U394 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U395 ( .A(G43GAT), .B(G134GAT), .Z(n453) );
  XNOR2_X1 U396 ( .A(n340), .B(n453), .ZN(n350) );
  XOR2_X1 U397 ( .A(KEYINPUT9), .B(KEYINPUT77), .Z(n342) );
  XNOR2_X1 U398 ( .A(G218GAT), .B(KEYINPUT65), .ZN(n341) );
  XNOR2_X1 U399 ( .A(n342), .B(n341), .ZN(n346) );
  XOR2_X1 U400 ( .A(KEYINPUT67), .B(KEYINPUT11), .Z(n344) );
  XNOR2_X1 U401 ( .A(KEYINPUT10), .B(KEYINPUT75), .ZN(n343) );
  XNOR2_X1 U402 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U403 ( .A(n346), .B(n345), .Z(n348) );
  INV_X1 U404 ( .A(G106GAT), .ZN(n347) );
  XNOR2_X1 U405 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n351) );
  XNOR2_X1 U406 ( .A(n351), .B(KEYINPUT7), .ZN(n379) );
  XNOR2_X1 U407 ( .A(n379), .B(G190GAT), .ZN(n352) );
  XNOR2_X1 U408 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U409 ( .A(n370), .B(n354), .ZN(n398) );
  XNOR2_X1 U410 ( .A(n355), .B(n398), .ZN(n592) );
  NOR2_X1 U411 ( .A1(n563), .A2(n592), .ZN(n358) );
  INV_X1 U412 ( .A(KEYINPUT66), .ZN(n356) );
  XNOR2_X1 U413 ( .A(n358), .B(n357), .ZN(n371) );
  XOR2_X1 U414 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n360) );
  XNOR2_X1 U415 ( .A(G120GAT), .B(KEYINPUT31), .ZN(n359) );
  XNOR2_X1 U416 ( .A(n360), .B(n359), .ZN(n364) );
  XOR2_X1 U417 ( .A(G78GAT), .B(G176GAT), .Z(n362) );
  NAND2_X1 U418 ( .A1(G230GAT), .A2(G233GAT), .ZN(n361) );
  XNOR2_X1 U419 ( .A(n362), .B(n361), .ZN(n363) );
  XOR2_X1 U420 ( .A(n364), .B(n363), .Z(n368) );
  XNOR2_X1 U421 ( .A(G106GAT), .B(G204GAT), .ZN(n365) );
  XNOR2_X1 U422 ( .A(n365), .B(G148GAT), .ZN(n432) );
  XNOR2_X1 U423 ( .A(n432), .B(n366), .ZN(n367) );
  XNOR2_X1 U424 ( .A(n368), .B(n367), .ZN(n369) );
  NOR2_X1 U425 ( .A1(n371), .A2(n582), .ZN(n372) );
  XNOR2_X1 U426 ( .A(n372), .B(KEYINPUT113), .ZN(n392) );
  XOR2_X1 U427 ( .A(G141GAT), .B(G197GAT), .Z(n374) );
  XNOR2_X1 U428 ( .A(G36GAT), .B(G22GAT), .ZN(n373) );
  XNOR2_X1 U429 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U430 ( .A(n375), .B(G43GAT), .Z(n378) );
  XNOR2_X1 U431 ( .A(n376), .B(G50GAT), .ZN(n377) );
  XNOR2_X1 U432 ( .A(n378), .B(n377), .ZN(n383) );
  XOR2_X1 U433 ( .A(n379), .B(KEYINPUT29), .Z(n381) );
  NAND2_X1 U434 ( .A1(G229GAT), .A2(G233GAT), .ZN(n380) );
  XNOR2_X1 U435 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U436 ( .A(n383), .B(n382), .Z(n391) );
  XOR2_X1 U437 ( .A(G8GAT), .B(G113GAT), .Z(n385) );
  XNOR2_X1 U438 ( .A(G169GAT), .B(G15GAT), .ZN(n384) );
  XNOR2_X1 U439 ( .A(n385), .B(n384), .ZN(n389) );
  XOR2_X1 U440 ( .A(KEYINPUT30), .B(KEYINPUT70), .Z(n387) );
  XNOR2_X1 U441 ( .A(KEYINPUT69), .B(KEYINPUT71), .ZN(n386) );
  XNOR2_X1 U442 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U443 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U444 ( .A(n391), .B(n390), .Z(n555) );
  INV_X1 U445 ( .A(n555), .ZN(n579) );
  NOR2_X1 U446 ( .A1(n392), .A2(n579), .ZN(n393) );
  XNOR2_X1 U447 ( .A(n393), .B(KEYINPUT114), .ZN(n403) );
  XNOR2_X1 U448 ( .A(KEYINPUT47), .B(KEYINPUT112), .ZN(n401) );
  XOR2_X1 U449 ( .A(KEYINPUT41), .B(n582), .Z(n558) );
  NAND2_X1 U450 ( .A1(n558), .A2(n579), .ZN(n395) );
  XNOR2_X1 U451 ( .A(n587), .B(KEYINPUT109), .ZN(n570) );
  NAND2_X1 U452 ( .A1(n396), .A2(n570), .ZN(n397) );
  XNOR2_X1 U453 ( .A(n397), .B(KEYINPUT111), .ZN(n399) );
  NAND2_X1 U454 ( .A1(n399), .A2(n398), .ZN(n400) );
  XNOR2_X1 U455 ( .A(n401), .B(n400), .ZN(n402) );
  NOR2_X1 U456 ( .A1(n403), .A2(n402), .ZN(n404) );
  XNOR2_X1 U457 ( .A(n404), .B(KEYINPUT48), .ZN(n552) );
  NOR2_X1 U458 ( .A1(n526), .A2(n552), .ZN(n405) );
  XNOR2_X1 U459 ( .A(n405), .B(KEYINPUT54), .ZN(n576) );
  XOR2_X1 U460 ( .A(G85GAT), .B(G148GAT), .Z(n407) );
  XNOR2_X1 U461 ( .A(G134GAT), .B(G155GAT), .ZN(n406) );
  XNOR2_X1 U462 ( .A(n407), .B(n406), .ZN(n409) );
  XOR2_X1 U463 ( .A(G29GAT), .B(G162GAT), .Z(n408) );
  XNOR2_X1 U464 ( .A(n409), .B(n408), .ZN(n423) );
  XOR2_X1 U465 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n411) );
  XNOR2_X1 U466 ( .A(KEYINPUT93), .B(KEYINPUT1), .ZN(n410) );
  XNOR2_X1 U467 ( .A(n411), .B(n410), .ZN(n415) );
  XOR2_X1 U468 ( .A(KEYINPUT6), .B(G57GAT), .Z(n413) );
  XNOR2_X1 U469 ( .A(G1GAT), .B(G127GAT), .ZN(n412) );
  XNOR2_X1 U470 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U471 ( .A(n415), .B(n414), .Z(n421) );
  XOR2_X1 U472 ( .A(G120GAT), .B(KEYINPUT81), .Z(n417) );
  XNOR2_X1 U473 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n416) );
  XNOR2_X1 U474 ( .A(n417), .B(n416), .ZN(n450) );
  XOR2_X1 U475 ( .A(KEYINPUT92), .B(KEYINPUT3), .Z(n419) );
  XNOR2_X1 U476 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n418) );
  XNOR2_X1 U477 ( .A(n419), .B(n418), .ZN(n431) );
  XNOR2_X1 U478 ( .A(n450), .B(n431), .ZN(n420) );
  XNOR2_X1 U479 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U480 ( .A(n423), .B(n422), .ZN(n425) );
  NAND2_X1 U481 ( .A1(G225GAT), .A2(G233GAT), .ZN(n424) );
  XNOR2_X1 U482 ( .A(n425), .B(n424), .ZN(n575) );
  XOR2_X1 U483 ( .A(n427), .B(n426), .Z(n440) );
  XOR2_X1 U484 ( .A(KEYINPUT90), .B(G211GAT), .Z(n429) );
  NAND2_X1 U485 ( .A1(G228GAT), .A2(G233GAT), .ZN(n428) );
  XNOR2_X1 U486 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U487 ( .A(n430), .B(KEYINPUT22), .Z(n434) );
  XNOR2_X1 U488 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U489 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U490 ( .A(n435), .B(KEYINPUT24), .Z(n438) );
  XNOR2_X1 U491 ( .A(n436), .B(KEYINPUT23), .ZN(n437) );
  XNOR2_X1 U492 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U493 ( .A(n440), .B(n439), .ZN(n482) );
  INV_X1 U494 ( .A(n482), .ZN(n441) );
  AND2_X1 U495 ( .A1(n575), .A2(n441), .ZN(n442) );
  XNOR2_X1 U496 ( .A(n443), .B(KEYINPUT55), .ZN(n461) );
  XOR2_X1 U497 ( .A(KEYINPUT20), .B(KEYINPUT83), .Z(n445) );
  XNOR2_X1 U498 ( .A(G71GAT), .B(KEYINPUT82), .ZN(n444) );
  XNOR2_X1 U499 ( .A(n445), .B(n444), .ZN(n458) );
  XOR2_X1 U500 ( .A(KEYINPUT88), .B(KEYINPUT87), .Z(n447) );
  XNOR2_X1 U501 ( .A(G99GAT), .B(KEYINPUT64), .ZN(n446) );
  XNOR2_X1 U502 ( .A(n447), .B(n446), .ZN(n449) );
  XOR2_X1 U503 ( .A(n449), .B(n448), .Z(n456) );
  XOR2_X1 U504 ( .A(n450), .B(KEYINPUT84), .Z(n452) );
  NAND2_X1 U505 ( .A1(G227GAT), .A2(G233GAT), .ZN(n451) );
  XNOR2_X1 U506 ( .A(n452), .B(n451), .ZN(n454) );
  XNOR2_X1 U507 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U508 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U509 ( .A(n458), .B(n457), .ZN(n460) );
  XOR2_X2 U510 ( .A(n460), .B(n459), .Z(n529) );
  NOR2_X1 U511 ( .A1(n461), .A2(n529), .ZN(n462) );
  XNOR2_X1 U512 ( .A(KEYINPUT121), .B(n462), .ZN(n466) );
  NOR2_X1 U513 ( .A1(n466), .A2(n398), .ZN(n465) );
  INV_X1 U514 ( .A(n466), .ZN(n569) );
  NAND2_X1 U515 ( .A1(n569), .A2(n558), .ZN(n470) );
  XOR2_X1 U516 ( .A(KEYINPUT122), .B(KEYINPUT57), .Z(n468) );
  XNOR2_X1 U517 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n467) );
  XNOR2_X1 U518 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U519 ( .A(n470), .B(n469), .ZN(G1349GAT) );
  XNOR2_X1 U520 ( .A(KEYINPUT34), .B(KEYINPUT99), .ZN(n490) );
  OR2_X1 U521 ( .A1(n555), .A2(n582), .ZN(n502) );
  NAND2_X1 U522 ( .A1(n398), .A2(n587), .ZN(n471) );
  XOR2_X1 U523 ( .A(KEYINPUT16), .B(n471), .Z(n487) );
  NOR2_X1 U524 ( .A1(n526), .A2(n529), .ZN(n472) );
  NOR2_X1 U525 ( .A1(n482), .A2(n472), .ZN(n473) );
  XOR2_X1 U526 ( .A(n473), .B(KEYINPUT25), .Z(n474) );
  XNOR2_X1 U527 ( .A(KEYINPUT96), .B(n474), .ZN(n477) );
  NAND2_X1 U528 ( .A1(n482), .A2(n529), .ZN(n475) );
  XNOR2_X1 U529 ( .A(n475), .B(KEYINPUT26), .ZN(n578) );
  XNOR2_X1 U530 ( .A(n526), .B(KEYINPUT27), .ZN(n480) );
  NOR2_X1 U531 ( .A1(n578), .A2(n480), .ZN(n476) );
  NOR2_X1 U532 ( .A1(n477), .A2(n476), .ZN(n478) );
  XNOR2_X1 U533 ( .A(n478), .B(KEYINPUT97), .ZN(n479) );
  NAND2_X1 U534 ( .A1(n479), .A2(n575), .ZN(n486) );
  NOR2_X1 U535 ( .A1(n575), .A2(n480), .ZN(n554) );
  XOR2_X1 U536 ( .A(KEYINPUT28), .B(KEYINPUT68), .Z(n481) );
  XNOR2_X1 U537 ( .A(n482), .B(n481), .ZN(n533) );
  NAND2_X1 U538 ( .A1(n554), .A2(n533), .ZN(n536) );
  XNOR2_X1 U539 ( .A(KEYINPUT95), .B(n536), .ZN(n484) );
  INV_X1 U540 ( .A(n529), .ZN(n538) );
  XNOR2_X1 U541 ( .A(KEYINPUT89), .B(n538), .ZN(n483) );
  NAND2_X1 U542 ( .A1(n484), .A2(n483), .ZN(n485) );
  NAND2_X1 U543 ( .A1(n486), .A2(n485), .ZN(n499) );
  NAND2_X1 U544 ( .A1(n487), .A2(n499), .ZN(n513) );
  NOR2_X1 U545 ( .A1(n502), .A2(n513), .ZN(n488) );
  XOR2_X1 U546 ( .A(KEYINPUT98), .B(n488), .Z(n497) );
  NOR2_X1 U547 ( .A1(n575), .A2(n497), .ZN(n489) );
  XNOR2_X1 U548 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U549 ( .A(G1GAT), .B(n491), .ZN(G1324GAT) );
  NOR2_X1 U550 ( .A1(n526), .A2(n497), .ZN(n492) );
  XOR2_X1 U551 ( .A(KEYINPUT100), .B(n492), .Z(n493) );
  XNOR2_X1 U552 ( .A(G8GAT), .B(n493), .ZN(G1325GAT) );
  NOR2_X1 U553 ( .A1(n497), .A2(n529), .ZN(n495) );
  XNOR2_X1 U554 ( .A(KEYINPUT101), .B(KEYINPUT35), .ZN(n494) );
  XNOR2_X1 U555 ( .A(n495), .B(n494), .ZN(n496) );
  XOR2_X1 U556 ( .A(G15GAT), .B(n496), .Z(G1326GAT) );
  NOR2_X1 U557 ( .A1(n533), .A2(n497), .ZN(n498) );
  XOR2_X1 U558 ( .A(G22GAT), .B(n498), .Z(G1327GAT) );
  NAND2_X1 U559 ( .A1(n563), .A2(n499), .ZN(n500) );
  NOR2_X1 U560 ( .A1(n500), .A2(n592), .ZN(n501) );
  XNOR2_X1 U561 ( .A(n501), .B(KEYINPUT37), .ZN(n524) );
  NOR2_X1 U562 ( .A1(n524), .A2(n502), .ZN(n503) );
  XOR2_X1 U563 ( .A(KEYINPUT38), .B(n503), .Z(n510) );
  NOR2_X1 U564 ( .A1(n575), .A2(n510), .ZN(n506) );
  XOR2_X1 U565 ( .A(G29GAT), .B(KEYINPUT103), .Z(n504) );
  XNOR2_X1 U566 ( .A(KEYINPUT39), .B(n504), .ZN(n505) );
  XNOR2_X1 U567 ( .A(n506), .B(n505), .ZN(G1328GAT) );
  NOR2_X1 U568 ( .A1(n526), .A2(n510), .ZN(n507) );
  XOR2_X1 U569 ( .A(G36GAT), .B(n507), .Z(G1329GAT) );
  NOR2_X1 U570 ( .A1(n510), .A2(n529), .ZN(n508) );
  XOR2_X1 U571 ( .A(KEYINPUT40), .B(n508), .Z(n509) );
  XNOR2_X1 U572 ( .A(G43GAT), .B(n509), .ZN(G1330GAT) );
  NOR2_X1 U573 ( .A1(n533), .A2(n510), .ZN(n511) );
  XOR2_X1 U574 ( .A(KEYINPUT104), .B(n511), .Z(n512) );
  XNOR2_X1 U575 ( .A(G50GAT), .B(n512), .ZN(G1331GAT) );
  NAND2_X1 U576 ( .A1(n558), .A2(n555), .ZN(n523) );
  NOR2_X1 U577 ( .A1(n523), .A2(n513), .ZN(n514) );
  XNOR2_X1 U578 ( .A(n514), .B(KEYINPUT105), .ZN(n520) );
  NOR2_X1 U579 ( .A1(n575), .A2(n520), .ZN(n515) );
  XOR2_X1 U580 ( .A(KEYINPUT42), .B(n515), .Z(n516) );
  XNOR2_X1 U581 ( .A(G57GAT), .B(n516), .ZN(G1332GAT) );
  NOR2_X1 U582 ( .A1(n526), .A2(n520), .ZN(n517) );
  XOR2_X1 U583 ( .A(G64GAT), .B(n517), .Z(G1333GAT) );
  NOR2_X1 U584 ( .A1(n529), .A2(n520), .ZN(n518) );
  XOR2_X1 U585 ( .A(KEYINPUT106), .B(n518), .Z(n519) );
  XNOR2_X1 U586 ( .A(G71GAT), .B(n519), .ZN(G1334GAT) );
  NOR2_X1 U587 ( .A1(n533), .A2(n520), .ZN(n522) );
  XNOR2_X1 U588 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n521) );
  XNOR2_X1 U589 ( .A(n522), .B(n521), .ZN(G1335GAT) );
  OR2_X1 U590 ( .A1(n524), .A2(n523), .ZN(n532) );
  NOR2_X1 U591 ( .A1(n575), .A2(n532), .ZN(n525) );
  XOR2_X1 U592 ( .A(G85GAT), .B(n525), .Z(G1336GAT) );
  NOR2_X1 U593 ( .A1(n526), .A2(n532), .ZN(n528) );
  XNOR2_X1 U594 ( .A(G92GAT), .B(KEYINPUT107), .ZN(n527) );
  XNOR2_X1 U595 ( .A(n528), .B(n527), .ZN(G1337GAT) );
  NOR2_X1 U596 ( .A1(n529), .A2(n532), .ZN(n530) );
  XOR2_X1 U597 ( .A(KEYINPUT108), .B(n530), .Z(n531) );
  XNOR2_X1 U598 ( .A(G99GAT), .B(n531), .ZN(G1338GAT) );
  NOR2_X1 U599 ( .A1(n533), .A2(n532), .ZN(n534) );
  XOR2_X1 U600 ( .A(KEYINPUT44), .B(n534), .Z(n535) );
  XNOR2_X1 U601 ( .A(G106GAT), .B(n535), .ZN(G1339GAT) );
  NOR2_X1 U602 ( .A1(n552), .A2(n536), .ZN(n537) );
  NAND2_X1 U603 ( .A1(n538), .A2(n537), .ZN(n539) );
  XOR2_X1 U604 ( .A(KEYINPUT115), .B(n539), .Z(n548) );
  INV_X1 U605 ( .A(n548), .ZN(n541) );
  NAND2_X1 U606 ( .A1(n579), .A2(n541), .ZN(n540) );
  XNOR2_X1 U607 ( .A(G113GAT), .B(n540), .ZN(G1340GAT) );
  XOR2_X1 U608 ( .A(G120GAT), .B(KEYINPUT49), .Z(n543) );
  NAND2_X1 U609 ( .A1(n541), .A2(n558), .ZN(n542) );
  XNOR2_X1 U610 ( .A(n543), .B(n542), .ZN(G1341GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n545) );
  XNOR2_X1 U612 ( .A(G127GAT), .B(KEYINPUT50), .ZN(n544) );
  XNOR2_X1 U613 ( .A(n545), .B(n544), .ZN(n547) );
  NOR2_X1 U614 ( .A1(n570), .A2(n548), .ZN(n546) );
  XOR2_X1 U615 ( .A(n547), .B(n546), .Z(G1342GAT) );
  NOR2_X1 U616 ( .A1(n398), .A2(n548), .ZN(n550) );
  XNOR2_X1 U617 ( .A(KEYINPUT118), .B(KEYINPUT51), .ZN(n549) );
  XNOR2_X1 U618 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U619 ( .A(G134GAT), .B(n551), .ZN(G1343GAT) );
  NOR2_X1 U620 ( .A1(n578), .A2(n552), .ZN(n553) );
  NAND2_X1 U621 ( .A1(n554), .A2(n553), .ZN(n566) );
  NOR2_X1 U622 ( .A1(n555), .A2(n566), .ZN(n557) );
  XNOR2_X1 U623 ( .A(G141GAT), .B(KEYINPUT119), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(G1344GAT) );
  INV_X1 U625 ( .A(n558), .ZN(n559) );
  NOR2_X1 U626 ( .A1(n559), .A2(n566), .ZN(n561) );
  XNOR2_X1 U627 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n560) );
  XNOR2_X1 U628 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U629 ( .A(G148GAT), .B(n562), .ZN(G1345GAT) );
  NOR2_X1 U630 ( .A1(n563), .A2(n566), .ZN(n564) );
  XOR2_X1 U631 ( .A(KEYINPUT120), .B(n564), .Z(n565) );
  XNOR2_X1 U632 ( .A(G155GAT), .B(n565), .ZN(G1346GAT) );
  NOR2_X1 U633 ( .A1(n398), .A2(n566), .ZN(n567) );
  XOR2_X1 U634 ( .A(G162GAT), .B(n567), .Z(G1347GAT) );
  NAND2_X1 U635 ( .A1(n579), .A2(n569), .ZN(n568) );
  XNOR2_X1 U636 ( .A(G169GAT), .B(n568), .ZN(G1348GAT) );
  NOR2_X1 U637 ( .A1(n570), .A2(n466), .ZN(n571) );
  XOR2_X1 U638 ( .A(G183GAT), .B(n571), .Z(G1350GAT) );
  XOR2_X1 U639 ( .A(KEYINPUT60), .B(KEYINPUT124), .Z(n573) );
  XNOR2_X1 U640 ( .A(G197GAT), .B(KEYINPUT123), .ZN(n572) );
  XNOR2_X1 U641 ( .A(n573), .B(n572), .ZN(n574) );
  XOR2_X1 U642 ( .A(KEYINPUT59), .B(n574), .Z(n581) );
  NAND2_X1 U643 ( .A1(n576), .A2(n575), .ZN(n577) );
  NOR2_X1 U644 ( .A1(n578), .A2(n577), .ZN(n590) );
  NAND2_X1 U645 ( .A1(n590), .A2(n579), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1352GAT) );
  XOR2_X1 U647 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n584) );
  NAND2_X1 U648 ( .A1(n590), .A2(n582), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(n586) );
  XOR2_X1 U650 ( .A(G204GAT), .B(KEYINPUT125), .Z(n585) );
  XNOR2_X1 U651 ( .A(n586), .B(n585), .ZN(G1353GAT) );
  XOR2_X1 U652 ( .A(G211GAT), .B(KEYINPUT127), .Z(n589) );
  NAND2_X1 U653 ( .A1(n590), .A2(n587), .ZN(n588) );
  XNOR2_X1 U654 ( .A(n589), .B(n588), .ZN(G1354GAT) );
  INV_X1 U655 ( .A(n590), .ZN(n591) );
  NOR2_X1 U656 ( .A1(n592), .A2(n591), .ZN(n593) );
  XOR2_X1 U657 ( .A(KEYINPUT62), .B(n593), .Z(n594) );
  XNOR2_X1 U658 ( .A(G218GAT), .B(n594), .ZN(G1355GAT) );
endmodule

