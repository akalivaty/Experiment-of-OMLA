//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 1 1 0 0 1 0 1 0 0 1 0 0 0 1 1 1 1 0 1 0 0 1 0 1 0 0 0 1 1 0 0 1 1 0 1 1 0 0 1 1 0 0 1 1 1 0 0 0 0 1 1 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:42 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n563, new_n564, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n610, new_n613, new_n614, new_n615, new_n616, new_n617, new_n619,
    new_n620, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1181, new_n1182, new_n1183, new_n1184;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT65), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n450), .A2(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n453), .B(new_n454), .ZN(new_n455));
  NAND4_X1  g030(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n455), .A2(new_n456), .ZN(G325));
  XOR2_X1   g032(.A(G325), .B(KEYINPUT68), .Z(G261));
  AOI22_X1  g033(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  OR2_X1    g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT69), .ZN(new_n461));
  NAND2_X1  g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(KEYINPUT69), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n463), .A2(new_n466), .A3(G125), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  INV_X1    g045(.A(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G101), .ZN(new_n473));
  INV_X1    g048(.A(G2105), .ZN(new_n474));
  OAI211_X1 g049(.A(G137), .B(new_n474), .C1(new_n464), .C2(new_n465), .ZN(new_n475));
  AND3_X1   g050(.A1(new_n470), .A2(new_n473), .A3(new_n475), .ZN(G160));
  NOR2_X1   g051(.A1(new_n464), .A2(new_n465), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n477), .A2(new_n474), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  OAI21_X1  g055(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(G112), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n481), .B1(new_n482), .B2(G2105), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT70), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n477), .A2(G2105), .ZN(new_n485));
  AOI211_X1 g060(.A(new_n480), .B(new_n484), .C1(G136), .C2(new_n485), .ZN(G162));
  NOR2_X1   g061(.A1(new_n474), .A2(G114), .ZN(new_n487));
  OAI21_X1  g062(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n488));
  OR2_X1    g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  OAI211_X1 g064(.A(G126), .B(G2105), .C1(new_n464), .C2(new_n465), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  OAI211_X1 g066(.A(G138), .B(new_n474), .C1(new_n464), .C2(new_n465), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n493));
  INV_X1    g068(.A(G138), .ZN(new_n494));
  NOR3_X1   g069(.A1(new_n494), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n463), .A2(new_n466), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n491), .B1(new_n493), .B2(new_n496), .ZN(G164));
  INV_X1    g072(.A(G543), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n498), .A2(KEYINPUT5), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT5), .ZN(new_n500));
  OAI21_X1  g075(.A(KEYINPUT71), .B1(new_n500), .B2(G543), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT71), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n502), .A2(new_n498), .A3(KEYINPUT5), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n499), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n504), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AND2_X1   g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  OAI21_X1  g084(.A(G543), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G50), .ZN(new_n512));
  XNOR2_X1  g087(.A(KEYINPUT6), .B(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n504), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G88), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n512), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n507), .A2(new_n516), .ZN(G166));
  NAND2_X1  g092(.A1(new_n510), .A2(KEYINPUT72), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT72), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n513), .A2(new_n519), .A3(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n521), .A2(G51), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n504), .A2(G63), .A3(G651), .ZN(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT7), .ZN(new_n525));
  INV_X1    g100(.A(G89), .ZN(new_n526));
  OAI211_X1 g101(.A(new_n523), .B(new_n525), .C1(new_n514), .C2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n522), .A2(new_n527), .ZN(G168));
  INV_X1    g103(.A(G52), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n529), .B1(new_n518), .B2(new_n520), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n501), .A2(new_n503), .ZN(new_n531));
  INV_X1    g106(.A(new_n499), .ZN(new_n532));
  AND4_X1   g107(.A1(G90), .A2(new_n531), .A3(new_n532), .A4(new_n513), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(G77), .A2(G543), .ZN(new_n535));
  INV_X1    g110(.A(new_n535), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n536), .B1(new_n504), .B2(G64), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT73), .ZN(new_n538));
  OAI21_X1  g113(.A(G651), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(G64), .ZN(new_n540));
  AOI211_X1 g115(.A(new_n540), .B(new_n499), .C1(new_n501), .C2(new_n503), .ZN(new_n541));
  NOR3_X1   g116(.A1(new_n541), .A2(KEYINPUT73), .A3(new_n536), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n534), .B1(new_n539), .B2(new_n542), .ZN(G301));
  INV_X1    g118(.A(G301), .ZN(G171));
  INV_X1    g119(.A(G43), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n545), .B1(new_n518), .B2(new_n520), .ZN(new_n546));
  AND2_X1   g121(.A1(KEYINPUT75), .A2(G81), .ZN(new_n547));
  NOR2_X1   g122(.A1(KEYINPUT75), .A2(G81), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  AND4_X1   g124(.A1(new_n531), .A2(new_n532), .A3(new_n513), .A4(new_n549), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n546), .A2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT74), .ZN(new_n552));
  AND2_X1   g127(.A1(G68), .A2(G543), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n553), .B1(new_n504), .B2(G56), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n552), .B1(new_n554), .B2(new_n506), .ZN(new_n555));
  INV_X1    g130(.A(G56), .ZN(new_n556));
  AOI211_X1 g131(.A(new_n556), .B(new_n499), .C1(new_n501), .C2(new_n503), .ZN(new_n557));
  OAI211_X1 g132(.A(KEYINPUT74), .B(G651), .C1(new_n557), .C2(new_n553), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n551), .A2(new_n555), .A3(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(G153));
  NAND4_X1  g136(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND4_X1  g139(.A1(G319), .A2(G483), .A3(G661), .A4(new_n564), .ZN(G188));
  INV_X1    g140(.A(new_n514), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G91), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n511), .A2(G53), .ZN(new_n568));
  AND2_X1   g143(.A1(KEYINPUT76), .A2(KEYINPUT9), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n568), .B(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(G78), .A2(G543), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT77), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n504), .B(new_n573), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n572), .B1(new_n574), .B2(G65), .ZN(new_n575));
  OAI211_X1 g150(.A(new_n567), .B(new_n570), .C1(new_n575), .C2(new_n506), .ZN(G299));
  INV_X1    g151(.A(G168), .ZN(G286));
  INV_X1    g152(.A(G166), .ZN(G303));
  NAND2_X1  g153(.A1(new_n566), .A2(G87), .ZN(new_n579));
  OAI21_X1  g154(.A(G651), .B1(new_n504), .B2(G74), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n511), .A2(G49), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(G288));
  AOI22_X1  g157(.A1(new_n504), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n583), .A2(new_n506), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n511), .A2(G48), .ZN(new_n585));
  INV_X1    g160(.A(G86), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n514), .B2(new_n586), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(G305));
  AOI22_X1  g164(.A1(new_n566), .A2(G85), .B1(new_n521), .B2(G47), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n504), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n506), .B2(new_n591), .ZN(G290));
  NOR2_X1   g167(.A1(new_n504), .A2(new_n573), .ZN(new_n593));
  AOI211_X1 g168(.A(KEYINPUT77), .B(new_n499), .C1(new_n501), .C2(new_n503), .ZN(new_n594));
  OAI21_X1  g169(.A(G66), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(G79), .A2(G543), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n506), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n504), .A2(G92), .A3(new_n513), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT10), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g175(.A1(new_n504), .A2(KEYINPUT10), .A3(G92), .A4(new_n513), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n521), .A2(G54), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n597), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n605), .B(KEYINPUT78), .ZN(new_n606));
  MUX2_X1   g181(.A(new_n606), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g182(.A(new_n606), .B(G301), .S(G868), .Z(G321));
  NAND2_X1  g183(.A1(G286), .A2(G868), .ZN(new_n609));
  INV_X1    g184(.A(G299), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(G868), .ZN(G297));
  OAI21_X1  g186(.A(new_n609), .B1(new_n610), .B2(G868), .ZN(G280));
  AOI22_X1  g187(.A1(new_n600), .A2(new_n601), .B1(G54), .B2(new_n521), .ZN(new_n613));
  AOI22_X1  g188(.A1(new_n574), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(new_n614), .B2(new_n506), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT78), .ZN(new_n616));
  XOR2_X1   g191(.A(KEYINPUT79), .B(G559), .Z(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(G860), .B2(new_n617), .ZN(G148));
  NAND2_X1  g193(.A1(new_n616), .A2(new_n617), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(G868), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(G868), .B2(new_n560), .ZN(G323));
  XNOR2_X1  g196(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g197(.A1(new_n485), .A2(G135), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(KEYINPUT81), .Z(new_n624));
  OAI21_X1  g199(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n625));
  INV_X1    g200(.A(G111), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n625), .B1(new_n626), .B2(G2105), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n627), .B1(new_n478), .B2(G123), .ZN(new_n628));
  AND2_X1   g203(.A1(new_n624), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2096), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n463), .A2(new_n466), .A3(new_n472), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT80), .B(KEYINPUT12), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n631), .B(new_n632), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT13), .ZN(new_n634));
  INV_X1    g209(.A(G2100), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n634), .A2(new_n635), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n630), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(KEYINPUT82), .Z(G156));
  INV_X1    g214(.A(KEYINPUT14), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2427), .B(G2438), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2430), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT15), .B(G2435), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n640), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n644), .B1(new_n643), .B2(new_n642), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2451), .B(G2454), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT16), .ZN(new_n647));
  XNOR2_X1  g222(.A(G1341), .B(G1348), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n645), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2443), .B(G2446), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n652), .A2(G14), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n650), .A2(new_n651), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n653), .A2(new_n654), .ZN(G401));
  XNOR2_X1  g230(.A(G2072), .B(G2078), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT83), .ZN(new_n657));
  XOR2_X1   g232(.A(KEYINPUT85), .B(KEYINPUT17), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2067), .B(G2678), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n660), .B(KEYINPUT84), .Z(new_n661));
  XOR2_X1   g236(.A(G2084), .B(G2090), .Z(new_n662));
  NAND3_X1  g237(.A1(new_n659), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT86), .ZN(new_n664));
  INV_X1    g239(.A(new_n657), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n662), .B1(new_n665), .B2(new_n661), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n666), .B1(new_n659), .B2(new_n661), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n657), .A2(new_n660), .A3(new_n662), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(KEYINPUT18), .Z(new_n669));
  NAND3_X1  g244(.A1(new_n664), .A2(new_n667), .A3(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G2096), .B(G2100), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(G227));
  XNOR2_X1  g247(.A(G1971), .B(G1976), .ZN(new_n673));
  INV_X1    g248(.A(KEYINPUT19), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G1956), .B(G2474), .Z(new_n676));
  XOR2_X1   g251(.A(G1961), .B(G1966), .Z(new_n677));
  AND2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(KEYINPUT20), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n676), .A2(new_n677), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  MUX2_X1   g258(.A(new_n683), .B(new_n682), .S(new_n675), .Z(new_n684));
  NOR2_X1   g259(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(G1991), .B(G1996), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1981), .B(G1986), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT87), .B(KEYINPUT88), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(G229));
  INV_X1    g268(.A(G16), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G23), .ZN(new_n695));
  INV_X1    g270(.A(G288), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n695), .B1(new_n696), .B2(new_n694), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT33), .B(G1976), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  NOR2_X1   g274(.A1(G6), .A2(G16), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(new_n588), .B2(G16), .ZN(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT32), .B(G1981), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n701), .B(new_n702), .Z(new_n703));
  NAND2_X1  g278(.A1(new_n694), .A2(G22), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(G166), .B2(new_n694), .ZN(new_n705));
  INV_X1    g280(.A(G1971), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n699), .A2(new_n703), .A3(new_n707), .ZN(new_n708));
  OR2_X1    g283(.A1(new_n708), .A2(KEYINPUT34), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n708), .A2(KEYINPUT34), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n485), .A2(G131), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n478), .A2(G119), .ZN(new_n712));
  OR2_X1    g287(.A1(G95), .A2(G2105), .ZN(new_n713));
  OAI211_X1 g288(.A(new_n713), .B(G2104), .C1(G107), .C2(new_n474), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n711), .A2(new_n712), .A3(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(G29), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n716), .A2(KEYINPUT89), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n716), .A2(KEYINPUT89), .ZN(new_n718));
  AND2_X1   g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(new_n720));
  MUX2_X1   g295(.A(G25), .B(new_n715), .S(new_n720), .Z(new_n721));
  XOR2_X1   g296(.A(KEYINPUT35), .B(G1991), .Z(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  NOR2_X1   g298(.A1(G16), .A2(G24), .ZN(new_n724));
  XNOR2_X1  g299(.A(G290), .B(KEYINPUT90), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n724), .B1(new_n725), .B2(G16), .ZN(new_n726));
  INV_X1    g301(.A(G1986), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NAND4_X1  g303(.A1(new_n709), .A2(new_n710), .A3(new_n723), .A4(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT36), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT31), .B(G11), .ZN(new_n732));
  INV_X1    g307(.A(G28), .ZN(new_n733));
  AOI21_X1  g308(.A(G29), .B1(new_n733), .B2(KEYINPUT30), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT97), .ZN(new_n735));
  OAI22_X1  g310(.A1(new_n734), .A2(new_n735), .B1(KEYINPUT30), .B2(new_n733), .ZN(new_n736));
  AND2_X1   g311(.A1(new_n734), .A2(new_n735), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n732), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(new_n629), .B2(new_n720), .ZN(new_n739));
  NOR2_X1   g314(.A1(G164), .A2(new_n719), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(G27), .B2(new_n719), .ZN(new_n741));
  INV_X1    g316(.A(G2078), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  AOI22_X1  g318(.A1(new_n485), .A2(G141), .B1(G105), .B2(new_n472), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n478), .A2(G129), .ZN(new_n745));
  NAND3_X1  g320(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT26), .Z(new_n747));
  AND3_X1   g322(.A1(new_n744), .A2(new_n745), .A3(new_n747), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n748), .A2(new_n716), .ZN(new_n749));
  AND2_X1   g324(.A1(new_n716), .A2(G32), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT27), .B(G1996), .ZN(new_n751));
  INV_X1    g326(.A(new_n751), .ZN(new_n752));
  OR3_X1    g327(.A1(new_n749), .A2(new_n750), .A3(new_n752), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n739), .A2(new_n743), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n719), .A2(G35), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G162), .B2(new_n719), .ZN(new_n756));
  XNOR2_X1  g331(.A(KEYINPUT29), .B(G2090), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n752), .B1(new_n749), .B2(new_n750), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n756), .A2(new_n757), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n741), .A2(new_n742), .ZN(new_n762));
  NOR4_X1   g337(.A1(new_n754), .A2(new_n760), .A3(new_n761), .A4(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n716), .A2(G33), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT93), .B(KEYINPUT25), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT94), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n474), .A2(G103), .A3(G2104), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n485), .A2(G139), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n770), .A2(KEYINPUT95), .ZN(new_n771));
  INV_X1    g346(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n770), .A2(KEYINPUT95), .ZN(new_n773));
  NAND3_X1  g348(.A1(new_n463), .A2(new_n466), .A3(G127), .ZN(new_n774));
  INV_X1    g349(.A(G115), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n774), .B1(new_n775), .B2(new_n471), .ZN(new_n776));
  AOI22_X1  g351(.A1(new_n772), .A2(new_n773), .B1(G2105), .B2(new_n776), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n764), .B1(new_n777), .B2(new_n716), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n778), .A2(G2072), .ZN(new_n779));
  INV_X1    g354(.A(KEYINPUT24), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n780), .A2(G34), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n719), .B1(new_n780), .B2(G34), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT96), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n781), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(new_n783), .B2(new_n782), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(G29), .B2(G160), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(G2084), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n694), .A2(G21), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G168), .B2(new_n694), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(G1966), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n787), .A2(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(G2072), .ZN(new_n792));
  OAI211_X1 g367(.A(new_n792), .B(new_n764), .C1(new_n777), .C2(new_n716), .ZN(new_n793));
  NAND4_X1  g368(.A1(new_n763), .A2(new_n779), .A3(new_n791), .A4(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n694), .A2(G20), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT23), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(new_n610), .B2(new_n694), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(G1956), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n694), .A2(G5), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G171), .B2(new_n694), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G1961), .ZN(new_n801));
  NOR3_X1   g376(.A1(new_n794), .A2(new_n798), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n694), .A2(G4), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(new_n616), .B2(new_n694), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n804), .A2(G1348), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n804), .A2(G1348), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n719), .A2(G26), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT91), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT28), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n808), .A2(new_n809), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n485), .A2(G140), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n478), .A2(G128), .ZN(new_n813));
  OR2_X1    g388(.A1(G104), .A2(G2105), .ZN(new_n814));
  OAI211_X1 g389(.A(new_n814), .B(G2104), .C1(G116), .C2(new_n474), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n812), .A2(new_n813), .A3(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(new_n816), .ZN(new_n817));
  OAI211_X1 g392(.A(new_n810), .B(new_n811), .C1(new_n716), .C2(new_n817), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(G2067), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n694), .A2(G19), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(new_n560), .B2(new_n694), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(G1341), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n805), .A2(new_n806), .A3(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT92), .ZN(new_n825));
  OR2_X1    g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n824), .A2(new_n825), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n802), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n731), .A2(new_n828), .ZN(G311));
  INV_X1    g404(.A(KEYINPUT98), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n830), .B1(new_n731), .B2(new_n828), .ZN(new_n831));
  AND2_X1   g406(.A1(new_n802), .A2(new_n827), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n729), .B(KEYINPUT36), .ZN(new_n833));
  NAND4_X1  g408(.A1(new_n832), .A2(new_n833), .A3(KEYINPUT98), .A4(new_n826), .ZN(new_n834));
  AND2_X1   g409(.A1(new_n831), .A2(new_n834), .ZN(G150));
  NAND2_X1  g410(.A1(new_n504), .A2(G67), .ZN(new_n836));
  NAND2_X1  g411(.A1(G80), .A2(G543), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n506), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(G55), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n839), .B1(new_n518), .B2(new_n520), .ZN(new_n840));
  AND3_X1   g415(.A1(new_n504), .A2(G93), .A3(new_n513), .ZN(new_n841));
  NOR3_X1   g416(.A1(new_n838), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n843), .A2(G860), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(KEYINPUT37), .Z(new_n845));
  XOR2_X1   g420(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n846));
  INV_X1    g421(.A(G559), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n846), .B1(new_n606), .B2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n846), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n616), .A2(G559), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n560), .A2(new_n842), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n843), .A2(new_n559), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n559), .B(new_n842), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n848), .A2(new_n856), .A3(new_n850), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n855), .A2(KEYINPUT39), .A3(new_n857), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n858), .B(KEYINPUT100), .Z(new_n859));
  INV_X1    g434(.A(KEYINPUT101), .ZN(new_n860));
  AOI21_X1  g435(.A(KEYINPUT39), .B1(new_n855), .B2(new_n857), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n861), .A2(G860), .ZN(new_n862));
  AND3_X1   g437(.A1(new_n859), .A2(new_n860), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n860), .B1(new_n859), .B2(new_n862), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n845), .B1(new_n863), .B2(new_n864), .ZN(G145));
  XNOR2_X1  g440(.A(new_n633), .B(new_n715), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n485), .A2(G142), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n478), .A2(G130), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n474), .A2(G118), .ZN(new_n869));
  OAI21_X1  g444(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n870));
  OAI211_X1 g445(.A(new_n867), .B(new_n868), .C1(new_n869), .C2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n866), .B(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n816), .B(G164), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n777), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n776), .A2(G2105), .ZN(new_n877));
  INV_X1    g452(.A(new_n773), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n877), .B1(new_n878), .B2(new_n771), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n879), .A2(new_n874), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n876), .A2(new_n748), .A3(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n748), .B1(new_n876), .B2(new_n880), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n873), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n883), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n885), .A2(new_n872), .A3(new_n881), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(G162), .B(G160), .ZN(new_n888));
  XOR2_X1   g463(.A(new_n888), .B(new_n629), .Z(new_n889));
  AOI21_X1  g464(.A(G37), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT102), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n886), .A2(new_n891), .ZN(new_n892));
  NAND4_X1  g467(.A1(new_n885), .A2(KEYINPUT102), .A3(new_n872), .A4(new_n881), .ZN(new_n893));
  INV_X1    g468(.A(new_n889), .ZN(new_n894));
  NAND4_X1  g469(.A1(new_n892), .A2(new_n893), .A3(new_n884), .A4(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n890), .A2(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g472(.A1(new_n619), .A2(new_n856), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n854), .B1(new_n616), .B2(new_n617), .ZN(new_n899));
  OAI21_X1  g474(.A(G65), .B1(new_n593), .B2(new_n594), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(new_n571), .ZN(new_n901));
  AOI22_X1  g476(.A1(new_n901), .A2(G651), .B1(G91), .B2(new_n566), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n615), .A2(new_n902), .A3(new_n570), .ZN(new_n903));
  NAND2_X1  g478(.A1(G299), .A2(new_n605), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  OR3_X1    g481(.A1(new_n898), .A2(new_n899), .A3(new_n906), .ZN(new_n907));
  AND3_X1   g482(.A1(new_n903), .A2(new_n904), .A3(KEYINPUT41), .ZN(new_n908));
  AOI21_X1  g483(.A(KEYINPUT41), .B1(new_n903), .B2(new_n904), .ZN(new_n909));
  OAI22_X1  g484(.A1(new_n898), .A2(new_n899), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(KEYINPUT104), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT103), .ZN(new_n913));
  XNOR2_X1  g488(.A(G288), .B(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(new_n588), .ZN(new_n915));
  XNOR2_X1  g490(.A(G288), .B(KEYINPUT103), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(G305), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(G303), .B(G290), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n915), .A2(new_n917), .A3(new_n919), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n923), .B(KEYINPUT42), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n912), .A2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT104), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n907), .A2(new_n926), .A3(new_n910), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n924), .B1(new_n912), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(G868), .B1(new_n925), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n929), .B1(G868), .B2(new_n842), .ZN(G295));
  OAI21_X1  g505(.A(new_n929), .B1(G868), .B2(new_n842), .ZN(G331));
  INV_X1    g506(.A(KEYINPUT105), .ZN(new_n932));
  OAI211_X1 g507(.A(new_n534), .B(new_n932), .C1(new_n539), .C2(new_n542), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(KEYINPUT73), .B1(new_n541), .B2(new_n536), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n504), .A2(G64), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n936), .A2(new_n538), .A3(new_n535), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n935), .A2(G651), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n932), .B1(new_n938), .B2(new_n534), .ZN(new_n939));
  NOR3_X1   g514(.A1(new_n934), .A2(new_n939), .A3(G168), .ZN(new_n940));
  NAND2_X1  g515(.A1(G301), .A2(KEYINPUT105), .ZN(new_n941));
  AOI21_X1  g516(.A(G286), .B1(new_n941), .B2(new_n933), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n854), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(G168), .B1(new_n934), .B2(new_n939), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n941), .A2(G286), .A3(new_n933), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n944), .A2(new_n856), .A3(new_n945), .ZN(new_n946));
  OAI211_X1 g521(.A(new_n943), .B(new_n946), .C1(new_n908), .C2(new_n909), .ZN(new_n947));
  AND3_X1   g522(.A1(new_n944), .A2(new_n856), .A3(new_n945), .ZN(new_n948));
  AOI22_X1  g523(.A1(new_n944), .A2(new_n945), .B1(new_n853), .B2(new_n852), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n905), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n947), .A2(new_n950), .ZN(new_n951));
  AND2_X1   g526(.A1(new_n921), .A2(new_n922), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(G37), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n923), .A2(new_n947), .A3(new_n950), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n956), .B(KEYINPUT43), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n957), .A2(KEYINPUT44), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n956), .A2(KEYINPUT106), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT107), .ZN(new_n960));
  AOI21_X1  g535(.A(G37), .B1(new_n951), .B2(new_n952), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT106), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n961), .A2(new_n962), .A3(new_n955), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n959), .A2(new_n960), .A3(KEYINPUT43), .A4(new_n963), .ZN(new_n964));
  AND3_X1   g539(.A1(new_n961), .A2(new_n962), .A3(new_n955), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n962), .B1(new_n961), .B2(new_n955), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT43), .ZN(new_n967));
  NOR3_X1   g542(.A1(new_n965), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n956), .A2(KEYINPUT43), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n969), .A2(KEYINPUT107), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n964), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n958), .B1(new_n971), .B2(KEYINPUT44), .ZN(G397));
  XNOR2_X1  g547(.A(KEYINPUT108), .B(G40), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n475), .A2(new_n473), .A3(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT109), .B1(new_n470), .B2(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n474), .B1(new_n467), .B2(new_n468), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT109), .ZN(new_n978));
  NOR3_X1   g553(.A1(new_n977), .A2(new_n974), .A3(new_n978), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n976), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT45), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n981), .B1(G164), .B2(G1384), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n748), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n983), .A2(G1996), .A3(new_n984), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n985), .B(KEYINPUT110), .ZN(new_n986));
  INV_X1    g561(.A(G2067), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n816), .B(new_n987), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n988), .B1(G1996), .B2(new_n984), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n986), .B1(new_n983), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(new_n722), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n715), .A2(new_n991), .ZN(new_n992));
  AND2_X1   g567(.A1(new_n715), .A2(new_n991), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n983), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n990), .A2(new_n994), .ZN(new_n995));
  XNOR2_X1  g570(.A(G290), .B(G1986), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n995), .B1(new_n983), .B2(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n496), .A2(new_n493), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n999), .A2(new_n490), .A3(new_n489), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT50), .ZN(new_n1001));
  INV_X1    g576(.A(G1384), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1000), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  OAI211_X1 g578(.A(new_n998), .B(new_n1003), .C1(new_n976), .C2(new_n979), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  OR2_X1    g580(.A1(new_n1005), .A2(G1961), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1000), .A2(KEYINPUT45), .A3(new_n1002), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(new_n982), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT53), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1010), .A2(G2078), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n1009), .A2(G40), .A3(G160), .A4(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(KEYINPUT111), .B1(new_n980), .B2(new_n1008), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n470), .A2(KEYINPUT109), .A3(new_n975), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n978), .B1(new_n977), .B2(new_n974), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT111), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n1016), .A2(new_n1017), .A3(new_n982), .A4(new_n1007), .ZN(new_n1018));
  AOI21_X1  g593(.A(G2078), .B1(new_n1013), .B2(new_n1018), .ZN(new_n1019));
  OAI211_X1 g594(.A(new_n1006), .B(new_n1012), .C1(new_n1019), .C2(KEYINPUT53), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT127), .ZN(new_n1021));
  AOI21_X1  g596(.A(G301), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  AND2_X1   g597(.A1(new_n1013), .A2(new_n1018), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1010), .B1(new_n1023), .B2(G2078), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1024), .A2(KEYINPUT127), .A3(new_n1006), .A4(new_n1012), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1022), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT54), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n980), .A2(new_n1008), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(new_n1011), .ZN(new_n1029));
  OAI211_X1 g604(.A(new_n1006), .B(new_n1029), .C1(new_n1019), .C2(KEYINPUT53), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1027), .B1(new_n1031), .B2(G301), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1026), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(G303), .A2(G8), .ZN(new_n1034));
  XNOR2_X1  g609(.A(new_n1034), .B(KEYINPUT55), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1013), .A2(new_n706), .A3(new_n1018), .ZN(new_n1036));
  OR2_X1    g611(.A1(KEYINPUT112), .A2(G2090), .ZN(new_n1037));
  NAND2_X1  g612(.A1(KEYINPUT112), .A2(G2090), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1005), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT115), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1036), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(G8), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1040), .B1(new_n1036), .B2(new_n1039), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1035), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(G8), .ZN(new_n1045));
  NOR2_X1   g620(.A1(G164), .A2(G1384), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1045), .B1(new_n1016), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n696), .A2(G1976), .ZN(new_n1048));
  INV_X1    g623(.A(G1976), .ZN(new_n1049));
  AOI21_X1  g624(.A(KEYINPUT52), .B1(G288), .B2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1047), .A2(new_n1048), .A3(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT113), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1052), .A2(KEYINPUT49), .ZN(new_n1053));
  OAI21_X1  g628(.A(G1981), .B1(new_n584), .B2(new_n587), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  NOR3_X1   g630(.A1(new_n584), .A2(new_n587), .A3(G1981), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1053), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1056), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1053), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1058), .A2(new_n1054), .A3(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1057), .A2(new_n1060), .A3(new_n1047), .ZN(new_n1061));
  AND2_X1   g636(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT52), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n1051), .B(new_n1061), .C1(new_n1062), .C2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1035), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1045), .B1(new_n1036), .B2(new_n1039), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1064), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  AND2_X1   g642(.A1(new_n1044), .A2(new_n1067), .ZN(new_n1068));
  AND2_X1   g643(.A1(new_n1030), .A2(G171), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1020), .A2(G171), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1027), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(KEYINPUT116), .B1(new_n1004), .B2(G2084), .ZN(new_n1072));
  AND2_X1   g647(.A1(new_n1003), .A2(new_n998), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT116), .ZN(new_n1074));
  INV_X1    g649(.A(G2084), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .A4(new_n1016), .ZN(new_n1076));
  INV_X1    g651(.A(G1966), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1077), .B1(new_n980), .B2(new_n1008), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1072), .A2(new_n1076), .A3(new_n1078), .ZN(new_n1079));
  AND2_X1   g654(.A1(new_n1079), .A2(G286), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1072), .A2(new_n1076), .A3(G168), .A4(new_n1078), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(G8), .ZN(new_n1082));
  OAI21_X1  g657(.A(KEYINPUT51), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1083));
  OR2_X1    g658(.A1(new_n1082), .A2(KEYINPUT51), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1033), .A2(new_n1068), .A3(new_n1071), .A4(new_n1085), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n616), .A2(KEYINPUT60), .ZN(new_n1087));
  OR2_X1    g662(.A1(new_n1005), .A2(G1348), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1016), .A2(new_n987), .A3(new_n1046), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT122), .ZN(new_n1090));
  OR2_X1    g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1088), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1093), .A2(KEYINPUT60), .A3(new_n616), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n616), .A2(KEYINPUT60), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1095), .A2(new_n1092), .A3(new_n1091), .A4(new_n1088), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1087), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT125), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(KEYINPUT59), .ZN(new_n1099));
  XOR2_X1   g674(.A(new_n1099), .B(KEYINPUT126), .Z(new_n1100));
  INV_X1    g675(.A(new_n1100), .ZN(new_n1101));
  XOR2_X1   g676(.A(KEYINPUT123), .B(G1996), .Z(new_n1102));
  NAND2_X1  g677(.A1(new_n1016), .A2(new_n1046), .ZN(new_n1103));
  XOR2_X1   g678(.A(KEYINPUT58), .B(G1341), .Z(new_n1104));
  AOI22_X1  g679(.A1(new_n1028), .A2(new_n1102), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  AND2_X1   g680(.A1(new_n1105), .A2(KEYINPUT124), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n560), .B1(new_n1105), .B2(KEYINPUT124), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1098), .A2(KEYINPUT59), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1101), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  OAI221_X1 g685(.A(new_n1100), .B1(new_n1098), .B2(KEYINPUT59), .C1(new_n1106), .C2(new_n1107), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1097), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT61), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n610), .A2(KEYINPUT57), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT119), .ZN(new_n1115));
  XNOR2_X1  g690(.A(new_n570), .B(new_n1115), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n567), .B1(new_n575), .B2(new_n506), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT120), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n902), .A2(KEYINPUT120), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1116), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  XNOR2_X1  g696(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1122), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1114), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT121), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  OAI211_X1 g701(.A(KEYINPUT121), .B(new_n1114), .C1(new_n1121), .C2(new_n1123), .ZN(new_n1127));
  XNOR2_X1  g702(.A(KEYINPUT56), .B(G2072), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1028), .A2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1129), .B1(new_n1005), .B2(G1956), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1126), .A2(new_n1127), .A3(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1130), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1113), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1130), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1137), .A2(KEYINPUT61), .A3(new_n1131), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1112), .A2(new_n1134), .A3(new_n1138), .ZN(new_n1139));
  AND2_X1   g714(.A1(new_n1093), .A2(new_n616), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1132), .B1(new_n1137), .B2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1086), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1085), .A2(KEYINPUT62), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT62), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1083), .A2(new_n1084), .A3(new_n1144), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1143), .A2(new_n1068), .A3(new_n1069), .A4(new_n1145), .ZN(new_n1146));
  AND3_X1   g721(.A1(new_n1079), .A2(G8), .A3(G168), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1044), .A2(new_n1067), .A3(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT63), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  AND2_X1   g725(.A1(new_n1147), .A2(KEYINPUT63), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT117), .ZN(new_n1152));
  AND2_X1   g727(.A1(new_n1066), .A2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1035), .B1(new_n1066), .B2(new_n1152), .ZN(new_n1154));
  OAI211_X1 g729(.A(new_n1151), .B(new_n1067), .C1(new_n1153), .C2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1150), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1066), .A2(new_n1065), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1157), .A2(new_n1064), .ZN(new_n1158));
  AND2_X1   g733(.A1(new_n1057), .A2(new_n1060), .ZN(new_n1159));
  NOR2_X1   g734(.A1(G288), .A2(G1976), .ZN(new_n1160));
  XOR2_X1   g735(.A(new_n1160), .B(KEYINPUT114), .Z(new_n1161));
  OAI21_X1  g736(.A(new_n1058), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1158), .B1(new_n1047), .B2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1146), .A2(new_n1156), .A3(new_n1163), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n997), .B1(new_n1142), .B2(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(new_n983), .ZN(new_n1166));
  OR3_X1    g741(.A1(new_n1166), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1167));
  OAI21_X1  g742(.A(KEYINPUT46), .B1(new_n1166), .B2(G1996), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n988), .A2(new_n748), .ZN(new_n1169));
  AOI22_X1  g744(.A1(new_n1167), .A2(new_n1168), .B1(new_n983), .B2(new_n1169), .ZN(new_n1170));
  XNOR2_X1  g745(.A(new_n1170), .B(KEYINPUT47), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n990), .A2(new_n992), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n817), .A2(new_n987), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1166), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(new_n995), .ZN(new_n1175));
  NOR3_X1   g750(.A1(new_n1166), .A2(G1986), .A3(G290), .ZN(new_n1176));
  XOR2_X1   g751(.A(new_n1176), .B(KEYINPUT48), .Z(new_n1177));
  AOI211_X1 g752(.A(new_n1171), .B(new_n1174), .C1(new_n1175), .C2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1165), .A2(new_n1178), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g754(.A(G229), .ZN(new_n1181));
  OAI21_X1  g755(.A(G319), .B1(new_n653), .B2(new_n654), .ZN(new_n1182));
  OR2_X1    g756(.A1(G227), .A2(new_n1182), .ZN(new_n1183));
  INV_X1    g757(.A(new_n1183), .ZN(new_n1184));
  AND4_X1   g758(.A1(new_n1181), .A2(new_n896), .A3(new_n957), .A4(new_n1184), .ZN(G308));
  NAND4_X1  g759(.A1(new_n1181), .A2(new_n896), .A3(new_n957), .A4(new_n1184), .ZN(G225));
endmodule


