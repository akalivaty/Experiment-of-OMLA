//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 0 0 0 0 0 0 1 0 0 0 0 1 1 0 1 0 1 0 1 0 0 1 1 0 0 1 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 0 1 1 1 0 0 1 0 1 0 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:30 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1295, new_n1296, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G250), .ZN(new_n205));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(G257), .ZN(new_n212));
  INV_X1    g0012(.A(G264), .ZN(new_n213));
  AOI211_X1 g0013(.A(new_n205), .B(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n207), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n202), .A2(G50), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(new_n214), .A2(KEYINPUT0), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n219), .B1(KEYINPUT0), .B2(new_n214), .ZN(new_n220));
  XOR2_X1   g0020(.A(new_n220), .B(KEYINPUT64), .Z(new_n221));
  XOR2_X1   g0021(.A(KEYINPUT65), .B(G244), .Z(new_n222));
  INV_X1    g0022(.A(G77), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G107), .A2(G264), .ZN(new_n228));
  NAND4_X1  g0028(.A1(new_n225), .A2(new_n226), .A3(new_n227), .A4(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n209), .B1(new_n224), .B2(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT1), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n221), .A2(new_n231), .ZN(G361));
  XOR2_X1   g0032(.A(G238), .B(G244), .Z(new_n233));
  XNOR2_X1  g0033(.A(G226), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XOR2_X1   g0042(.A(G107), .B(G116), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  AND2_X1   g0048(.A1(KEYINPUT3), .A2(G33), .ZN(new_n249));
  NOR2_X1   g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT67), .ZN(new_n251));
  NOR3_X1   g0051(.A1(new_n249), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT3), .ZN(new_n253));
  INV_X1    g0053(.A(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  AOI21_X1  g0056(.A(KEYINPUT67), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n252), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G1698), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n258), .A2(G222), .A3(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n258), .A2(G223), .A3(G1698), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n251), .B1(new_n249), .B2(new_n250), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n255), .A2(KEYINPUT67), .A3(new_n256), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G77), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n260), .A2(new_n261), .A3(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n215), .ZN(new_n267));
  NAND2_X1  g0067(.A1(G33), .A2(G41), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n266), .A2(new_n270), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n269), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n275), .B1(new_n267), .B2(new_n268), .ZN(new_n276));
  INV_X1    g0076(.A(new_n272), .ZN(new_n277));
  AOI22_X1  g0077(.A1(new_n274), .A2(G226), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n271), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G200), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n271), .A2(G190), .A3(new_n278), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT9), .ZN(new_n282));
  NAND3_X1  g0082(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(new_n215), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(KEYINPUT68), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT68), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n283), .A2(new_n286), .A3(new_n215), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  XNOR2_X1  g0088(.A(KEYINPUT8), .B(G58), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n207), .A2(G33), .ZN(new_n290));
  INV_X1    g0090(.A(G150), .ZN(new_n291));
  NOR2_X1   g0091(.A1(G20), .A2(G33), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  OAI22_X1  g0093(.A1(new_n289), .A2(new_n290), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G50), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n207), .B1(new_n201), .B2(new_n295), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n288), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(KEYINPUT69), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n288), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n295), .B1(new_n206), .B2(G20), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n298), .A2(new_n303), .ZN(new_n304));
  OAI22_X1  g0104(.A1(new_n297), .A2(KEYINPUT69), .B1(G50), .B2(new_n299), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n282), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n304), .ZN(new_n307));
  INV_X1    g0107(.A(new_n305), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n307), .A2(KEYINPUT9), .A3(new_n308), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n280), .A2(new_n281), .A3(new_n306), .A4(new_n309), .ZN(new_n310));
  XNOR2_X1  g0110(.A(new_n310), .B(KEYINPUT10), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n307), .A2(new_n308), .ZN(new_n312));
  INV_X1    g0112(.A(new_n279), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n312), .B1(new_n313), .B2(G169), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n279), .A2(G179), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n311), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n262), .A2(new_n263), .A3(G232), .A4(G1698), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(KEYINPUT70), .ZN(new_n321));
  NAND2_X1  g0121(.A1(G33), .A2(G97), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n262), .A2(new_n263), .A3(G226), .A4(new_n259), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n321), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n320), .A2(KEYINPUT70), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n270), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n269), .A2(new_n277), .A3(G274), .ZN(new_n327));
  INV_X1    g0127(.A(G238), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n327), .B1(new_n273), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n326), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(KEYINPUT13), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT13), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n326), .A2(new_n333), .A3(new_n330), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n332), .A2(G190), .A3(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT70), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n258), .A2(new_n336), .A3(G232), .A4(G1698), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n337), .A2(new_n321), .A3(new_n322), .A4(new_n323), .ZN(new_n338));
  AOI211_X1 g0138(.A(KEYINPUT13), .B(new_n329), .C1(new_n338), .C2(new_n270), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n333), .B1(new_n326), .B2(new_n330), .ZN(new_n340));
  OAI21_X1  g0140(.A(G200), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n207), .A2(G68), .ZN(new_n342));
  INV_X1    g0142(.A(G13), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n343), .A2(G1), .ZN(new_n344));
  NAND2_X1  g0144(.A1(KEYINPUT71), .A2(KEYINPUT12), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n342), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  NOR2_X1   g0146(.A1(KEYINPUT71), .A2(KEYINPUT12), .ZN(new_n347));
  XOR2_X1   g0147(.A(new_n346), .B(new_n347), .Z(new_n348));
  AOI21_X1  g0148(.A(new_n342), .B1(G50), .B2(new_n292), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n349), .B1(new_n223), .B2(new_n290), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n350), .A2(KEYINPUT11), .A3(new_n288), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n299), .A2(new_n215), .A3(new_n283), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n353), .B(G68), .C1(G1), .C2(new_n207), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n348), .A2(new_n351), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(KEYINPUT11), .B1(new_n350), .B2(new_n288), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n335), .A2(new_n341), .A3(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n339), .A2(new_n340), .ZN(new_n360));
  INV_X1    g0160(.A(G169), .ZN(new_n361));
  OAI21_X1  g0161(.A(KEYINPUT14), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT14), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n363), .B(G169), .C1(new_n339), .C2(new_n340), .ZN(new_n364));
  AOI21_X1  g0164(.A(KEYINPUT72), .B1(new_n360), .B2(G179), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT72), .ZN(new_n366));
  INV_X1    g0166(.A(G179), .ZN(new_n367));
  NOR4_X1   g0167(.A1(new_n339), .A2(new_n340), .A3(new_n366), .A4(new_n367), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n362), .B(new_n364), .C1(new_n365), .C2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n357), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n359), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n284), .ZN(new_n372));
  INV_X1    g0172(.A(G58), .ZN(new_n373));
  INV_X1    g0173(.A(G68), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(G20), .B1(new_n375), .B2(new_n201), .ZN(new_n376));
  INV_X1    g0176(.A(G159), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n376), .B1(new_n377), .B2(new_n293), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT7), .ZN(new_n379));
  XNOR2_X1  g0179(.A(KEYINPUT3), .B(G33), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n379), .B1(new_n380), .B2(G20), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n249), .A2(new_n250), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n382), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n378), .B1(new_n384), .B2(G68), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n372), .B1(new_n385), .B2(KEYINPUT16), .ZN(new_n386));
  AOI21_X1  g0186(.A(G20), .B1(new_n262), .B2(new_n263), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n383), .B1(new_n387), .B2(KEYINPUT7), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n378), .B1(new_n388), .B2(G68), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n386), .B1(KEYINPUT16), .B2(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n289), .B1(new_n206), .B2(G20), .ZN(new_n391));
  AOI22_X1  g0191(.A1(new_n301), .A2(new_n391), .B1(new_n300), .B2(new_n289), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  OR2_X1    g0193(.A1(G223), .A2(G1698), .ZN(new_n394));
  OAI221_X1 g0194(.A(new_n394), .B1(G226), .B2(new_n259), .C1(new_n249), .C2(new_n250), .ZN(new_n395));
  NAND2_X1  g0195(.A1(G33), .A2(G87), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n269), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(G232), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n327), .B1(new_n273), .B2(new_n398), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(G179), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n401), .B1(new_n361), .B2(new_n400), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n393), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(KEYINPUT18), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT18), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n393), .A2(new_n405), .A3(new_n402), .ZN(new_n406));
  INV_X1    g0206(.A(G200), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n400), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(G190), .ZN(new_n409));
  NOR3_X1   g0209(.A1(new_n397), .A2(new_n399), .A3(new_n409), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n390), .A2(new_n411), .A3(new_n392), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT17), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n392), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT16), .ZN(new_n416));
  INV_X1    g0216(.A(new_n383), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n207), .B1(new_n252), .B2(new_n257), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n417), .B1(new_n418), .B2(new_n379), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n419), .A2(new_n374), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n416), .B1(new_n420), .B2(new_n378), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n415), .B1(new_n421), .B2(new_n386), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n422), .A2(KEYINPUT17), .A3(new_n411), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n404), .A2(new_n406), .A3(new_n414), .A4(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n327), .B1(new_n273), .B2(new_n222), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n258), .A2(G232), .A3(new_n259), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n258), .A2(G238), .A3(G1698), .ZN(new_n428));
  INV_X1    g0228(.A(G107), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n427), .B(new_n428), .C1(new_n429), .C2(new_n258), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n426), .B1(new_n430), .B2(new_n270), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  OAI22_X1  g0232(.A1(new_n289), .A2(new_n293), .B1(new_n207), .B2(new_n223), .ZN(new_n433));
  XNOR2_X1  g0233(.A(KEYINPUT15), .B(G87), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n434), .A2(new_n290), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n284), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n223), .B1(new_n206), .B2(G20), .ZN(new_n437));
  AOI22_X1  g0237(.A1(new_n353), .A2(new_n437), .B1(new_n223), .B2(new_n300), .ZN(new_n438));
  AOI22_X1  g0238(.A1(new_n432), .A2(new_n361), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n431), .A2(new_n367), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n436), .A2(new_n438), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n442), .B1(new_n431), .B2(G190), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n443), .B1(new_n407), .B2(new_n431), .ZN(new_n444));
  AND2_X1   g0244(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n319), .A2(new_n371), .A3(new_n425), .A4(new_n445), .ZN(new_n446));
  NAND3_X1  g0246(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(new_n207), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT75), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n447), .A2(KEYINPUT75), .A3(new_n207), .ZN(new_n451));
  INV_X1    g0251(.A(G87), .ZN(new_n452));
  INV_X1    g0252(.A(G97), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n452), .A2(new_n453), .A3(new_n429), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n450), .A2(new_n451), .A3(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n380), .A2(new_n207), .A3(G68), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT19), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n457), .B1(new_n290), .B2(new_n453), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n455), .A2(new_n456), .A3(new_n458), .ZN(new_n459));
  AOI22_X1  g0259(.A1(new_n459), .A2(new_n284), .B1(new_n300), .B2(new_n434), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n206), .A2(G33), .ZN(new_n461));
  AND4_X1   g0261(.A1(new_n285), .A2(new_n287), .A3(new_n299), .A4(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n434), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(G244), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(G1698), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n466), .B1(G238), .B2(G1698), .ZN(new_n467));
  INV_X1    g0267(.A(G116), .ZN(new_n468));
  OAI22_X1  g0268(.A1(new_n467), .A2(new_n382), .B1(new_n254), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(new_n270), .ZN(new_n470));
  INV_X1    g0270(.A(G45), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n205), .B1(new_n471), .B2(G1), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n206), .A2(new_n275), .A3(G45), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n269), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  AND2_X1   g0274(.A1(new_n470), .A2(new_n474), .ZN(new_n475));
  AOI22_X1  g0275(.A1(new_n460), .A2(new_n464), .B1(new_n475), .B2(new_n367), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n470), .A2(new_n474), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(new_n361), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n407), .B1(new_n470), .B2(new_n474), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n254), .A2(new_n468), .ZN(new_n480));
  NOR2_X1   g0280(.A1(G238), .A2(G1698), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n481), .B1(new_n465), .B2(G1698), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n480), .B1(new_n482), .B2(new_n380), .ZN(new_n483));
  OAI211_X1 g0283(.A(G190), .B(new_n474), .C1(new_n483), .C2(new_n269), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT76), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n470), .A2(KEYINPUT76), .A3(G190), .A4(new_n474), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n479), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n459), .A2(new_n284), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n434), .A2(new_n300), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n462), .A2(G87), .ZN(new_n491));
  AND3_X1   g0291(.A1(new_n489), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  AOI22_X1  g0292(.A1(new_n476), .A2(new_n478), .B1(new_n488), .B2(new_n492), .ZN(new_n493));
  XNOR2_X1  g0293(.A(G97), .B(G107), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT6), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NOR3_X1   g0296(.A1(new_n495), .A2(new_n453), .A3(G107), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  AOI22_X1  g0299(.A1(new_n499), .A2(G20), .B1(G77), .B2(new_n292), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n500), .B1(new_n419), .B2(new_n429), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(new_n284), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n299), .A2(G97), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n503), .B1(new_n462), .B2(G97), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n262), .A2(new_n263), .A3(G250), .A4(G1698), .ZN(new_n505));
  NAND2_X1  g0305(.A1(G33), .A2(G283), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n465), .A2(G1698), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n508), .B1(new_n249), .B2(new_n250), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT4), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n507), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n510), .A2(new_n465), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n262), .A2(new_n263), .A3(new_n259), .A4(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n505), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n270), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT5), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(KEYINPUT74), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT74), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(KEYINPUT5), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(G41), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n516), .A2(G41), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n523), .A2(KEYINPUT73), .A3(new_n206), .A4(G45), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n206), .B(G45), .C1(new_n521), .C2(KEYINPUT5), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT73), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n522), .A2(new_n276), .A3(new_n524), .A4(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(G41), .B1(new_n517), .B2(new_n519), .ZN(new_n529));
  OAI211_X1 g0329(.A(G257), .B(new_n269), .C1(new_n529), .C2(new_n525), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  AND3_X1   g0332(.A1(new_n515), .A2(new_n409), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g0333(.A(G200), .B1(new_n515), .B2(new_n532), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n502), .B(new_n504), .C1(new_n533), .C2(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n497), .B1(new_n495), .B2(new_n494), .ZN(new_n536));
  OAI22_X1  g0336(.A1(new_n536), .A2(new_n207), .B1(new_n223), .B2(new_n293), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n537), .B1(new_n388), .B2(G107), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n504), .B1(new_n538), .B2(new_n372), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n515), .A2(new_n532), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n361), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n531), .B1(new_n270), .B2(new_n514), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n367), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n539), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n493), .A2(new_n535), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(KEYINPUT77), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT77), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n493), .A2(new_n535), .A3(new_n544), .A4(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n213), .A2(G1698), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n380), .B(new_n549), .C1(G257), .C2(G1698), .ZN(new_n550));
  INV_X1    g0350(.A(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(G303), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n552), .B1(new_n262), .B2(new_n263), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n270), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  OAI211_X1 g0354(.A(G270), .B(new_n269), .C1(new_n529), .C2(new_n525), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n554), .A2(new_n528), .A3(new_n555), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n506), .B(new_n207), .C1(G33), .C2(new_n453), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n468), .A2(G20), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n557), .A2(new_n284), .A3(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT20), .ZN(new_n560));
  XNOR2_X1  g0360(.A(new_n559), .B(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT78), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n461), .A2(G116), .ZN(new_n563));
  OR3_X1    g0363(.A1(new_n352), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n562), .B1(new_n352), .B2(new_n563), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n300), .A2(new_n468), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n561), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n556), .A2(new_n568), .A3(KEYINPUT21), .A4(G169), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n264), .A2(G303), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n269), .B1(new_n570), .B2(new_n550), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n528), .A2(new_n555), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n573), .A2(new_n568), .A3(G179), .ZN(new_n574));
  AND2_X1   g0374(.A1(new_n569), .A2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT79), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT21), .ZN(new_n577));
  INV_X1    g0377(.A(new_n568), .ZN(new_n578));
  OAI21_X1  g0378(.A(G169), .B1(new_n571), .B2(new_n572), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n577), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  OAI21_X1  g0380(.A(G200), .B1(new_n571), .B2(new_n572), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n554), .A2(G190), .A3(new_n528), .A4(new_n555), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n578), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n575), .A2(new_n576), .A3(new_n580), .A4(new_n583), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n580), .A2(new_n583), .A3(new_n574), .A4(new_n569), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(KEYINPUT79), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n546), .A2(new_n548), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n480), .A2(new_n207), .ZN(new_n588));
  OR3_X1    g0388(.A1(new_n207), .A2(KEYINPUT23), .A3(G107), .ZN(new_n589));
  NAND2_X1  g0389(.A1(KEYINPUT82), .A2(KEYINPUT24), .ZN(new_n590));
  OAI21_X1  g0390(.A(KEYINPUT23), .B1(new_n207), .B2(G107), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n588), .A2(new_n589), .A3(new_n590), .A4(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n207), .B(G87), .C1(new_n249), .C2(new_n250), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT80), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n380), .A2(KEYINPUT80), .A3(new_n207), .A4(G87), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n596), .A2(new_n597), .A3(KEYINPUT22), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT81), .ZN(new_n599));
  NOR3_X1   g0399(.A1(new_n452), .A2(KEYINPUT22), .A3(G20), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n262), .A2(new_n263), .A3(new_n600), .ZN(new_n601));
  AND3_X1   g0401(.A1(new_n598), .A2(new_n599), .A3(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n599), .B1(new_n598), .B2(new_n601), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n593), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NOR2_X1   g0404(.A1(KEYINPUT82), .A2(KEYINPUT24), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n593), .B(new_n605), .C1(new_n602), .C2(new_n603), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n372), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n300), .A2(new_n429), .ZN(new_n610));
  XNOR2_X1  g0410(.A(new_n610), .B(KEYINPUT25), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n611), .B1(G107), .B2(new_n462), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  OAI211_X1 g0414(.A(G264), .B(new_n269), .C1(new_n529), .C2(new_n525), .ZN(new_n615));
  NOR2_X1   g0415(.A1(G250), .A2(G1698), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n616), .B1(new_n212), .B2(G1698), .ZN(new_n617));
  XNOR2_X1  g0417(.A(KEYINPUT83), .B(G294), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n617), .A2(new_n380), .B1(new_n618), .B2(G33), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n528), .B(new_n615), .C1(new_n619), .C2(new_n269), .ZN(new_n620));
  AND2_X1   g0420(.A1(new_n620), .A2(KEYINPUT84), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n620), .A2(KEYINPUT84), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g0423(.A(KEYINPUT86), .B1(new_n623), .B2(G190), .ZN(new_n624));
  XNOR2_X1  g0424(.A(new_n620), .B(KEYINPUT84), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT86), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n625), .A2(new_n626), .A3(new_n409), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n620), .A2(new_n407), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n624), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n614), .A2(new_n629), .ZN(new_n630));
  OAI22_X1  g0430(.A1(new_n625), .A2(new_n361), .B1(new_n367), .B2(new_n620), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n631), .B1(new_n609), .B2(new_n613), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT85), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  OAI211_X1 g0434(.A(KEYINPUT85), .B(new_n631), .C1(new_n609), .C2(new_n613), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n587), .A2(new_n630), .A3(new_n634), .A4(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n446), .A2(new_n636), .ZN(G372));
  AND3_X1   g0437(.A1(new_n393), .A2(new_n405), .A3(new_n402), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n405), .B1(new_n393), .B2(new_n402), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g0440(.A(new_n412), .B(KEYINPUT17), .ZN(new_n641));
  INV_X1    g0441(.A(new_n441), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n369), .A2(new_n370), .B1(new_n358), .B2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT89), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n641), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n369), .A2(new_n370), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n642), .A2(new_n358), .ZN(new_n647));
  AND3_X1   g0447(.A1(new_n646), .A2(new_n644), .A3(new_n647), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n640), .B1(new_n645), .B2(new_n648), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n316), .B1(new_n649), .B2(new_n311), .ZN(new_n650));
  INV_X1    g0450(.A(new_n446), .ZN(new_n651));
  INV_X1    g0451(.A(new_n544), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n493), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(KEYINPUT26), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n474), .A2(KEYINPUT87), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n474), .A2(KEYINPUT87), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n470), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(new_n361), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n476), .A2(new_n658), .ZN(new_n659));
  AOI22_X1  g0459(.A1(new_n486), .A2(new_n487), .B1(new_n657), .B2(G200), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(new_n492), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT88), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n544), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT26), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n539), .A2(new_n541), .A3(new_n543), .A4(KEYINPUT88), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n662), .A2(new_n664), .A3(new_n665), .A4(new_n666), .ZN(new_n667));
  AND3_X1   g0467(.A1(new_n654), .A2(new_n667), .A3(new_n659), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n575), .A2(new_n580), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n632), .A2(new_n669), .ZN(new_n670));
  AND3_X1   g0470(.A1(new_n662), .A2(new_n544), .A3(new_n535), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n670), .A2(new_n630), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n651), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n650), .A2(new_n674), .ZN(G369));
  AND3_X1   g0475(.A1(new_n634), .A2(new_n630), .A3(new_n635), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n344), .A2(new_n207), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n678));
  XOR2_X1   g0478(.A(new_n678), .B(KEYINPUT90), .Z(new_n679));
  INV_X1    g0479(.A(G213), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n680), .B1(new_n677), .B2(KEYINPUT27), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(G343), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n676), .B1(new_n614), .B2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n632), .ZN(new_n686));
  INV_X1    g0486(.A(new_n684), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n586), .A2(new_n584), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n687), .A2(new_n568), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n669), .A2(new_n691), .ZN(new_n693));
  OAI21_X1  g0493(.A(G330), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n689), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n686), .A2(new_n684), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n669), .A2(new_n687), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n676), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n696), .A2(new_n697), .A3(new_n699), .ZN(G399));
  NOR2_X1   g0500(.A1(new_n211), .A2(G41), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n454), .A2(G116), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n702), .A2(G1), .A3(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(new_n217), .B2(new_n702), .ZN(new_n705));
  XNOR2_X1  g0505(.A(new_n705), .B(KEYINPUT28), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n687), .B1(new_n668), .B2(new_n672), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(KEYINPUT29), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n634), .A2(new_n635), .A3(new_n669), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(KEYINPUT93), .ZN(new_n710));
  AND2_X1   g0510(.A1(new_n630), .A2(new_n671), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT93), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n634), .A2(new_n712), .A3(new_n635), .A4(new_n669), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n710), .A2(new_n711), .A3(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n659), .B1(new_n653), .B2(KEYINPUT26), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n662), .A2(new_n664), .A3(new_n666), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n715), .B1(KEYINPUT26), .B2(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n687), .B1(new_n714), .B2(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n708), .B1(new_n718), .B2(KEYINPUT29), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n598), .A2(new_n601), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(KEYINPUT81), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n598), .A2(new_n599), .A3(new_n601), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n605), .B1(new_n723), .B2(new_n593), .ZN(new_n724));
  INV_X1    g0524(.A(new_n608), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n284), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(new_n612), .ZN(new_n727));
  AOI21_X1  g0527(.A(KEYINPUT85), .B1(new_n727), .B2(new_n631), .ZN(new_n728));
  INV_X1    g0528(.A(new_n635), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n730), .A2(new_n630), .A3(new_n587), .A4(new_n684), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n615), .B1(new_n619), .B2(new_n269), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n477), .A2(new_n732), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n542), .A2(new_n573), .A3(new_n733), .A4(G179), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT30), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n657), .A2(new_n620), .A3(new_n367), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(new_n573), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(new_n540), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n736), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n556), .A2(new_n367), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n741), .A2(KEYINPUT30), .A3(new_n542), .A4(new_n733), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(KEYINPUT92), .B1(new_n740), .B2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT31), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT92), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n736), .A2(new_n739), .A3(new_n742), .A4(new_n746), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n744), .A2(new_n745), .A3(new_n687), .A4(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n743), .B1(new_n740), .B2(KEYINPUT91), .ZN(new_n749));
  AOI22_X1  g0549(.A1(new_n735), .A2(new_n734), .B1(new_n738), .B2(new_n540), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT91), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n684), .B1(new_n749), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n748), .B1(new_n753), .B2(new_n745), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n731), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(G330), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n719), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n706), .B1(new_n758), .B2(G1), .ZN(new_n759));
  XNOR2_X1  g0559(.A(new_n759), .B(KEYINPUT94), .ZN(G364));
  XOR2_X1   g0560(.A(new_n694), .B(KEYINPUT96), .Z(new_n761));
  NOR2_X1   g0561(.A1(new_n343), .A2(G20), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n206), .B1(new_n762), .B2(G45), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n701), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AND2_X1   g0566(.A1(new_n761), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NOR3_X1   g0568(.A1(new_n692), .A2(G330), .A3(new_n693), .ZN(new_n769));
  XNOR2_X1  g0569(.A(new_n769), .B(KEYINPUT95), .ZN(new_n770));
  NOR2_X1   g0570(.A1(G13), .A2(G33), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(G20), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR3_X1   g0574(.A1(new_n692), .A2(new_n693), .A3(new_n774), .ZN(new_n775));
  NOR3_X1   g0575(.A1(new_n409), .A2(G179), .A3(G200), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(new_n207), .ZN(new_n777));
  INV_X1    g0577(.A(new_n618), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n207), .A2(new_n367), .ZN(new_n779));
  NOR2_X1   g0579(.A1(G190), .A2(G200), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(G311), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n777), .A2(new_n778), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n779), .A2(G200), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(new_n409), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n783), .B1(G326), .B2(new_n785), .ZN(new_n786));
  XOR2_X1   g0586(.A(new_n786), .B(KEYINPUT98), .Z(new_n787));
  NOR2_X1   g0587(.A1(new_n207), .A2(G179), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(new_n780), .ZN(new_n789));
  OR2_X1    g0589(.A1(new_n789), .A2(KEYINPUT99), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n789), .A2(KEYINPUT99), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(G329), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n779), .A2(G190), .A3(new_n407), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n258), .B1(G322), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n784), .A2(G190), .ZN(new_n798));
  INV_X1    g0598(.A(G317), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(KEYINPUT33), .ZN(new_n800));
  OR2_X1    g0600(.A1(new_n799), .A2(KEYINPUT33), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n798), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n788), .A2(G190), .A3(G200), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n788), .A2(new_n409), .A3(G200), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n804), .A2(G303), .B1(new_n806), .B2(G283), .ZN(new_n807));
  NAND4_X1  g0607(.A1(new_n794), .A2(new_n797), .A3(new_n802), .A4(new_n807), .ZN(new_n808));
  AOI22_X1  g0608(.A1(G50), .A2(new_n785), .B1(new_n798), .B2(G68), .ZN(new_n809));
  INV_X1    g0609(.A(new_n777), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(G97), .ZN(new_n811));
  INV_X1    g0611(.A(new_n789), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(G159), .ZN(new_n813));
  OAI211_X1 g0613(.A(new_n809), .B(new_n811), .C1(KEYINPUT32), .C2(new_n813), .ZN(new_n814));
  OAI22_X1  g0614(.A1(new_n795), .A2(new_n373), .B1(new_n781), .B2(new_n223), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n815), .B(KEYINPUT97), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n264), .B1(G87), .B2(new_n804), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n813), .A2(KEYINPUT32), .B1(G107), .B2(new_n806), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n816), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  OAI22_X1  g0619(.A1(new_n787), .A2(new_n808), .B1(new_n814), .B2(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n215), .B1(G20), .B2(new_n361), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n773), .A2(new_n821), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n211), .A2(new_n380), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n824), .B1(G45), .B2(new_n217), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n825), .B1(G45), .B2(new_n247), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n258), .A2(new_n210), .ZN(new_n827));
  INV_X1    g0627(.A(G355), .ZN(new_n828));
  OAI22_X1  g0628(.A1(new_n827), .A2(new_n828), .B1(G116), .B2(new_n210), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n823), .B1(new_n826), .B2(new_n829), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n822), .A2(new_n765), .A3(new_n830), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n768), .A2(new_n770), .B1(new_n775), .B2(new_n831), .ZN(G396));
  NAND2_X1  g0632(.A1(new_n673), .A2(new_n684), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n687), .A2(new_n442), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n444), .A2(new_n834), .B1(new_n439), .B2(new_n440), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n439), .A2(new_n440), .A3(new_n684), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n833), .A2(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(KEYINPUT103), .B1(new_n835), .B2(new_n837), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n444), .A2(new_n834), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(new_n441), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT103), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n843), .A2(new_n844), .A3(new_n836), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n841), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n840), .B1(new_n833), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(new_n757), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n848), .B(KEYINPUT104), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n849), .B(new_n766), .C1(new_n757), .C2(new_n847), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n821), .A2(new_n771), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n765), .B1(G77), .B2(new_n852), .ZN(new_n853));
  XNOR2_X1  g0653(.A(new_n853), .B(KEYINPUT100), .ZN(new_n854));
  INV_X1    g0654(.A(new_n821), .ZN(new_n855));
  INV_X1    g0655(.A(new_n798), .ZN(new_n856));
  XOR2_X1   g0656(.A(KEYINPUT101), .B(G283), .Z(new_n857));
  INV_X1    g0657(.A(new_n785), .ZN(new_n858));
  OAI22_X1  g0658(.A1(new_n856), .A2(new_n857), .B1(new_n858), .B2(new_n552), .ZN(new_n859));
  INV_X1    g0659(.A(new_n781), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n796), .A2(G294), .B1(new_n860), .B2(G116), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n861), .B(new_n811), .C1(new_n792), .C2(new_n782), .ZN(new_n862));
  AOI211_X1 g0662(.A(new_n859), .B(new_n862), .C1(G87), .C2(new_n806), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n264), .B1(new_n429), .B2(new_n803), .ZN(new_n864));
  XOR2_X1   g0664(.A(new_n864), .B(KEYINPUT102), .Z(new_n865));
  AOI22_X1  g0665(.A1(new_n796), .A2(G143), .B1(new_n860), .B2(G159), .ZN(new_n866));
  INV_X1    g0666(.A(G137), .ZN(new_n867));
  OAI221_X1 g0667(.A(new_n866), .B1(new_n858), .B2(new_n867), .C1(new_n291), .C2(new_n856), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT34), .ZN(new_n869));
  OR2_X1    g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  AOI22_X1  g0670(.A1(new_n810), .A2(G58), .B1(new_n804), .B2(G50), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n382), .B1(new_n806), .B2(G68), .ZN(new_n872));
  INV_X1    g0672(.A(G132), .ZN(new_n873));
  OAI211_X1 g0673(.A(new_n871), .B(new_n872), .C1(new_n792), .C2(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n874), .B1(new_n868), .B2(new_n869), .ZN(new_n875));
  AOI22_X1  g0675(.A1(new_n863), .A2(new_n865), .B1(new_n870), .B2(new_n875), .ZN(new_n876));
  OAI221_X1 g0676(.A(new_n854), .B1(new_n855), .B2(new_n876), .C1(new_n838), .C2(new_n772), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n850), .A2(new_n877), .ZN(G384));
  NOR2_X1   g0678(.A1(new_n762), .A2(new_n206), .ZN(new_n879));
  INV_X1    g0679(.A(G330), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n385), .A2(KEYINPUT16), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n374), .B1(new_n381), .B2(new_n383), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n416), .B1(new_n882), .B2(new_n378), .ZN(new_n883));
  AND3_X1   g0683(.A1(new_n881), .A2(new_n288), .A3(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n884), .A2(new_n415), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n885), .A2(new_n682), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n424), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT37), .ZN(new_n888));
  OAI22_X1  g0688(.A1(new_n884), .A2(new_n415), .B1(new_n402), .B2(new_n683), .ZN(new_n889));
  AOI211_X1 g0689(.A(KEYINPUT107), .B(new_n888), .C1(new_n889), .C2(new_n412), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n889), .A2(new_n412), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(KEYINPUT37), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n393), .A2(new_n683), .ZN(new_n894));
  NAND4_X1  g0694(.A1(new_n403), .A2(new_n894), .A3(new_n888), .A4(new_n412), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n893), .A2(new_n895), .A3(KEYINPUT107), .ZN(new_n896));
  NAND4_X1  g0696(.A1(new_n887), .A2(new_n891), .A3(KEYINPUT38), .A4(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n890), .B1(new_n424), .B2(new_n886), .ZN(new_n899));
  AOI21_X1  g0699(.A(KEYINPUT38), .B1(new_n899), .B2(new_n896), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n684), .A2(new_n357), .ZN(new_n902));
  XNOR2_X1  g0702(.A(new_n902), .B(KEYINPUT105), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n646), .A2(new_n358), .A3(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n332), .A2(G179), .A3(new_n334), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(new_n366), .ZN(new_n907));
  NAND4_X1  g0707(.A1(new_n332), .A2(KEYINPUT72), .A3(new_n334), .A4(G179), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n909), .A2(new_n362), .A3(new_n358), .A4(new_n364), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n902), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n905), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n745), .A2(KEYINPUT109), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n747), .A2(new_n687), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n746), .B1(new_n750), .B2(new_n742), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n913), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(new_n913), .ZN(new_n917));
  NAND4_X1  g0717(.A1(new_n744), .A2(new_n687), .A3(new_n747), .A4(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n919), .B1(new_n636), .B2(new_n687), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n912), .A2(new_n920), .A3(new_n838), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT110), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n901), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n839), .B1(new_n905), .B2(new_n911), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n924), .A2(KEYINPUT110), .A3(new_n920), .ZN(new_n925));
  AOI21_X1  g0725(.A(KEYINPUT40), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT40), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT38), .ZN(new_n928));
  INV_X1    g0728(.A(new_n402), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n412), .B1(new_n422), .B2(new_n929), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n422), .A2(new_n682), .ZN(new_n931));
  OAI21_X1  g0731(.A(KEYINPUT37), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  AND2_X1   g0732(.A1(new_n932), .A2(new_n895), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n894), .B1(new_n640), .B2(new_n641), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n928), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n927), .B1(new_n935), .B2(new_n897), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n924), .A2(new_n936), .A3(new_n920), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n926), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n546), .A2(new_n548), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(new_n690), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n634), .A2(new_n630), .A3(new_n635), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  AOI22_X1  g0743(.A1(new_n943), .A2(new_n684), .B1(new_n916), .B2(new_n918), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n944), .A2(new_n446), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n880), .B1(new_n939), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n939), .B2(new_n945), .ZN(new_n947));
  XOR2_X1   g0747(.A(new_n947), .B(KEYINPUT111), .Z(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n836), .B1(new_n833), .B2(new_n835), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(new_n912), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(KEYINPUT106), .ZN(new_n952));
  OR2_X1    g0752(.A1(new_n898), .A2(new_n900), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT106), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n950), .A2(new_n954), .A3(new_n912), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n952), .A2(new_n953), .A3(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n682), .B1(new_n638), .B2(new_n639), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT108), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n953), .A2(new_n958), .A3(KEYINPUT39), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT39), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n935), .A2(new_n960), .A3(new_n897), .ZN(new_n961));
  OAI211_X1 g0761(.A(KEYINPUT108), .B(new_n961), .C1(new_n901), .C2(new_n960), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n369), .A2(new_n370), .A3(new_n684), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n959), .A2(new_n962), .A3(new_n964), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n956), .A2(new_n957), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n714), .A2(new_n717), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n967), .A2(KEYINPUT29), .A3(new_n684), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n708), .A2(new_n446), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n650), .A2(new_n970), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n966), .B(new_n971), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n879), .B1(new_n949), .B2(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(new_n949), .B2(new_n972), .ZN(new_n974));
  OR2_X1    g0774(.A1(new_n499), .A2(KEYINPUT35), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n499), .A2(KEYINPUT35), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n975), .A2(G116), .A3(new_n216), .A4(new_n976), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT36), .ZN(new_n978));
  NOR3_X1   g0778(.A1(new_n217), .A2(new_n223), .A3(new_n375), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n374), .A2(G50), .ZN(new_n980));
  OAI211_X1 g0780(.A(G1), .B(new_n343), .C1(new_n979), .C2(new_n980), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n974), .A2(new_n978), .A3(new_n981), .ZN(G367));
  INV_X1    g0782(.A(new_n539), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n535), .B(new_n544), .C1(new_n983), .C2(new_n684), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n652), .A2(new_n687), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n676), .A2(new_n698), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(KEYINPUT42), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n544), .B1(new_n730), .B2(new_n984), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(new_n684), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n991), .A2(KEYINPUT112), .B1(KEYINPUT42), .B2(new_n987), .ZN(new_n992));
  AND2_X1   g0792(.A1(new_n991), .A2(KEYINPUT112), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n684), .A2(new_n492), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n995), .A2(new_n476), .A3(new_n658), .ZN(new_n996));
  INV_X1    g0796(.A(new_n662), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n996), .B1(new_n997), .B2(new_n995), .ZN(new_n998));
  INV_X1    g0798(.A(new_n986), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n696), .A2(new_n999), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n994), .A2(new_n998), .B1(KEYINPUT114), .B2(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n998), .B(KEYINPUT43), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT113), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1003), .B1(new_n994), .B2(new_n1004), .ZN(new_n1005));
  OAI211_X1 g0805(.A(KEYINPUT113), .B(new_n1002), .C1(new_n992), .C2(new_n993), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1001), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1007), .B1(KEYINPUT114), .B2(new_n1000), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n1000), .A2(KEYINPUT114), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n1001), .A2(new_n1005), .A3(new_n1009), .A4(new_n1006), .ZN(new_n1010));
  XOR2_X1   g0810(.A(new_n701), .B(KEYINPUT41), .Z(new_n1011));
  OAI211_X1 g0811(.A(new_n685), .B(new_n688), .C1(new_n669), .C2(new_n687), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(new_n699), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n761), .A2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1012), .A2(new_n695), .A3(new_n699), .ZN(new_n1015));
  AND3_X1   g0815(.A1(new_n758), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n699), .A2(new_n697), .A3(new_n986), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT45), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1017), .B(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n699), .A2(new_n697), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT44), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n986), .B1(KEYINPUT115), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n1021), .A2(KEYINPUT115), .ZN(new_n1024));
  OR2_X1    g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n1019), .A2(new_n1025), .A3(new_n696), .A4(new_n1026), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1019), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n696), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1016), .A2(new_n1027), .A3(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1011), .B1(new_n1031), .B2(new_n758), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1008), .B(new_n1010), .C1(new_n1032), .C2(new_n764), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n823), .B1(new_n210), .B2(new_n434), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(new_n824), .B2(new_n240), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n766), .A2(new_n1035), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n796), .A2(G150), .B1(new_n812), .B2(G137), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n295), .B2(new_n781), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n805), .A2(new_n223), .ZN(new_n1039));
  NOR3_X1   g0839(.A1(new_n1038), .A2(new_n264), .A3(new_n1039), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n777), .A2(new_n374), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(G159), .B2(new_n798), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n785), .A2(G143), .B1(new_n804), .B2(G58), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1040), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n798), .A2(new_n618), .B1(new_n806), .B2(G97), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1045), .B1(new_n429), .B2(new_n777), .C1(new_n782), .C2(new_n858), .ZN(new_n1046));
  AOI21_X1  g0846(.A(KEYINPUT46), .B1(new_n804), .B2(G116), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n795), .A2(new_n552), .B1(new_n789), .B2(new_n799), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n382), .B1(new_n857), .B2(new_n781), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT46), .ZN(new_n1050));
  NOR3_X1   g0850(.A1(new_n803), .A2(new_n1050), .A3(new_n468), .ZN(new_n1051));
  OR4_X1    g0851(.A1(new_n1047), .A2(new_n1048), .A3(new_n1049), .A4(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1044), .B1(new_n1046), .B2(new_n1052), .ZN(new_n1053));
  XOR2_X1   g0853(.A(new_n1053), .B(KEYINPUT47), .Z(new_n1054));
  OAI221_X1 g0854(.A(new_n1036), .B1(new_n998), .B2(new_n774), .C1(new_n1054), .C2(new_n855), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1033), .A2(new_n1055), .ZN(G387));
  AND2_X1   g0856(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n1057), .A2(new_n758), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1016), .A2(new_n702), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1058), .B1(new_n1059), .B2(KEYINPUT117), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT117), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1061), .B1(new_n1016), .B2(new_n702), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1057), .A2(new_n764), .ZN(new_n1064));
  AND2_X1   g0864(.A1(new_n237), .A2(G45), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n824), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n1065), .A2(new_n1066), .B1(new_n703), .B2(new_n827), .ZN(new_n1067));
  OR3_X1    g0867(.A1(new_n289), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1068));
  OAI21_X1  g0868(.A(KEYINPUT50), .B1(new_n289), .B2(G50), .ZN(new_n1069));
  AOI21_X1  g0869(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1070));
  NAND4_X1  g0870(.A1(new_n1068), .A2(new_n703), .A3(new_n1069), .A4(new_n1070), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n1067), .A2(new_n1071), .B1(new_n429), .B2(new_n211), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n823), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n765), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n781), .A2(new_n374), .B1(new_n789), .B2(new_n291), .ZN(new_n1075));
  AOI211_X1 g0875(.A(new_n382), .B(new_n1075), .C1(G50), .C2(new_n796), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n804), .A2(G77), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n289), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n463), .A2(new_n810), .B1(new_n798), .B2(new_n1078), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n785), .A2(G159), .B1(new_n806), .B2(G97), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n1076), .A2(new_n1077), .A3(new_n1079), .A4(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n380), .B1(new_n812), .B2(G326), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n777), .A2(new_n857), .B1(new_n778), .B2(new_n803), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n796), .A2(G317), .B1(new_n860), .B2(G303), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n785), .A2(G322), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1084), .B(new_n1085), .C1(new_n782), .C2(new_n856), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT48), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1083), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n1087), .B2(new_n1086), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT49), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n1082), .B1(new_n468), .B2(new_n805), .C1(new_n1089), .C2(new_n1090), .ZN(new_n1091));
  AND2_X1   g0891(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1081), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(KEYINPUT116), .ZN(new_n1094));
  OR2_X1    g0894(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n855), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1074), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1097), .B1(new_n689), .B2(new_n774), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1064), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1063), .A2(new_n1100), .ZN(G393));
  NAND2_X1  g0901(.A1(new_n1030), .A2(new_n1027), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n1102), .A2(new_n763), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n999), .A2(new_n773), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n823), .B1(new_n453), .B2(new_n210), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(new_n824), .B2(new_n244), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n858), .A2(new_n799), .B1(new_n782), .B2(new_n795), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(new_n1107), .B(KEYINPUT52), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(G294), .A2(new_n860), .B1(new_n812), .B2(G322), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n856), .A2(new_n552), .B1(new_n805), .B2(new_n429), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n777), .A2(new_n468), .B1(new_n857), .B2(new_n803), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n1108), .A2(new_n264), .A3(new_n1109), .A4(new_n1112), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n777), .A2(new_n223), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(new_n1078), .B2(new_n860), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1115), .B1(new_n295), .B2(new_n856), .ZN(new_n1116));
  INV_X1    g0916(.A(KEYINPUT119), .ZN(new_n1117));
  OR2_X1    g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n858), .A2(new_n291), .B1(new_n377), .B2(new_n795), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n1119), .B(KEYINPUT51), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1118), .A2(new_n1120), .A3(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n382), .B1(new_n812), .B2(G143), .ZN(new_n1123));
  OAI221_X1 g0923(.A(new_n1123), .B1(new_n374), .B2(new_n803), .C1(new_n452), .C2(new_n805), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1124), .B(KEYINPUT118), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1113), .B1(new_n1122), .B2(new_n1125), .ZN(new_n1126));
  AOI211_X1 g0926(.A(new_n766), .B(new_n1106), .C1(new_n1126), .C2(new_n821), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1103), .B1(new_n1104), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1057), .A2(new_n758), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1102), .A2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1130), .A2(new_n701), .A3(new_n1031), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1128), .A2(new_n1131), .ZN(G390));
  NAND2_X1  g0932(.A1(new_n959), .A2(new_n962), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n951), .A2(new_n963), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n964), .B1(new_n935), .B2(new_n897), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n837), .B1(new_n718), .B2(new_n843), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n912), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1136), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n912), .A2(new_n755), .A3(G330), .A4(new_n838), .ZN(new_n1140));
  AND3_X1   g0940(.A1(new_n1135), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n880), .B1(new_n731), .B2(new_n919), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n924), .A2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(new_n1135), .B2(new_n1139), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1141), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(new_n764), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n765), .B1(new_n1078), .B2(new_n852), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n805), .A2(new_n295), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n856), .A2(new_n867), .B1(new_n377), .B2(new_n777), .ZN(new_n1149));
  AOI211_X1 g0949(.A(new_n1148), .B(new_n1149), .C1(G128), .C2(new_n785), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n803), .A2(new_n291), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1151), .B(KEYINPUT53), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n793), .A2(G125), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(KEYINPUT54), .B(G143), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n795), .A2(new_n873), .B1(new_n781), .B2(new_n1154), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1155), .A2(new_n264), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1150), .A2(new_n1152), .A3(new_n1153), .A4(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1114), .B1(G107), .B2(new_n798), .ZN(new_n1158));
  INV_X1    g0958(.A(G283), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1158), .B1(new_n1159), .B2(new_n858), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n793), .A2(G294), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n796), .A2(G116), .B1(new_n860), .B2(G97), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n804), .A2(G87), .B1(new_n806), .B2(G68), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1161), .A2(new_n264), .A3(new_n1162), .A4(new_n1163), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1157), .B1(new_n1160), .B2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1147), .B1(new_n1165), .B2(new_n821), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1133), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1166), .B1(new_n1167), .B2(new_n772), .ZN(new_n1168));
  NOR3_X1   g0968(.A1(new_n941), .A2(new_n942), .A3(new_n687), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n754), .ZN(new_n1170));
  OAI211_X1 g0970(.A(G330), .B(new_n838), .C1(new_n1169), .C2(new_n1170), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1171), .A2(new_n1138), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n846), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n912), .B1(new_n1142), .B2(new_n1173), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1171), .A2(new_n1138), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(new_n1143), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n1175), .A2(new_n1137), .B1(new_n1177), .B2(new_n950), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n651), .A2(new_n1142), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n650), .A2(new_n970), .A3(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(KEYINPUT120), .B1(new_n1178), .B2(new_n1180), .ZN(new_n1181));
  AND3_X1   g0981(.A1(new_n650), .A2(new_n970), .A3(new_n1179), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n880), .B(new_n846), .C1(new_n731), .C2(new_n919), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1140), .B1(new_n1183), .B2(new_n912), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n967), .A2(new_n684), .A3(new_n843), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(new_n836), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n1171), .A2(new_n1138), .B1(new_n924), .B2(new_n1142), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n950), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n1184), .A2(new_n1186), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT120), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1182), .A2(new_n1189), .A3(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1181), .A2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n701), .B1(new_n1192), .B2(new_n1145), .ZN(new_n1193));
  AND3_X1   g0993(.A1(new_n1182), .A2(new_n1189), .A3(new_n1190), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1190), .B1(new_n1182), .B2(new_n1189), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1135), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1197));
  AND2_X1   g0997(.A1(new_n1135), .A2(new_n1139), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1197), .B1(new_n1198), .B2(new_n1143), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1196), .A2(new_n1199), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1146), .B(new_n1168), .C1(new_n1193), .C2(new_n1200), .ZN(G378));
  NOR2_X1   g1001(.A1(new_n380), .A2(G41), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(G33), .A2(G41), .ZN(new_n1203));
  NOR3_X1   g1003(.A1(new_n1202), .A2(G50), .A3(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n785), .A2(G125), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1205), .B1(new_n856), .B2(new_n873), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1206), .B1(G150), .B2(new_n810), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n796), .A2(G128), .B1(new_n860), .B2(G137), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1207), .B(new_n1208), .C1(new_n803), .C2(new_n1154), .ZN(new_n1209));
  OR2_X1    g1009(.A1(new_n1209), .A2(KEYINPUT59), .ZN(new_n1210));
  INV_X1    g1010(.A(G124), .ZN(new_n1211));
  OAI221_X1 g1011(.A(new_n1203), .B1(new_n789), .B2(new_n1211), .C1(new_n377), .C2(new_n805), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(new_n1209), .B2(KEYINPUT59), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1204), .B1(new_n1210), .B2(new_n1213), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n795), .A2(new_n429), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT122), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n1215), .A2(new_n1216), .B1(new_n798), .B2(G97), .ZN(new_n1217));
  OAI221_X1 g1017(.A(new_n1217), .B1(new_n1216), .B2(new_n1215), .C1(new_n468), .C2(new_n858), .ZN(new_n1218));
  AOI211_X1 g1018(.A(new_n1041), .B(new_n1218), .C1(new_n463), .C2(new_n860), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n805), .A2(new_n373), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1077), .A2(new_n1202), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n1220), .B(new_n1221), .C1(new_n793), .C2(G283), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(new_n1222), .B(KEYINPUT121), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1219), .A2(new_n1223), .A3(KEYINPUT58), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1214), .A2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(KEYINPUT58), .B1(new_n1219), .B2(new_n1223), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n821), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n766), .B1(new_n295), .B2(new_n851), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n312), .A2(new_n683), .ZN(new_n1229));
  XNOR2_X1  g1029(.A(new_n318), .B(new_n1229), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1231));
  XNOR2_X1  g1031(.A(new_n1230), .B(new_n1231), .ZN(new_n1232));
  OAI211_X1 g1032(.A(new_n1227), .B(new_n1228), .C1(new_n1232), .C2(new_n772), .ZN(new_n1233));
  XOR2_X1   g1033(.A(new_n1233), .B(KEYINPUT123), .Z(new_n1234));
  NAND2_X1  g1034(.A1(new_n937), .A2(G330), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1232), .B1(new_n926), .B2(new_n1235), .ZN(new_n1236));
  AOI211_X1 g1036(.A(new_n359), .B(new_n903), .C1(new_n369), .C2(new_n370), .ZN(new_n1237));
  AND2_X1   g1037(.A1(new_n910), .A2(new_n902), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n838), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n922), .B1(new_n1239), .B2(new_n944), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1240), .A2(new_n925), .A3(new_n953), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(new_n927), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1235), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1232), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1242), .A2(new_n1243), .A3(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1236), .A2(new_n1245), .A3(KEYINPUT124), .ZN(new_n1246));
  AND3_X1   g1046(.A1(new_n956), .A2(new_n957), .A3(new_n965), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1236), .A2(new_n1245), .A3(new_n966), .A4(KEYINPUT124), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1234), .B1(new_n1250), .B2(new_n764), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1182), .B1(new_n1196), .B2(new_n1199), .ZN(new_n1252));
  AOI21_X1  g1052(.A(KEYINPUT57), .B1(new_n1252), .B2(new_n1250), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1180), .B1(new_n1192), .B2(new_n1145), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1244), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1255));
  AOI211_X1 g1055(.A(new_n1232), .B(new_n1235), .C1(new_n1241), .C2(new_n927), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n966), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1247), .A2(new_n1236), .A3(new_n1245), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1257), .A2(KEYINPUT57), .A3(new_n1258), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n701), .B1(new_n1254), .B2(new_n1259), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1251), .B1(new_n1253), .B2(new_n1260), .ZN(G375));
  OAI21_X1  g1061(.A(new_n765), .B1(G68), .B2(new_n852), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n785), .A2(G132), .ZN(new_n1263));
  OAI221_X1 g1063(.A(new_n1263), .B1(new_n867), .B2(new_n795), .C1(new_n856), .C2(new_n1154), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(KEYINPUT126), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n793), .A2(G128), .ZN(new_n1267));
  AOI211_X1 g1067(.A(new_n382), .B(new_n1220), .C1(G150), .C2(new_n860), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n810), .A2(G50), .B1(new_n804), .B2(G159), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1266), .A2(new_n1267), .A3(new_n1268), .A4(new_n1269), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1265), .A2(KEYINPUT126), .ZN(new_n1271));
  OAI22_X1  g1071(.A1(new_n777), .A2(new_n434), .B1(new_n795), .B2(new_n1159), .ZN(new_n1272));
  XNOR2_X1  g1072(.A(new_n1272), .B(KEYINPUT125), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n793), .A2(G303), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n258), .B1(G107), .B2(new_n860), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1039), .B1(G294), .B2(new_n785), .ZN(new_n1276));
  AOI22_X1  g1076(.A1(new_n798), .A2(G116), .B1(new_n804), .B2(G97), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1274), .A2(new_n1275), .A3(new_n1276), .A4(new_n1277), .ZN(new_n1278));
  OAI22_X1  g1078(.A1(new_n1270), .A2(new_n1271), .B1(new_n1273), .B2(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1262), .B1(new_n1279), .B2(new_n821), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1280), .B1(new_n912), .B2(new_n772), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1281), .B1(new_n1178), .B2(new_n763), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1178), .A2(new_n1180), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1181), .A2(new_n1191), .A3(new_n1284), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1283), .B1(new_n1285), .B2(new_n1011), .ZN(G381));
  INV_X1    g1086(.A(G375), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1146), .A2(new_n1168), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n702), .B1(new_n1196), .B2(new_n1199), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1192), .A2(new_n1145), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1288), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1291));
  NOR3_X1   g1091(.A1(G387), .A2(G384), .A3(G390), .ZN(new_n1292));
  NOR3_X1   g1092(.A1(G393), .A2(G396), .A3(G381), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1287), .A2(new_n1291), .A3(new_n1292), .A4(new_n1293), .ZN(G407));
  NOR2_X1   g1094(.A1(new_n680), .A2(G343), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1287), .A2(new_n1291), .A3(new_n1295), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(G407), .A2(new_n1296), .A3(G213), .ZN(G409));
  INV_X1    g1097(.A(KEYINPUT63), .ZN(new_n1298));
  OAI211_X1 g1098(.A(G378), .B(new_n1251), .C1(new_n1253), .C2(new_n1260), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1011), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1252), .A2(new_n1300), .A3(new_n1250), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1257), .A2(new_n764), .A3(new_n1258), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1234), .ZN(new_n1303));
  AND2_X1   g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1301), .A2(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(new_n1291), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1299), .A2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1295), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1285), .A2(KEYINPUT60), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1182), .A2(new_n1189), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n701), .B1(new_n1311), .B2(KEYINPUT60), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1310), .A2(new_n1313), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1314), .A2(G384), .A3(new_n1283), .ZN(new_n1315));
  AND2_X1   g1115(.A1(new_n850), .A2(new_n877), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1312), .B1(new_n1285), .B2(KEYINPUT60), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1316), .B1(new_n1317), .B2(new_n1282), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1315), .A2(new_n1318), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1298), .B1(new_n1309), .B2(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1295), .A2(G2897), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1321), .ZN(new_n1322));
  AOI21_X1  g1122(.A(G384), .B1(new_n1314), .B2(new_n1283), .ZN(new_n1323));
  NOR3_X1   g1123(.A1(new_n1317), .A2(new_n1316), .A3(new_n1282), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1322), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1315), .A2(new_n1318), .A3(new_n1321), .ZN(new_n1326));
  AND2_X1   g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  AOI21_X1  g1127(.A(KEYINPUT61), .B1(new_n1309), .B2(new_n1327), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1033), .A2(G390), .A3(new_n1055), .ZN(new_n1329));
  INV_X1    g1129(.A(new_n1329), .ZN(new_n1330));
  AOI21_X1  g1130(.A(G390), .B1(new_n1033), .B2(new_n1055), .ZN(new_n1331));
  AOI211_X1 g1131(.A(G396), .B(new_n1099), .C1(new_n1060), .C2(new_n1062), .ZN(new_n1332));
  INV_X1    g1132(.A(G396), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1333), .B1(new_n1063), .B2(new_n1100), .ZN(new_n1334));
  OAI22_X1  g1134(.A1(new_n1330), .A2(new_n1331), .B1(new_n1332), .B2(new_n1334), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(G387), .A2(new_n1131), .A3(new_n1128), .ZN(new_n1336));
  NOR2_X1   g1136(.A1(new_n1334), .A2(new_n1332), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1336), .A2(new_n1337), .A3(new_n1329), .ZN(new_n1338));
  AND2_X1   g1138(.A1(new_n1335), .A2(new_n1338), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1295), .B1(new_n1299), .B2(new_n1306), .ZN(new_n1340));
  INV_X1    g1140(.A(new_n1319), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1340), .A2(KEYINPUT63), .A3(new_n1341), .ZN(new_n1342));
  NAND4_X1  g1142(.A1(new_n1320), .A2(new_n1328), .A3(new_n1339), .A4(new_n1342), .ZN(new_n1343));
  INV_X1    g1143(.A(KEYINPUT62), .ZN(new_n1344));
  AND3_X1   g1144(.A1(new_n1340), .A2(new_n1344), .A3(new_n1341), .ZN(new_n1345));
  INV_X1    g1145(.A(KEYINPUT61), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1347));
  OAI21_X1  g1147(.A(new_n1346), .B1(new_n1340), .B2(new_n1347), .ZN(new_n1348));
  AOI21_X1  g1148(.A(new_n1344), .B1(new_n1340), .B2(new_n1341), .ZN(new_n1349));
  NOR3_X1   g1149(.A1(new_n1345), .A2(new_n1348), .A3(new_n1349), .ZN(new_n1350));
  OAI21_X1  g1150(.A(new_n1343), .B1(new_n1350), .B2(new_n1339), .ZN(G405));
  NAND2_X1  g1151(.A1(new_n1319), .A2(KEYINPUT127), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1339), .A2(new_n1352), .ZN(new_n1353));
  OAI21_X1  g1153(.A(new_n1299), .B1(new_n1319), .B2(KEYINPUT127), .ZN(new_n1354));
  AOI21_X1  g1154(.A(new_n1354), .B1(new_n1291), .B2(G375), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1335), .A2(new_n1338), .ZN(new_n1356));
  NAND3_X1  g1156(.A1(new_n1356), .A2(KEYINPUT127), .A3(new_n1319), .ZN(new_n1357));
  AND3_X1   g1157(.A1(new_n1353), .A2(new_n1355), .A3(new_n1357), .ZN(new_n1358));
  AOI21_X1  g1158(.A(new_n1355), .B1(new_n1353), .B2(new_n1357), .ZN(new_n1359));
  NOR2_X1   g1159(.A1(new_n1358), .A2(new_n1359), .ZN(G402));
endmodule


