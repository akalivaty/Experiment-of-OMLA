//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 0 1 0 0 1 0 0 1 0 0 0 1 0 0 0 1 1 1 1 1 1 1 0 0 0 0 0 0 0 1 1 1 0 0 0 0 0 1 0 1 0 1 1 1 1 0 0 1 0 0 0 0 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:13 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n550, new_n552, new_n553,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n576, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n597, new_n598, new_n599, new_n602, new_n604, new_n605,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n813, new_n814, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1188;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT65), .B(G2066), .ZN(G411));
  XNOR2_X1  g006(.A(KEYINPUT66), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n461), .A2(new_n463), .A3(G125), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n459), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n461), .A2(new_n463), .A3(G137), .ZN(new_n467));
  NAND2_X1  g042(.A1(G101), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(G2105), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n466), .A2(new_n469), .ZN(G160));
  NAND2_X1  g045(.A1(new_n461), .A2(new_n463), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n471), .A2(new_n459), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G124), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n471), .A2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G136), .ZN(new_n475));
  NOR2_X1   g050(.A1(G100), .A2(G2105), .ZN(new_n476));
  OAI21_X1  g051(.A(G2104), .B1(new_n459), .B2(G112), .ZN(new_n477));
  OAI211_X1 g052(.A(new_n473), .B(new_n475), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G162));
  NAND4_X1  g054(.A1(new_n461), .A2(new_n463), .A3(G126), .A4(G2105), .ZN(new_n480));
  OR2_X1    g055(.A1(G102), .A2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(G114), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n481), .A2(new_n483), .A3(G2104), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n480), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(KEYINPUT67), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n461), .A2(new_n463), .A3(G138), .A4(new_n459), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  XNOR2_X1  g064(.A(KEYINPUT3), .B(G2104), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n490), .A2(KEYINPUT4), .A3(G138), .A4(new_n459), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT67), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n480), .A2(new_n492), .A3(new_n484), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n486), .A2(new_n489), .A3(new_n491), .A4(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(G164));
  NAND2_X1  g070(.A1(G75), .A2(G543), .ZN(new_n496));
  INV_X1    g071(.A(G543), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT5), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT5), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(G543), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(G62), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n496), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(G651), .ZN(new_n505));
  OAI21_X1  g080(.A(KEYINPUT70), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT70), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n503), .A2(new_n507), .A3(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT6), .ZN(new_n510));
  OAI21_X1  g085(.A(KEYINPUT68), .B1(new_n510), .B2(G651), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT68), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n512), .A2(new_n505), .A3(KEYINPUT6), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n510), .A2(G651), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT5), .B(G543), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT69), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND4_X1  g094(.A1(new_n514), .A2(KEYINPUT69), .A3(new_n515), .A4(new_n516), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n519), .A2(G88), .A3(new_n520), .ZN(new_n521));
  AND3_X1   g096(.A1(new_n514), .A2(G543), .A3(new_n515), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G50), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n509), .A2(new_n521), .A3(new_n523), .ZN(G303));
  INV_X1    g099(.A(G303), .ZN(G166));
  NAND2_X1  g100(.A1(new_n519), .A2(new_n520), .ZN(new_n526));
  INV_X1    g101(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G89), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT7), .ZN(new_n530));
  AND2_X1   g105(.A1(new_n516), .A2(G63), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n522), .A2(G51), .B1(G651), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n528), .A2(new_n530), .A3(new_n532), .ZN(G286));
  INV_X1    g108(.A(G286), .ZN(G168));
  NAND2_X1  g109(.A1(new_n527), .A2(G90), .ZN(new_n535));
  NAND2_X1  g110(.A1(G77), .A2(G543), .ZN(new_n536));
  INV_X1    g111(.A(G64), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n536), .B1(new_n501), .B2(new_n537), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n522), .A2(G52), .B1(G651), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n535), .A2(new_n539), .ZN(G301));
  INV_X1    g115(.A(G301), .ZN(G171));
  NAND3_X1  g116(.A1(new_n519), .A2(G81), .A3(new_n520), .ZN(new_n542));
  NAND2_X1  g117(.A1(G68), .A2(G543), .ZN(new_n543));
  INV_X1    g118(.A(G56), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n543), .B1(new_n501), .B2(new_n544), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n522), .A2(G43), .B1(G651), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n542), .A2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  AND3_X1   g124(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G36), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n550), .A2(new_n553), .ZN(G188));
  AND3_X1   g129(.A1(new_n519), .A2(G91), .A3(new_n520), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n522), .A2(G53), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT71), .ZN(new_n558));
  AOI21_X1  g133(.A(KEYINPUT72), .B1(new_n558), .B2(KEYINPUT9), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(G78), .A2(G543), .ZN(new_n561));
  XOR2_X1   g136(.A(KEYINPUT73), .B(G65), .Z(new_n562));
  OAI21_X1  g137(.A(new_n561), .B1(new_n562), .B2(new_n501), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G651), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n559), .B1(KEYINPUT72), .B2(KEYINPUT9), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n522), .A2(G53), .A3(new_n565), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n556), .A2(new_n560), .A3(new_n564), .A4(new_n566), .ZN(G299));
  OR2_X1    g142(.A1(new_n516), .A2(G74), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n522), .A2(G49), .B1(new_n568), .B2(G651), .ZN(new_n569));
  INV_X1    g144(.A(G87), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n526), .B2(new_n570), .ZN(G288));
  NAND3_X1  g146(.A1(new_n519), .A2(G86), .A3(new_n520), .ZN(new_n572));
  NAND2_X1  g147(.A1(G73), .A2(G543), .ZN(new_n573));
  INV_X1    g148(.A(G61), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n501), .B2(new_n574), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n522), .A2(G48), .B1(G651), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n572), .A2(new_n576), .ZN(G305));
  NAND2_X1  g152(.A1(new_n527), .A2(G85), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n516), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n579), .A2(new_n505), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n580), .B(KEYINPUT74), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n522), .A2(G47), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n578), .A2(new_n581), .A3(new_n582), .ZN(G290));
  NAND2_X1  g158(.A1(G301), .A2(G868), .ZN(new_n584));
  INV_X1    g159(.A(G92), .ZN(new_n585));
  OR3_X1    g160(.A1(new_n526), .A2(KEYINPUT10), .A3(new_n585), .ZN(new_n586));
  OAI21_X1  g161(.A(KEYINPUT10), .B1(new_n526), .B2(new_n585), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(G79), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G66), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n501), .B2(new_n590), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n522), .A2(G54), .B1(G651), .B2(new_n591), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n592), .B(KEYINPUT75), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n588), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n584), .B1(new_n594), .B2(G868), .ZN(G284));
  OAI21_X1  g170(.A(new_n584), .B1(new_n594), .B2(G868), .ZN(G321));
  NAND2_X1  g171(.A1(G286), .A2(G868), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n560), .A2(new_n564), .A3(new_n566), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n598), .A2(new_n555), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n597), .B1(new_n599), .B2(G868), .ZN(G297));
  OAI21_X1  g175(.A(new_n597), .B1(new_n599), .B2(G868), .ZN(G280));
  XOR2_X1   g176(.A(KEYINPUT76), .B(G559), .Z(new_n602));
  OAI21_X1  g177(.A(new_n594), .B1(G860), .B2(new_n602), .ZN(G148));
  NAND2_X1  g178(.A1(new_n594), .A2(new_n602), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n604), .A2(G868), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(G868), .B2(new_n548), .ZN(G323));
  XNOR2_X1  g181(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g182(.A1(new_n474), .A2(G2104), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT12), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT13), .ZN(new_n610));
  XOR2_X1   g185(.A(KEYINPUT77), .B(G2100), .Z(new_n611));
  XNOR2_X1  g186(.A(new_n610), .B(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n474), .A2(G135), .ZN(new_n613));
  OR2_X1    g188(.A1(G99), .A2(G2105), .ZN(new_n614));
  OAI211_X1 g189(.A(new_n614), .B(G2104), .C1(G111), .C2(new_n459), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n616), .B1(G123), .B2(new_n472), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(G2096), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n612), .A2(new_n618), .ZN(G156));
  XNOR2_X1  g194(.A(G2451), .B(G2454), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT78), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT16), .ZN(new_n622));
  XOR2_X1   g197(.A(G2443), .B(G2446), .Z(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XOR2_X1   g199(.A(G1341), .B(G1348), .Z(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(G2427), .B(G2438), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2430), .ZN(new_n628));
  XOR2_X1   g203(.A(KEYINPUT15), .B(G2435), .Z(new_n629));
  XOR2_X1   g204(.A(new_n628), .B(new_n629), .Z(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(KEYINPUT14), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n626), .B(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(G14), .ZN(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(G401));
  XOR2_X1   g209(.A(G2072), .B(G2078), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT79), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT81), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT17), .ZN(new_n638));
  XOR2_X1   g213(.A(G2067), .B(G2678), .Z(new_n639));
  XOR2_X1   g214(.A(G2084), .B(G2090), .Z(new_n640));
  NAND3_X1  g215(.A1(new_n638), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  INV_X1    g216(.A(new_n639), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n636), .A2(new_n642), .A3(new_n640), .ZN(new_n643));
  XOR2_X1   g218(.A(KEYINPUT80), .B(KEYINPUT18), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  INV_X1    g220(.A(new_n640), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n646), .B1(new_n638), .B2(new_n639), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n636), .A2(new_n642), .ZN(new_n648));
  OAI211_X1 g223(.A(new_n641), .B(new_n645), .C1(new_n647), .C2(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2096), .B(G2100), .ZN(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n649), .A2(new_n651), .ZN(new_n653));
  AND2_X1   g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(G227));
  INV_X1    g230(.A(KEYINPUT20), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1956), .B(G2474), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT82), .ZN(new_n658));
  XOR2_X1   g233(.A(G1961), .B(G1966), .Z(new_n659));
  NAND2_X1  g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1971), .B(G1976), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT19), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n656), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n658), .A2(new_n659), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n665), .A2(new_n662), .A3(new_n660), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n660), .A2(new_n656), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n667), .A2(new_n664), .ZN(new_n668));
  OAI211_X1 g243(.A(new_n663), .B(new_n666), .C1(new_n668), .C2(new_n662), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(G1991), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(G1981), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1986), .B(G1996), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n670), .B(new_n674), .ZN(G229));
  AND2_X1   g250(.A1(KEYINPUT24), .A2(G34), .ZN(new_n676));
  NOR2_X1   g251(.A1(KEYINPUT24), .A2(G34), .ZN(new_n677));
  NOR3_X1   g252(.A1(new_n676), .A2(new_n677), .A3(G29), .ZN(new_n678));
  INV_X1    g253(.A(G160), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n678), .B1(new_n679), .B2(G29), .ZN(new_n680));
  INV_X1    g255(.A(G2084), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(G29), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n684), .A2(G26), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT28), .ZN(new_n686));
  AOI22_X1  g261(.A1(G128), .A2(new_n472), .B1(new_n474), .B2(G140), .ZN(new_n687));
  OR2_X1    g262(.A1(G104), .A2(G2105), .ZN(new_n688));
  INV_X1    g263(.A(KEYINPUT85), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n460), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  OAI221_X1 g265(.A(new_n690), .B1(new_n689), .B2(new_n688), .C1(G116), .C2(new_n459), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n687), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(G29), .ZN(new_n693));
  AND2_X1   g268(.A1(new_n693), .A2(KEYINPUT86), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n693), .A2(KEYINPUT86), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n686), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(G2067), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(G16), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G19), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(new_n548), .B2(new_n699), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n594), .A2(new_n699), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n702), .B1(G4), .B2(new_n699), .ZN(new_n703));
  INV_X1    g278(.A(G1348), .ZN(new_n704));
  OAI221_X1 g279(.A(new_n698), .B1(G1341), .B2(new_n701), .C1(new_n703), .C2(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n617), .A2(G29), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(KEYINPUT92), .Z(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT31), .B(G11), .ZN(new_n708));
  INV_X1    g283(.A(KEYINPUT30), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n709), .A2(G28), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(G28), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n710), .A2(new_n711), .A3(new_n684), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n707), .A2(new_n708), .A3(new_n712), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(KEYINPUT93), .Z(new_n714));
  AOI211_X1 g289(.A(new_n705), .B(new_n714), .C1(new_n704), .C2(new_n703), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n684), .A2(G33), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(KEYINPUT25), .Z(new_n718));
  NAND2_X1  g293(.A1(new_n474), .A2(G139), .ZN(new_n719));
  AOI22_X1  g294(.A1(new_n490), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n720));
  OAI211_X1 g295(.A(new_n718), .B(new_n719), .C1(new_n459), .C2(new_n720), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT87), .Z(new_n722));
  OAI21_X1  g297(.A(new_n716), .B1(new_n722), .B2(new_n684), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(G2072), .Z(new_n724));
  NAND2_X1  g299(.A1(new_n472), .A2(G129), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n474), .A2(G141), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n459), .A2(G105), .A3(G2104), .ZN(new_n727));
  NAND3_X1  g302(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT26), .Z(new_n729));
  NAND4_X1  g304(.A1(new_n725), .A2(new_n726), .A3(new_n727), .A4(new_n729), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT89), .Z(new_n731));
  NOR2_X1   g306(.A1(new_n731), .A2(new_n684), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(new_n684), .B2(G32), .ZN(new_n733));
  XNOR2_X1  g308(.A(KEYINPUT27), .B(G1996), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n680), .A2(new_n681), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT88), .Z(new_n737));
  NAND3_X1  g312(.A1(new_n724), .A2(new_n735), .A3(new_n737), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT90), .Z(new_n739));
  NAND2_X1  g314(.A1(new_n699), .A2(G20), .ZN(new_n740));
  OAI211_X1 g315(.A(KEYINPUT23), .B(new_n740), .C1(new_n599), .C2(new_n699), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(KEYINPUT23), .B2(new_n740), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(G1956), .ZN(new_n743));
  NAND2_X1  g318(.A1(G168), .A2(G16), .ZN(new_n744));
  NOR2_X1   g319(.A1(G16), .A2(G21), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n744), .B1(KEYINPUT91), .B2(new_n745), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(KEYINPUT91), .B2(new_n744), .ZN(new_n747));
  INV_X1    g322(.A(G1966), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  NOR2_X1   g324(.A1(G164), .A2(new_n684), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(G27), .B2(new_n684), .ZN(new_n751));
  INV_X1    g326(.A(new_n751), .ZN(new_n752));
  OAI22_X1  g327(.A1(new_n733), .A2(new_n734), .B1(G2078), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n684), .A2(G35), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G162), .B2(new_n684), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT29), .B(G2090), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(G5), .A2(G16), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(G171), .B2(G16), .ZN(new_n759));
  AOI22_X1  g334(.A1(G1961), .A2(new_n759), .B1(new_n752), .B2(G2078), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n701), .A2(G1341), .ZN(new_n761));
  OAI211_X1 g336(.A(new_n760), .B(new_n761), .C1(G1961), .C2(new_n759), .ZN(new_n762));
  NOR4_X1   g337(.A1(new_n749), .A2(new_n753), .A3(new_n757), .A4(new_n762), .ZN(new_n763));
  NAND4_X1  g338(.A1(new_n715), .A2(new_n739), .A3(new_n743), .A4(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n684), .A2(G25), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n472), .A2(G119), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n474), .A2(G131), .ZN(new_n767));
  OR2_X1    g342(.A1(G95), .A2(G2105), .ZN(new_n768));
  OAI211_X1 g343(.A(new_n768), .B(G2104), .C1(G107), .C2(new_n459), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n766), .A2(new_n767), .A3(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n765), .B1(new_n771), .B2(new_n684), .ZN(new_n772));
  XNOR2_X1  g347(.A(KEYINPUT35), .B(G1991), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(G290), .A2(G16), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n699), .A2(G24), .ZN(new_n776));
  AND2_X1   g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(new_n777), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n774), .B1(new_n778), .B2(G1986), .ZN(new_n779));
  INV_X1    g354(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n699), .A2(G23), .ZN(new_n781));
  INV_X1    g356(.A(G288), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n781), .B1(new_n782), .B2(new_n699), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT33), .ZN(new_n784));
  INV_X1    g359(.A(G1976), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n699), .A2(G22), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(G166), .B2(new_n699), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT83), .B(G1971), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  MUX2_X1   g365(.A(G6), .B(G305), .S(G16), .Z(new_n791));
  XOR2_X1   g366(.A(KEYINPUT32), .B(G1981), .Z(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  OR2_X1    g368(.A1(new_n783), .A2(KEYINPUT33), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n783), .A2(KEYINPUT33), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n794), .A2(G1976), .A3(new_n795), .ZN(new_n796));
  NAND4_X1  g371(.A1(new_n786), .A2(new_n790), .A3(new_n793), .A4(new_n796), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT84), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n780), .B1(new_n798), .B2(KEYINPUT34), .ZN(new_n799));
  INV_X1    g374(.A(G1986), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n777), .A2(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT84), .ZN(new_n802));
  OR2_X1    g377(.A1(new_n797), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n797), .A2(new_n802), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT34), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n799), .A2(new_n801), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n808), .A2(KEYINPUT36), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT36), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n799), .A2(new_n810), .A3(new_n807), .A4(new_n801), .ZN(new_n811));
  AOI211_X1 g386(.A(new_n683), .B(new_n764), .C1(new_n809), .C2(new_n811), .ZN(G311));
  NAND2_X1  g387(.A1(new_n809), .A2(new_n811), .ZN(new_n813));
  INV_X1    g388(.A(new_n764), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n813), .A2(new_n682), .A3(new_n814), .ZN(G150));
  NAND2_X1  g390(.A1(new_n522), .A2(G55), .ZN(new_n816));
  AOI22_X1  g391(.A1(new_n516), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n817));
  XNOR2_X1  g392(.A(KEYINPUT94), .B(G93), .ZN(new_n818));
  OAI221_X1 g393(.A(new_n816), .B1(new_n505), .B2(new_n817), .C1(new_n526), .C2(new_n818), .ZN(new_n819));
  XOR2_X1   g394(.A(KEYINPUT97), .B(G860), .Z(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(KEYINPUT37), .Z(new_n822));
  NAND2_X1  g397(.A1(new_n594), .A2(G559), .ZN(new_n823));
  XOR2_X1   g398(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n824));
  XNOR2_X1  g399(.A(new_n823), .B(new_n824), .ZN(new_n825));
  OR3_X1    g400(.A1(new_n547), .A2(KEYINPUT95), .A3(KEYINPUT96), .ZN(new_n826));
  OAI21_X1  g401(.A(KEYINPUT96), .B1(new_n547), .B2(KEYINPUT95), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n547), .A2(KEYINPUT95), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(new_n819), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  NAND4_X1  g406(.A1(new_n826), .A2(new_n829), .A3(new_n819), .A4(new_n827), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n825), .B(new_n833), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n822), .B1(new_n834), .B2(new_n820), .ZN(G145));
  NAND4_X1  g410(.A1(new_n489), .A2(new_n491), .A3(new_n480), .A4(new_n484), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT99), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(new_n770), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n472), .A2(G130), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n474), .A2(G142), .ZN(new_n840));
  NOR2_X1   g415(.A1(G106), .A2(G2105), .ZN(new_n841));
  OAI21_X1  g416(.A(G2104), .B1(new_n459), .B2(G118), .ZN(new_n842));
  OAI211_X1 g417(.A(new_n839), .B(new_n840), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT98), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n838), .B(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n609), .B(new_n692), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n730), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n722), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n849), .B1(new_n731), .B2(new_n722), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n617), .B(new_n679), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(G162), .ZN(new_n853));
  OR2_X1    g428(.A1(new_n845), .A2(new_n846), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n845), .A2(new_n846), .ZN(new_n855));
  INV_X1    g430(.A(new_n850), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  AND3_X1   g432(.A1(new_n851), .A2(new_n853), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n853), .B1(new_n851), .B2(new_n857), .ZN(new_n859));
  OR3_X1    g434(.A1(new_n858), .A2(new_n859), .A3(G37), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g436(.A1(new_n819), .A2(G868), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT42), .ZN(new_n863));
  XOR2_X1   g438(.A(G288), .B(G305), .Z(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(G303), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(G290), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT103), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(G290), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n865), .B(new_n869), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n870), .A2(KEYINPUT103), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n863), .B1(new_n868), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n870), .A2(KEYINPUT103), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n866), .A2(new_n867), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n873), .A2(new_n874), .A3(KEYINPUT42), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT104), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n833), .B(new_n604), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  OAI21_X1  g454(.A(G299), .B1(new_n588), .B2(new_n593), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT75), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n592), .B(new_n881), .ZN(new_n882));
  NAND4_X1  g457(.A1(new_n599), .A2(new_n882), .A3(new_n587), .A4(new_n586), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(KEYINPUT100), .ZN(new_n885));
  OR2_X1    g460(.A1(new_n879), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT101), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT41), .ZN(new_n888));
  NAND4_X1  g463(.A1(new_n880), .A2(new_n883), .A3(new_n887), .A4(new_n888), .ZN(new_n889));
  OAI21_X1  g464(.A(KEYINPUT101), .B1(new_n884), .B2(KEYINPUT41), .ZN(new_n890));
  AOI21_X1  g465(.A(KEYINPUT102), .B1(new_n884), .B2(KEYINPUT41), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT102), .ZN(new_n892));
  AOI211_X1 g467(.A(new_n892), .B(new_n888), .C1(new_n880), .C2(new_n883), .ZN(new_n893));
  OAI211_X1 g468(.A(new_n889), .B(new_n890), .C1(new_n891), .C2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n886), .B1(new_n895), .B2(new_n878), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n876), .A2(new_n877), .A3(new_n896), .ZN(new_n897));
  OAI211_X1 g472(.A(new_n886), .B(KEYINPUT104), .C1(new_n878), .C2(new_n895), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n895), .A2(new_n878), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n879), .A2(new_n885), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n877), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND4_X1  g476(.A1(new_n898), .A2(new_n875), .A3(new_n872), .A4(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n897), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n862), .B1(new_n903), .B2(G868), .ZN(G295));
  AOI21_X1  g479(.A(new_n862), .B1(new_n903), .B2(G868), .ZN(G331));
  AOI21_X1  g480(.A(G286), .B1(G171), .B2(KEYINPUT105), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  OR2_X1    g482(.A1(G171), .A2(KEYINPUT105), .ZN(new_n908));
  AND3_X1   g483(.A1(new_n831), .A2(new_n832), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n908), .B1(new_n831), .B2(new_n832), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n907), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n908), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n833), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n831), .A2(new_n832), .A3(new_n908), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n913), .A2(new_n906), .A3(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n911), .A2(new_n915), .A3(new_n884), .ZN(new_n916));
  AND2_X1   g491(.A1(new_n911), .A2(new_n915), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n916), .B1(new_n917), .B2(new_n894), .ZN(new_n918));
  AOI21_X1  g493(.A(G37), .B1(new_n918), .B2(new_n870), .ZN(new_n919));
  OAI211_X1 g494(.A(new_n866), .B(new_n916), .C1(new_n917), .C2(new_n894), .ZN(new_n920));
  AOI21_X1  g495(.A(KEYINPUT43), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n894), .B1(new_n915), .B2(new_n911), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n911), .A2(new_n915), .A3(new_n884), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n870), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(G37), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n911), .A2(new_n915), .A3(new_n885), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n884), .B(KEYINPUT41), .ZN(new_n927));
  OAI211_X1 g502(.A(new_n926), .B(new_n866), .C1(new_n917), .C2(new_n927), .ZN(new_n928));
  AND4_X1   g503(.A1(KEYINPUT43), .A2(new_n924), .A3(new_n925), .A4(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(KEYINPUT44), .B1(new_n921), .B2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT44), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT43), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n932), .B1(new_n919), .B2(new_n920), .ZN(new_n933));
  AND4_X1   g508(.A1(new_n932), .A2(new_n924), .A3(new_n925), .A4(new_n928), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n931), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n930), .A2(new_n935), .ZN(G397));
  INV_X1    g511(.A(G1384), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n836), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n938), .B(KEYINPUT106), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT45), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n464), .A2(new_n465), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(G2105), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n467), .A2(new_n468), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(new_n459), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n943), .A2(new_n945), .A3(G40), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT107), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(G160), .A2(KEYINPUT107), .A3(G40), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n941), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(G1996), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n848), .A2(new_n952), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n692), .B(new_n697), .ZN(new_n954));
  INV_X1    g529(.A(new_n954), .ZN(new_n955));
  AOI211_X1 g530(.A(new_n953), .B(new_n955), .C1(new_n952), .C2(new_n731), .ZN(new_n956));
  INV_X1    g531(.A(new_n773), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n771), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n770), .A2(new_n773), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n956), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  XNOR2_X1  g535(.A(G290), .B(G1986), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n951), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT108), .ZN(new_n963));
  AND3_X1   g538(.A1(new_n480), .A2(new_n492), .A3(new_n484), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n492), .B1(new_n480), .B2(new_n484), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n489), .A2(new_n491), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(G1384), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n963), .B1(new_n969), .B2(KEYINPUT45), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n836), .A2(KEYINPUT45), .A3(new_n937), .ZN(new_n971));
  AND3_X1   g546(.A1(new_n948), .A2(new_n949), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n494), .A2(new_n937), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n973), .A2(KEYINPUT108), .A3(new_n940), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n970), .A2(new_n972), .A3(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(G1971), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT50), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n977), .B1(new_n494), .B2(new_n937), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n938), .A2(KEYINPUT50), .ZN(new_n979));
  NOR3_X1   g554(.A1(new_n950), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(G2090), .ZN(new_n981));
  AOI22_X1  g556(.A1(new_n975), .A2(new_n976), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(KEYINPUT109), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT55), .ZN(new_n986));
  INV_X1    g561(.A(G8), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n986), .B1(G166), .B2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT109), .ZN(new_n989));
  NAND4_X1  g564(.A1(G303), .A2(new_n989), .A3(KEYINPUT55), .A4(G8), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n985), .A2(new_n988), .A3(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n983), .A2(G8), .A3(new_n991), .ZN(new_n992));
  AND3_X1   g567(.A1(new_n985), .A2(new_n988), .A3(new_n990), .ZN(new_n993));
  AOI21_X1  g568(.A(KEYINPUT107), .B1(G160), .B2(G40), .ZN(new_n994));
  AND4_X1   g569(.A1(KEYINPUT107), .A2(new_n943), .A3(new_n945), .A4(G40), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n938), .A2(KEYINPUT50), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n494), .A2(new_n977), .A3(new_n937), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n996), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  AOI22_X1  g575(.A1(new_n981), .A2(new_n1000), .B1(new_n975), .B2(new_n976), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n993), .B1(new_n1001), .B2(new_n987), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT111), .ZN(new_n1003));
  INV_X1    g578(.A(new_n938), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1004), .A2(new_n948), .A3(new_n949), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT52), .ZN(new_n1006));
  OAI211_X1 g581(.A(new_n569), .B(G1976), .C1(new_n526), .C2(new_n570), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n1005), .A2(new_n1006), .A3(G8), .A4(new_n1007), .ZN(new_n1008));
  XOR2_X1   g583(.A(KEYINPUT110), .B(G1976), .Z(new_n1009));
  AND2_X1   g584(.A1(G288), .A2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1003), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n987), .B1(new_n996), .B2(new_n1004), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT113), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1013), .A2(KEYINPUT49), .ZN(new_n1014));
  INV_X1    g589(.A(G1981), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n572), .A2(new_n576), .A3(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g591(.A(KEYINPUT112), .B(G86), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n519), .A2(new_n520), .A3(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1015), .B1(new_n1018), .B2(new_n576), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1014), .B1(new_n1016), .B2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n572), .A2(new_n576), .A3(new_n1015), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1014), .ZN(new_n1022));
  AND2_X1   g597(.A1(new_n1018), .A2(new_n576), .ZN(new_n1023));
  OAI211_X1 g598(.A(new_n1021), .B(new_n1022), .C1(new_n1023), .C2(new_n1015), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1012), .A2(new_n1020), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1005), .A2(G8), .A3(new_n1007), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(KEYINPUT52), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1028), .B1(new_n1010), .B2(new_n1008), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1026), .B1(new_n1029), .B2(KEYINPUT111), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n992), .A2(new_n1002), .A3(new_n1011), .A4(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT51), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT115), .ZN(new_n1034));
  AOI21_X1  g609(.A(KEYINPUT45), .B1(new_n836), .B2(new_n937), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1034), .B1(new_n950), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n969), .A2(KEYINPUT45), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1035), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1038), .A2(KEYINPUT115), .A3(new_n948), .A4(new_n949), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1036), .A2(new_n1037), .A3(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(new_n748), .ZN(new_n1041));
  XOR2_X1   g616(.A(KEYINPUT116), .B(G2084), .Z(new_n1042));
  NAND2_X1  g617(.A1(new_n980), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1041), .A2(G168), .A3(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1033), .B1(new_n1044), .B2(G8), .ZN(new_n1045));
  AOI22_X1  g620(.A1(new_n1040), .A2(new_n748), .B1(new_n980), .B2(new_n1042), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n987), .B1(new_n1046), .B2(G168), .ZN(new_n1047));
  OAI21_X1  g622(.A(KEYINPUT51), .B1(new_n1046), .B2(G168), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1045), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT62), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1032), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1048), .A2(new_n1047), .ZN(new_n1052));
  AOI221_X4 g627(.A(G286), .B1(new_n980), .B2(new_n1042), .C1(new_n1040), .C2(new_n748), .ZN(new_n1053));
  OAI21_X1  g628(.A(KEYINPUT51), .B1(new_n1053), .B2(new_n987), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1052), .A2(new_n1054), .A3(new_n1050), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n980), .A2(G1961), .ZN(new_n1056));
  OR2_X1    g631(.A1(new_n975), .A2(G2078), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT53), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1056), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1058), .A2(G2078), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1036), .A2(new_n1060), .A3(new_n1037), .A4(new_n1039), .ZN(new_n1061));
  AOI21_X1  g636(.A(G301), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1055), .A2(new_n1062), .ZN(new_n1063));
  NOR3_X1   g638(.A1(new_n1051), .A2(KEYINPUT125), .A3(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT125), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1062), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1066), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1031), .B1(new_n1068), .B2(KEYINPUT62), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1065), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT117), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT63), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1000), .A2(new_n981), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n975), .A2(new_n976), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n987), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1072), .B1(new_n1075), .B2(new_n991), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1077), .A2(G8), .A3(G168), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n992), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1079));
  AND2_X1   g654(.A1(new_n1030), .A2(new_n1011), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NOR3_X1   g656(.A1(new_n1046), .A2(new_n987), .A3(G286), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n993), .B1(new_n982), .B2(new_n987), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1082), .A2(new_n1083), .A3(new_n1011), .A4(new_n1030), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(KEYINPUT63), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1025), .A2(new_n785), .A3(new_n782), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT114), .ZN(new_n1087));
  AND3_X1   g662(.A1(new_n1086), .A2(new_n1087), .A3(new_n1021), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1087), .B1(new_n1086), .B2(new_n1021), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(new_n1012), .ZN(new_n1091));
  AND4_X1   g666(.A1(new_n1071), .A2(new_n1081), .A3(new_n1085), .A4(new_n1091), .ZN(new_n1092));
  AOI22_X1  g667(.A1(KEYINPUT63), .A2(new_n1084), .B1(new_n1090), .B2(new_n1012), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1071), .B1(new_n1093), .B2(new_n1081), .ZN(new_n1094));
  OAI22_X1  g669(.A1(new_n1064), .A2(new_n1070), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT54), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1059), .A2(G301), .A3(new_n1061), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1096), .B1(new_n1097), .B2(KEYINPUT124), .ZN(new_n1098));
  INV_X1    g673(.A(new_n946), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n941), .A2(new_n1099), .A3(new_n971), .A4(new_n1060), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1059), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(G171), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT124), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1059), .A2(new_n1103), .A3(new_n1061), .A4(G301), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1098), .A2(new_n1102), .A3(new_n1104), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1101), .A2(G171), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1096), .B1(new_n1106), .B2(new_n1062), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1105), .A2(new_n1107), .A3(new_n1032), .A4(new_n1068), .ZN(new_n1108));
  AOI21_X1  g683(.A(KEYINPUT108), .B1(new_n973), .B2(new_n940), .ZN(new_n1109));
  AOI211_X1 g684(.A(new_n963), .B(KEYINPUT45), .C1(new_n494), .C2(new_n937), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT119), .ZN(new_n1112));
  XNOR2_X1  g687(.A(KEYINPUT56), .B(G2072), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1111), .A2(new_n1112), .A3(new_n1113), .A4(new_n972), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n970), .A2(new_n972), .A3(new_n1113), .A4(new_n974), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(KEYINPUT119), .ZN(new_n1116));
  INV_X1    g691(.A(G1956), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n999), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1114), .A2(new_n1116), .A3(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT118), .ZN(new_n1120));
  AOI21_X1  g695(.A(KEYINPUT57), .B1(G299), .B2(new_n1120), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n1120), .B(KEYINPUT57), .C1(new_n598), .C2(new_n555), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1122), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1119), .A2(new_n1125), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1124), .A2(new_n1114), .A3(new_n1116), .A4(new_n1118), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  XOR2_X1   g703(.A(KEYINPUT122), .B(KEYINPUT61), .Z(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT122), .ZN(new_n1131));
  OAI211_X1 g706(.A(new_n1126), .B(new_n1127), .C1(new_n1131), .C2(KEYINPUT61), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT120), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(KEYINPUT59), .ZN(new_n1134));
  XNOR2_X1  g709(.A(new_n1134), .B(KEYINPUT121), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1111), .A2(new_n952), .A3(new_n972), .ZN(new_n1136));
  XOR2_X1   g711(.A(KEYINPUT58), .B(G1341), .Z(new_n1137));
  NAND2_X1  g712(.A1(new_n1005), .A2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n547), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1133), .A2(KEYINPUT59), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1135), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1138), .B1(new_n975), .B2(G1996), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1140), .B1(new_n1142), .B2(new_n548), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1135), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1141), .A2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1130), .A2(new_n1132), .A3(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1147), .A2(KEYINPUT123), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT123), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1130), .A2(new_n1149), .A3(new_n1132), .A4(new_n1146), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1005), .A2(G2067), .ZN(new_n1151));
  INV_X1    g726(.A(new_n980), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1151), .B1(new_n1152), .B2(new_n704), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1153), .B1(KEYINPUT60), .B2(new_n594), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n594), .A2(KEYINPUT60), .ZN(new_n1155));
  XNOR2_X1  g730(.A(new_n1154), .B(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1148), .A2(new_n1150), .A3(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(new_n594), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1126), .B1(new_n1158), .B2(new_n1153), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1159), .A2(new_n1127), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1108), .B1(new_n1157), .B2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n962), .B1(new_n1095), .B2(new_n1161), .ZN(new_n1162));
  NOR3_X1   g737(.A1(new_n941), .A2(G1996), .A3(new_n950), .ZN(new_n1163));
  OR2_X1    g738(.A1(new_n1163), .A2(KEYINPUT46), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n951), .B1(new_n730), .B2(new_n955), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1163), .A2(KEYINPUT46), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1164), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1167));
  XOR2_X1   g742(.A(KEYINPUT126), .B(KEYINPUT47), .Z(new_n1168));
  XNOR2_X1  g743(.A(new_n1167), .B(new_n1168), .ZN(new_n1169));
  AND3_X1   g744(.A1(new_n956), .A2(new_n957), .A3(new_n771), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n692), .A2(G2067), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n951), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n960), .A2(new_n951), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n951), .A2(new_n800), .A3(new_n869), .ZN(new_n1174));
  XNOR2_X1  g749(.A(new_n1174), .B(KEYINPUT48), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1173), .A2(new_n1175), .ZN(new_n1176));
  AND3_X1   g751(.A1(new_n1169), .A2(new_n1172), .A3(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1162), .A2(new_n1177), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g753(.A(new_n860), .B1(new_n933), .B2(new_n934), .ZN(new_n1180));
  INV_X1    g754(.A(KEYINPUT127), .ZN(new_n1181));
  NAND2_X1  g755(.A1(new_n633), .A2(G319), .ZN(new_n1182));
  OAI21_X1  g756(.A(new_n1181), .B1(G227), .B2(new_n1182), .ZN(new_n1183));
  INV_X1    g757(.A(G229), .ZN(new_n1184));
  NAND4_X1  g758(.A1(new_n654), .A2(new_n633), .A3(KEYINPUT127), .A4(G319), .ZN(new_n1185));
  NAND3_X1  g759(.A1(new_n1183), .A2(new_n1184), .A3(new_n1185), .ZN(new_n1186));
  NOR2_X1   g760(.A1(new_n1180), .A2(new_n1186), .ZN(G308));
  INV_X1    g761(.A(new_n1186), .ZN(new_n1188));
  OAI211_X1 g762(.A(new_n1188), .B(new_n860), .C1(new_n933), .C2(new_n934), .ZN(G225));
endmodule


