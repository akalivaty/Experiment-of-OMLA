//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 1 1 0 1 1 1 0 1 0 0 1 1 0 0 0 0 0 1 1 0 0 1 1 0 0 0 0 1 1 0 0 1 0 0 1 1 0 1 0 1 1 1 1 1 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n709, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n738,
    new_n739, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n790, new_n791, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n816, new_n817,
    new_n818, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n883, new_n884,
    new_n885, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n995,
    new_n996;
  NAND2_X1  g000(.A1(G225gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(KEYINPUT2), .ZN(new_n205));
  INV_X1    g004(.A(G141gat), .ZN(new_n206));
  INV_X1    g005(.A(G148gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(G141gat), .A2(G148gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n205), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  OR2_X1    g009(.A1(G155gat), .A2(G162gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT74), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n211), .A2(new_n212), .A3(new_n204), .ZN(new_n213));
  AND2_X1   g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(G155gat), .A2(G162gat), .ZN(new_n215));
  OAI21_X1  g014(.A(KEYINPUT74), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n210), .A2(new_n213), .A3(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT75), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND4_X1  g018(.A1(new_n210), .A2(new_n213), .A3(new_n216), .A4(KEYINPUT75), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(G127gat), .B(G134gat), .ZN(new_n222));
  INV_X1    g021(.A(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(G113gat), .B(G120gat), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n223), .B1(KEYINPUT1), .B2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(new_n224), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT1), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n226), .A2(new_n227), .A3(new_n222), .ZN(new_n228));
  AND2_X1   g027(.A1(new_n225), .A2(new_n228), .ZN(new_n229));
  AND3_X1   g028(.A1(new_n204), .A2(KEYINPUT77), .A3(KEYINPUT2), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n214), .A2(new_n215), .ZN(new_n231));
  AOI21_X1  g030(.A(KEYINPUT77), .B1(new_n204), .B2(KEYINPUT2), .ZN(new_n232));
  NOR3_X1   g031(.A1(new_n230), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n208), .A2(new_n209), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(KEYINPUT76), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT76), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n208), .A2(new_n236), .A3(new_n209), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n233), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n221), .A2(new_n229), .A3(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  AOI22_X1  g040(.A1(new_n219), .A2(new_n220), .B1(new_n238), .B2(new_n233), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n242), .A2(new_n229), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n203), .B1(new_n241), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT4), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n240), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n242), .A2(KEYINPUT4), .A3(new_n229), .ZN(new_n247));
  INV_X1    g046(.A(new_n229), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT3), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n248), .B1(new_n242), .B2(new_n249), .ZN(new_n250));
  AND3_X1   g049(.A1(new_n221), .A2(new_n249), .A3(new_n239), .ZN(new_n251));
  OAI211_X1 g050(.A(new_n246), .B(new_n247), .C1(new_n250), .C2(new_n251), .ZN(new_n252));
  OAI211_X1 g051(.A(KEYINPUT5), .B(new_n244), .C1(new_n252), .C2(new_n203), .ZN(new_n253));
  AND2_X1   g052(.A1(new_n246), .A2(new_n247), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT5), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n221), .A2(new_n239), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(KEYINPUT3), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n242), .A2(new_n249), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n257), .A2(new_n258), .A3(new_n248), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n254), .A2(new_n255), .A3(new_n202), .A4(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n253), .A2(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(G1gat), .B(G29gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n262), .B(KEYINPUT0), .ZN(new_n263));
  XNOR2_X1  g062(.A(G57gat), .B(G85gat), .ZN(new_n264));
  XOR2_X1   g063(.A(new_n263), .B(new_n264), .Z(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  XOR2_X1   g065(.A(KEYINPUT78), .B(KEYINPUT6), .Z(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  AND4_X1   g067(.A1(KEYINPUT82), .A2(new_n261), .A3(new_n266), .A4(new_n268), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n265), .B1(new_n253), .B2(new_n260), .ZN(new_n270));
  AOI21_X1  g069(.A(KEYINPUT82), .B1(new_n270), .B2(new_n268), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT80), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n261), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n253), .A2(KEYINPUT80), .A3(new_n260), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n274), .A2(new_n266), .A3(new_n275), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n253), .A2(new_n265), .A3(new_n260), .ZN(new_n277));
  AND2_X1   g076(.A1(new_n277), .A2(new_n267), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n272), .A2(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(G8gat), .B(G36gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(G64gat), .B(G92gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n281), .B(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(KEYINPUT72), .B(KEYINPUT73), .ZN(new_n284));
  XOR2_X1   g083(.A(new_n283), .B(new_n284), .Z(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(G197gat), .B(G204gat), .ZN(new_n287));
  INV_X1    g086(.A(G211gat), .ZN(new_n288));
  INV_X1    g087(.A(G218gat), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n287), .B1(KEYINPUT22), .B2(new_n290), .ZN(new_n291));
  XOR2_X1   g090(.A(G211gat), .B(G218gat), .Z(new_n292));
  XNOR2_X1  g091(.A(new_n291), .B(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT71), .ZN(new_n294));
  NAND2_X1  g093(.A1(G226gat), .A2(G233gat), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(KEYINPUT27), .B(G183gat), .ZN(new_n297));
  INV_X1    g096(.A(G190gat), .ZN(new_n298));
  AND2_X1   g097(.A1(new_n298), .A2(KEYINPUT28), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n297), .A2(KEYINPUT68), .A3(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  AOI21_X1  g100(.A(KEYINPUT68), .B1(new_n297), .B2(new_n299), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  XOR2_X1   g102(.A(KEYINPUT67), .B(KEYINPUT28), .Z(new_n304));
  NOR2_X1   g103(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n305));
  INV_X1    g104(.A(G183gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(KEYINPUT66), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT66), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(G183gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n305), .B1(new_n310), .B2(KEYINPUT27), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n304), .B1(new_n311), .B2(G190gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n303), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(G169gat), .ZN(new_n314));
  INV_X1    g113(.A(G176gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT26), .ZN(new_n317));
  NAND2_X1  g116(.A1(G169gat), .A2(G176gat), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n316), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  NOR2_X1   g118(.A1(G169gat), .A2(G176gat), .ZN(new_n320));
  AOI22_X1  g119(.A1(new_n320), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT69), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n319), .A2(new_n321), .A3(KEYINPUT69), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n313), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(G183gat), .A2(G190gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(KEYINPUT24), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT24), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n330), .A2(G183gat), .A3(G190gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n306), .A2(new_n298), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n318), .A2(KEYINPUT23), .ZN(new_n334));
  AOI22_X1  g133(.A1(new_n332), .A2(new_n333), .B1(new_n316), .B2(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n314), .A2(new_n315), .A3(KEYINPUT23), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(KEYINPUT64), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT64), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n320), .A2(new_n338), .A3(KEYINPUT23), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(KEYINPUT25), .B1(new_n335), .B2(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n307), .A2(new_n309), .A3(new_n298), .ZN(new_n342));
  AND2_X1   g141(.A1(new_n342), .A2(new_n332), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n334), .A2(new_n316), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n344), .A2(KEYINPUT25), .A3(new_n336), .ZN(new_n345));
  OAI22_X1  g144(.A1(new_n341), .A2(KEYINPUT65), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n332), .A2(new_n333), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n340), .A2(new_n347), .A3(new_n344), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT25), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT65), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n327), .B1(new_n346), .B2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT29), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n296), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  AOI22_X1  g154(.A1(new_n303), .A2(new_n312), .B1(new_n324), .B2(new_n325), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n343), .A2(new_n345), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n357), .B1(new_n350), .B2(new_n351), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n341), .A2(KEYINPUT65), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n356), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n360), .A2(new_n295), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n294), .B1(new_n355), .B2(new_n361), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n295), .B1(new_n360), .B2(KEYINPUT29), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT71), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n293), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n293), .ZN(new_n366));
  NOR3_X1   g165(.A1(new_n355), .A2(new_n361), .A3(new_n366), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n286), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n296), .ZN(new_n369));
  AOI21_X1  g168(.A(KEYINPUT71), .B1(new_n363), .B2(new_n369), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n355), .A2(new_n294), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n366), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n367), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n372), .A2(new_n373), .A3(new_n285), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n368), .A2(new_n374), .A3(KEYINPUT30), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n365), .A2(new_n367), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT30), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n376), .A2(new_n377), .A3(new_n285), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n375), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT35), .ZN(new_n380));
  AND3_X1   g179(.A1(new_n280), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  XNOR2_X1  g180(.A(G78gat), .B(G106gat), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n382), .B(G22gat), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n293), .A2(KEYINPUT79), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n291), .A2(KEYINPUT79), .A3(new_n292), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(new_n354), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n249), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  AOI22_X1  g187(.A1(new_n388), .A2(new_n256), .B1(G228gat), .B2(G233gat), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n293), .B1(new_n258), .B2(new_n354), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n293), .A2(new_n354), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n242), .B1(new_n393), .B2(new_n249), .ZN(new_n394));
  OAI211_X1 g193(.A(G228gat), .B(G233gat), .C1(new_n390), .C2(new_n394), .ZN(new_n395));
  XNOR2_X1  g194(.A(KEYINPUT31), .B(G50gat), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n392), .A2(new_n395), .A3(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n397), .B1(new_n392), .B2(new_n395), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n384), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n400), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n402), .A2(new_n383), .A3(new_n398), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n353), .A2(new_n248), .ZN(new_n405));
  OAI211_X1 g204(.A(new_n327), .B(new_n229), .C1(new_n346), .C2(new_n352), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(G227gat), .A2(G233gat), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(KEYINPUT34), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT34), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n405), .A2(new_n411), .A3(new_n408), .A4(new_n406), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  XOR2_X1   g213(.A(G15gat), .B(G43gat), .Z(new_n415));
  XNOR2_X1  g214(.A(G71gat), .B(G99gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n415), .B(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n408), .B1(new_n405), .B2(new_n406), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n417), .B1(new_n418), .B2(KEYINPUT33), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT32), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  AOI221_X4 g221(.A(new_n420), .B1(KEYINPUT33), .B2(new_n417), .C1(new_n407), .C2(new_n409), .ZN(new_n423));
  OAI211_X1 g222(.A(KEYINPUT70), .B(new_n414), .C1(new_n422), .C2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT70), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n413), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n407), .A2(new_n409), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(KEYINPUT32), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT33), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n428), .A2(new_n430), .A3(new_n417), .ZN(new_n431));
  INV_X1    g230(.A(new_n423), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n410), .A2(KEYINPUT70), .A3(new_n412), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n426), .A2(new_n431), .A3(new_n432), .A4(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n404), .B1(new_n424), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n381), .A2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n270), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n278), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n270), .A2(new_n268), .ZN(new_n439));
  AOI22_X1  g238(.A1(new_n375), .A2(new_n378), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n435), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(KEYINPUT35), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n436), .A2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT39), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n252), .A2(new_n444), .A3(new_n203), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n202), .B1(new_n254), .B2(new_n259), .ZN(new_n446));
  OR2_X1    g245(.A1(new_n241), .A2(new_n243), .ZN(new_n447));
  OAI21_X1  g246(.A(KEYINPUT39), .B1(new_n447), .B2(new_n203), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n265), .B(new_n445), .C1(new_n446), .C2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT40), .ZN(new_n450));
  OAI21_X1  g249(.A(KEYINPUT81), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  OR2_X1    g250(.A1(new_n446), .A2(new_n448), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT81), .ZN(new_n453));
  AND2_X1   g252(.A1(new_n445), .A2(new_n265), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n452), .A2(new_n453), .A3(KEYINPUT40), .A4(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n451), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n265), .B1(new_n261), .B2(new_n273), .ZN(new_n457));
  AOI22_X1  g256(.A1(new_n457), .A2(new_n275), .B1(new_n450), .B2(new_n449), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n375), .A2(new_n378), .A3(new_n456), .A4(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n404), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n293), .B1(new_n370), .B2(new_n371), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT37), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n355), .A2(new_n361), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n462), .B1(new_n463), .B2(new_n366), .ZN(new_n464));
  AOI21_X1  g263(.A(KEYINPUT38), .B1(new_n461), .B2(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n285), .B1(new_n372), .B2(new_n373), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n285), .A2(new_n462), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n468), .A2(new_n272), .A3(new_n374), .A4(new_n279), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT38), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n285), .B1(new_n376), .B2(new_n462), .ZN(new_n471));
  OAI21_X1  g270(.A(KEYINPUT37), .B1(new_n365), .B2(new_n367), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  OAI211_X1 g272(.A(new_n459), .B(new_n460), .C1(new_n469), .C2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n434), .A2(new_n424), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT36), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n434), .A2(new_n424), .A3(KEYINPUT36), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n478), .B(new_n479), .C1(new_n440), .C2(new_n460), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n443), .B1(new_n475), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g280(.A1(G71gat), .A2(G78gat), .ZN(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT94), .ZN(new_n484));
  NAND2_X1  g283(.A1(G71gat), .A2(G78gat), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n485), .ZN(new_n487));
  OAI21_X1  g286(.A(KEYINPUT94), .B1(new_n487), .B2(new_n482), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(G57gat), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(G64gat), .ZN(new_n491));
  INV_X1    g290(.A(G64gat), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(G57gat), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT9), .ZN(new_n494));
  AOI22_X1  g293(.A1(new_n491), .A2(new_n493), .B1(new_n494), .B2(new_n485), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n489), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n491), .A2(new_n493), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n485), .A2(new_n494), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OR2_X1    g298(.A1(new_n485), .A2(KEYINPUT93), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n482), .B1(KEYINPUT93), .B2(new_n485), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n496), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT21), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(G231gat), .A2(G233gat), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n505), .B(new_n506), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n507), .B(KEYINPUT20), .ZN(new_n508));
  INV_X1    g307(.A(G1gat), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(KEYINPUT16), .ZN(new_n510));
  XNOR2_X1  g309(.A(G15gat), .B(G22gat), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT89), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(G22gat), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(G15gat), .ZN(new_n515));
  INV_X1    g314(.A(G15gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(G22gat), .ZN(new_n517));
  AND3_X1   g316(.A1(new_n515), .A2(new_n517), .A3(new_n512), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n510), .B1(new_n513), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n515), .A2(new_n517), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(KEYINPUT89), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n511), .A2(new_n512), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n521), .A2(new_n522), .A3(new_n509), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(G8gat), .ZN(new_n525));
  INV_X1    g324(.A(G8gat), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n519), .A2(new_n526), .A3(new_n523), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n529), .B1(new_n504), .B2(new_n503), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n508), .B(new_n530), .ZN(new_n531));
  XOR2_X1   g330(.A(KEYINPUT95), .B(KEYINPUT19), .Z(new_n532));
  XNOR2_X1  g331(.A(new_n532), .B(KEYINPUT96), .ZN(new_n533));
  XOR2_X1   g332(.A(G127gat), .B(G155gat), .Z(new_n534));
  XNOR2_X1  g333(.A(new_n533), .B(new_n534), .ZN(new_n535));
  XOR2_X1   g334(.A(G183gat), .B(G211gat), .Z(new_n536));
  XNOR2_X1  g335(.A(new_n535), .B(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n531), .B(new_n537), .ZN(new_n538));
  AND2_X1   g337(.A1(G232gat), .A2(G233gat), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n539), .A2(KEYINPUT41), .ZN(new_n540));
  XNOR2_X1  g339(.A(G134gat), .B(G162gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n540), .B(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT88), .ZN(new_n544));
  XNOR2_X1  g343(.A(G43gat), .B(G50gat), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT84), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(G43gat), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n548), .A2(G50gat), .ZN(new_n549));
  INV_X1    g348(.A(G50gat), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n550), .A2(G43gat), .ZN(new_n551));
  OAI21_X1  g350(.A(KEYINPUT84), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n547), .A2(new_n552), .A3(KEYINPUT15), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT15), .ZN(new_n554));
  OR2_X1    g353(.A1(KEYINPUT87), .A2(G50gat), .ZN(new_n555));
  NAND2_X1  g354(.A1(KEYINPUT87), .A2(G50gat), .ZN(new_n556));
  AOI21_X1  g355(.A(G43gat), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n554), .B1(new_n557), .B2(new_n549), .ZN(new_n558));
  INV_X1    g357(.A(G29gat), .ZN(new_n559));
  INV_X1    g358(.A(G36gat), .ZN(new_n560));
  OAI21_X1  g359(.A(KEYINPUT86), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT86), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n562), .A2(G29gat), .A3(G36gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n559), .A2(new_n560), .A3(KEYINPUT14), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT14), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n566), .B1(G29gat), .B2(G36gat), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n564), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n553), .A2(new_n558), .A3(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT85), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n564), .B1(new_n572), .B2(new_n568), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n565), .A2(new_n567), .A3(KEYINPUT85), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n553), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n544), .B1(new_n571), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n573), .A2(new_n574), .ZN(new_n577));
  INV_X1    g376(.A(new_n553), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n579), .A2(KEYINPUT88), .A3(new_n570), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT17), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n576), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n579), .A2(KEYINPUT17), .A3(new_n570), .ZN(new_n583));
  NAND2_X1  g382(.A1(G99gat), .A2(G106gat), .ZN(new_n584));
  INV_X1    g383(.A(G85gat), .ZN(new_n585));
  INV_X1    g384(.A(G92gat), .ZN(new_n586));
  AOI22_X1  g385(.A1(KEYINPUT8), .A2(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(G85gat), .A2(G92gat), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT7), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n587), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(G99gat), .B(G106gat), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  AND2_X1   g394(.A1(new_n590), .A2(new_n591), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n596), .A2(new_n593), .A3(new_n587), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n582), .A2(new_n583), .A3(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n539), .A2(KEYINPUT41), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n576), .A2(new_n580), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n601), .B1(new_n602), .B2(new_n598), .ZN(new_n603));
  XOR2_X1   g402(.A(G190gat), .B(G218gat), .Z(new_n604));
  NOR3_X1   g403(.A1(new_n600), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n604), .ZN(new_n606));
  INV_X1    g405(.A(new_n603), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n606), .B1(new_n607), .B2(new_n599), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n543), .B1(new_n605), .B2(new_n608), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n604), .B1(new_n600), .B2(new_n603), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n607), .A2(new_n606), .A3(new_n599), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n610), .A2(new_n611), .A3(new_n542), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n538), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n503), .A2(new_n598), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT10), .ZN(new_n617));
  NAND4_X1  g416(.A1(new_n496), .A2(new_n595), .A3(new_n502), .A4(new_n597), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  AND2_X1   g418(.A1(new_n496), .A2(new_n502), .ZN(new_n620));
  AND2_X1   g419(.A1(new_n595), .A2(new_n597), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT97), .ZN(new_n622));
  NAND4_X1  g421(.A1(new_n620), .A2(new_n621), .A3(new_n622), .A4(KEYINPUT10), .ZN(new_n623));
  OAI21_X1  g422(.A(KEYINPUT97), .B1(new_n618), .B2(new_n617), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n619), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(G230gat), .A2(G233gat), .ZN(new_n626));
  XOR2_X1   g425(.A(new_n626), .B(KEYINPUT98), .Z(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT101), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n625), .A2(KEYINPUT101), .A3(new_n628), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n616), .A2(new_n618), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(new_n627), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  XOR2_X1   g435(.A(G120gat), .B(G148gat), .Z(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(KEYINPUT99), .ZN(new_n638));
  XNOR2_X1  g437(.A(G176gat), .B(G204gat), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n638), .B(new_n639), .Z(new_n640));
  XOR2_X1   g439(.A(new_n640), .B(KEYINPUT100), .Z(new_n641));
  NAND2_X1  g440(.A1(new_n636), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n640), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n629), .A2(new_n635), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n615), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(G113gat), .B(G141gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(KEYINPUT83), .B(G197gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(KEYINPUT11), .B(G169gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(KEYINPUT12), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n582), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT90), .ZN(new_n656));
  INV_X1    g455(.A(new_n527), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n526), .B1(new_n519), .B2(new_n523), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n656), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n525), .A2(KEYINPUT90), .A3(new_n527), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n659), .A2(new_n660), .A3(new_n583), .ZN(new_n661));
  OAI21_X1  g460(.A(KEYINPUT91), .B1(new_n655), .B2(new_n661), .ZN(new_n662));
  AND2_X1   g461(.A1(new_n659), .A2(new_n660), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT91), .ZN(new_n664));
  NAND4_X1  g463(.A1(new_n663), .A2(new_n582), .A3(new_n664), .A4(new_n583), .ZN(new_n665));
  NAND2_X1  g464(.A1(G229gat), .A2(G233gat), .ZN(new_n666));
  NOR3_X1   g465(.A1(new_n571), .A2(new_n575), .A3(new_n544), .ZN(new_n667));
  AOI21_X1  g466(.A(KEYINPUT88), .B1(new_n579), .B2(new_n570), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(new_n528), .ZN(new_n670));
  NAND4_X1  g469(.A1(new_n662), .A2(new_n665), .A3(new_n666), .A4(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT18), .ZN(new_n672));
  AND2_X1   g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n602), .A2(new_n529), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n670), .A2(new_n674), .ZN(new_n675));
  XOR2_X1   g474(.A(new_n666), .B(KEYINPUT13), .Z(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n677), .B1(new_n671), .B2(new_n672), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n654), .B1(new_n673), .B2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT92), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n680), .B1(new_n671), .B2(new_n672), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n671), .A2(new_n680), .A3(new_n672), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  OAI211_X1 g483(.A(new_n677), .B(new_n653), .C1(new_n671), .C2(new_n672), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n679), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n647), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n481), .A2(new_n688), .ZN(new_n689));
  OR2_X1    g488(.A1(new_n689), .A2(KEYINPUT102), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(KEYINPUT102), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n438), .A2(new_n439), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(G1gat), .ZN(G1324gat));
  INV_X1    g495(.A(new_n379), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n526), .B1(new_n692), .B2(new_n697), .ZN(new_n698));
  XNOR2_X1  g497(.A(KEYINPUT104), .B(KEYINPUT16), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(new_n526), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n692), .A2(new_n697), .A3(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n698), .B1(new_n702), .B2(KEYINPUT42), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT105), .ZN(new_n704));
  XNOR2_X1  g503(.A(KEYINPUT103), .B(KEYINPUT42), .ZN(new_n705));
  AND3_X1   g504(.A1(new_n701), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n704), .B1(new_n701), .B2(new_n705), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n703), .B1(new_n706), .B2(new_n707), .ZN(G1325gat));
  NAND3_X1  g507(.A1(new_n692), .A2(new_n516), .A3(new_n476), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n478), .A2(new_n479), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n711), .B1(new_n690), .B2(new_n691), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n709), .B1(new_n516), .B2(new_n712), .ZN(G1326gat));
  NAND2_X1  g512(.A1(new_n692), .A2(new_n404), .ZN(new_n714));
  XNOR2_X1  g513(.A(KEYINPUT43), .B(G22gat), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n714), .B(new_n715), .ZN(G1327gat));
  INV_X1    g515(.A(KEYINPUT44), .ZN(new_n717));
  AOI22_X1  g516(.A1(new_n435), .A2(new_n381), .B1(new_n441), .B2(KEYINPUT35), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT106), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n719), .B1(new_n475), .B2(new_n480), .ZN(new_n720));
  INV_X1    g519(.A(new_n480), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n721), .A2(KEYINPUT106), .A3(new_n474), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n718), .B1(new_n720), .B2(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n717), .B1(new_n723), .B2(new_n613), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n481), .A2(KEYINPUT44), .A3(new_n614), .ZN(new_n725));
  AND2_X1   g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n538), .ZN(new_n727));
  NOR3_X1   g526(.A1(new_n687), .A2(new_n727), .A3(new_n645), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n726), .A2(new_n694), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(KEYINPUT107), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT107), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n726), .A2(new_n731), .A3(new_n694), .A4(new_n728), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n730), .A2(G29gat), .A3(new_n732), .ZN(new_n733));
  AND3_X1   g532(.A1(new_n481), .A2(new_n614), .A3(new_n728), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n734), .A2(new_n559), .A3(new_n694), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(KEYINPUT45), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n733), .A2(new_n736), .ZN(G1328gat));
  NAND2_X1  g536(.A1(new_n726), .A2(new_n728), .ZN(new_n738));
  OAI21_X1  g537(.A(G36gat), .B1(new_n738), .B2(new_n379), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n734), .A2(new_n560), .A3(new_n697), .ZN(new_n740));
  XOR2_X1   g539(.A(new_n740), .B(KEYINPUT46), .Z(new_n741));
  NAND2_X1  g540(.A1(new_n739), .A2(new_n741), .ZN(G1329gat));
  NAND2_X1  g541(.A1(new_n734), .A2(new_n476), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(new_n548), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n711), .A2(new_n548), .ZN(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n744), .B1(new_n738), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(KEYINPUT47), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT47), .ZN(new_n749));
  OAI211_X1 g548(.A(new_n744), .B(new_n749), .C1(new_n738), .C2(new_n746), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n748), .A2(new_n750), .ZN(G1330gat));
  NAND4_X1  g550(.A1(new_n724), .A2(new_n404), .A3(new_n728), .A4(new_n725), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n555), .A2(new_n556), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT108), .ZN(new_n755));
  AOI21_X1  g554(.A(KEYINPUT48), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n734), .A2(new_n404), .A3(new_n555), .A4(new_n556), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n754), .B(new_n757), .C1(new_n755), .C2(KEYINPUT48), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(G1331gat));
  NOR3_X1   g560(.A1(new_n475), .A2(new_n719), .A3(new_n480), .ZN(new_n762));
  AOI21_X1  g561(.A(KEYINPUT106), .B1(new_n721), .B2(new_n474), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n443), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n615), .A2(new_n645), .ZN(new_n765));
  INV_X1    g564(.A(new_n765), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n764), .A2(KEYINPUT109), .A3(new_n687), .A4(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT109), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n766), .A2(new_n687), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n768), .B1(new_n723), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n767), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n771), .A2(new_n693), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(new_n490), .ZN(G1332gat));
  AOI21_X1  g572(.A(new_n379), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n767), .A2(new_n770), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(KEYINPUT110), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT110), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n767), .A2(new_n770), .A3(new_n777), .A4(new_n774), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g578(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n779), .B(new_n780), .ZN(G1333gat));
  OAI21_X1  g580(.A(G71gat), .B1(new_n771), .B2(new_n711), .ZN(new_n782));
  INV_X1    g581(.A(G71gat), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n476), .A2(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n782), .B1(new_n771), .B2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT50), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  OAI211_X1 g586(.A(new_n782), .B(KEYINPUT50), .C1(new_n771), .C2(new_n784), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(G1334gat));
  NOR2_X1   g588(.A1(new_n771), .A2(new_n460), .ZN(new_n790));
  XOR2_X1   g589(.A(KEYINPUT111), .B(G78gat), .Z(new_n791));
  XNOR2_X1  g590(.A(new_n790), .B(new_n791), .ZN(G1335gat));
  NOR2_X1   g591(.A1(new_n727), .A2(new_n686), .ZN(new_n793));
  INV_X1    g592(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n794), .A2(new_n646), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n726), .A2(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(G85gat), .B1(new_n796), .B2(new_n693), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n720), .A2(new_n722), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n613), .B1(new_n798), .B2(new_n443), .ZN(new_n799));
  AOI21_X1  g598(.A(KEYINPUT51), .B1(new_n799), .B2(new_n793), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT51), .ZN(new_n801));
  NOR4_X1   g600(.A1(new_n723), .A2(new_n801), .A3(new_n613), .A4(new_n794), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n694), .A2(new_n585), .A3(new_n645), .ZN(new_n804));
  XNOR2_X1  g603(.A(new_n804), .B(KEYINPUT112), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n797), .B1(new_n803), .B2(new_n805), .ZN(G1336gat));
  NAND4_X1  g605(.A1(new_n724), .A2(new_n697), .A3(new_n725), .A4(new_n795), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(G92gat), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n379), .A2(G92gat), .A3(new_n646), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n809), .B(KEYINPUT113), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n808), .B1(new_n803), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(KEYINPUT52), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT52), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n808), .B(new_n813), .C1(new_n803), .C2(new_n810), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n812), .A2(new_n814), .ZN(G1337gat));
  OAI21_X1  g614(.A(G99gat), .B1(new_n796), .B2(new_n711), .ZN(new_n816));
  INV_X1    g615(.A(G99gat), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n476), .A2(new_n817), .A3(new_n645), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n816), .B1(new_n803), .B2(new_n818), .ZN(G1338gat));
  INV_X1    g618(.A(KEYINPUT115), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n820), .A2(KEYINPUT53), .ZN(new_n821));
  AND2_X1   g620(.A1(new_n820), .A2(KEYINPUT53), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n460), .A2(new_n646), .A3(G106gat), .ZN(new_n823));
  XNOR2_X1  g622(.A(new_n823), .B(KEYINPUT114), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n824), .B1(new_n800), .B2(new_n802), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n724), .A2(new_n404), .A3(new_n725), .A4(new_n795), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(G106gat), .ZN(new_n827));
  AOI211_X1 g626(.A(new_n821), .B(new_n822), .C1(new_n825), .C2(new_n827), .ZN(new_n828));
  AND4_X1   g627(.A1(new_n820), .A2(new_n825), .A3(new_n827), .A4(KEYINPUT53), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n828), .A2(new_n829), .ZN(G1339gat));
  INV_X1    g629(.A(KEYINPUT54), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n631), .A2(new_n831), .A3(new_n632), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT55), .ZN(new_n833));
  OR2_X1    g632(.A1(new_n625), .A2(new_n628), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n831), .B1(new_n625), .B2(new_n628), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n833), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n832), .A2(new_n836), .A3(new_n640), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(KEYINPUT116), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT116), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n832), .A2(new_n836), .A3(new_n839), .A4(new_n640), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n644), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(KEYINPUT117), .ZN(new_n843));
  INV_X1    g642(.A(new_n644), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n844), .B1(new_n838), .B2(new_n840), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT117), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n834), .A2(new_n835), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n832), .A2(new_n640), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(new_n833), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n843), .A2(new_n686), .A3(new_n847), .A4(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(new_n652), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n662), .A2(new_n665), .A3(new_n670), .ZN(new_n853));
  INV_X1    g652(.A(new_n666), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  OR2_X1    g654(.A1(new_n675), .A2(new_n676), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n852), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  AND3_X1   g656(.A1(new_n671), .A2(new_n680), .A3(new_n672), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n858), .A2(new_n681), .ZN(new_n859));
  INV_X1    g658(.A(new_n685), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n857), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n645), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n614), .B1(new_n851), .B2(new_n862), .ZN(new_n863));
  AOI22_X1  g662(.A1(new_n842), .A2(KEYINPUT117), .B1(new_n833), .B2(new_n849), .ZN(new_n864));
  AOI211_X1 g663(.A(new_n857), .B(new_n613), .C1(new_n859), .C2(new_n860), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n864), .A2(new_n865), .A3(new_n847), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n538), .B1(new_n863), .B2(new_n867), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n647), .A2(new_n686), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n404), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n871), .A2(new_n694), .A3(new_n379), .A4(new_n476), .ZN(new_n872));
  OAI21_X1  g671(.A(G113gat), .B1(new_n872), .B2(new_n687), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n693), .B1(new_n868), .B2(new_n870), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n874), .A2(new_n379), .A3(new_n435), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n687), .A2(G113gat), .ZN(new_n876));
  XOR2_X1   g675(.A(new_n876), .B(KEYINPUT118), .Z(new_n877));
  OAI21_X1  g676(.A(new_n873), .B1(new_n875), .B2(new_n877), .ZN(G1340gat));
  INV_X1    g677(.A(G120gat), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n872), .A2(new_n879), .A3(new_n646), .ZN(new_n880));
  OR2_X1    g679(.A1(new_n875), .A2(new_n646), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n880), .B1(new_n879), .B2(new_n881), .ZN(G1341gat));
  OAI21_X1  g681(.A(G127gat), .B1(new_n872), .B2(new_n538), .ZN(new_n883));
  OR2_X1    g682(.A1(new_n538), .A2(G127gat), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n883), .B1(new_n875), .B2(new_n884), .ZN(new_n885));
  XNOR2_X1  g684(.A(new_n885), .B(KEYINPUT119), .ZN(G1342gat));
  NAND2_X1  g685(.A1(new_n379), .A2(new_n614), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n887), .A2(G134gat), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n874), .A2(new_n435), .A3(new_n888), .ZN(new_n889));
  OR2_X1    g688(.A1(new_n889), .A2(KEYINPUT56), .ZN(new_n890));
  OAI21_X1  g689(.A(G134gat), .B1(new_n872), .B2(new_n613), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n889), .A2(KEYINPUT56), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(G1343gat));
  NOR2_X1   g692(.A1(KEYINPUT121), .A2(KEYINPUT58), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n710), .A2(new_n460), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n874), .A2(new_n379), .A3(new_n686), .A4(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n894), .B1(new_n896), .B2(new_n206), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n710), .A2(new_n693), .A3(new_n697), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n868), .A2(new_n870), .ZN(new_n899));
  AOI21_X1  g698(.A(KEYINPUT57), .B1(new_n899), .B2(new_n404), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT120), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n849), .A2(new_n901), .ZN(new_n902));
  NAND4_X1  g701(.A1(new_n832), .A2(KEYINPUT120), .A3(new_n640), .A4(new_n848), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n902), .A2(new_n833), .A3(new_n903), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n845), .A2(new_n904), .ZN(new_n905));
  AOI22_X1  g704(.A1(new_n905), .A2(new_n686), .B1(new_n861), .B2(new_n645), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n866), .B1(new_n906), .B2(new_n614), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n869), .B1(new_n907), .B2(new_n538), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT57), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n908), .A2(new_n909), .A3(new_n460), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n898), .B1(new_n900), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n686), .A2(G141gat), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n897), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(KEYINPUT121), .A2(KEYINPUT58), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n913), .B(new_n914), .ZN(G1344gat));
  NAND2_X1  g714(.A1(new_n898), .A2(new_n645), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n727), .B1(new_n907), .B2(KEYINPUT123), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT123), .ZN(new_n918));
  OAI211_X1 g717(.A(new_n866), .B(new_n918), .C1(new_n906), .C2(new_n614), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n869), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n909), .B1(new_n920), .B2(new_n460), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n899), .A2(KEYINPUT57), .A3(new_n404), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n916), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(KEYINPUT59), .B1(new_n923), .B2(new_n207), .ZN(new_n924));
  OAI211_X1 g723(.A(new_n645), .B(new_n898), .C1(new_n900), .C2(new_n910), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n207), .A2(KEYINPUT59), .ZN(new_n926));
  AND3_X1   g725(.A1(new_n925), .A2(KEYINPUT122), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g726(.A(KEYINPUT122), .B1(new_n925), .B2(new_n926), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n924), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n874), .A2(new_n895), .ZN(new_n930));
  OR4_X1    g729(.A1(G148gat), .A2(new_n930), .A3(new_n697), .A4(new_n646), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n929), .A2(new_n931), .ZN(G1345gat));
  INV_X1    g731(.A(G155gat), .ZN(new_n933));
  NOR3_X1   g732(.A1(new_n911), .A2(new_n933), .A3(new_n538), .ZN(new_n934));
  NOR3_X1   g733(.A1(new_n930), .A2(new_n697), .A3(new_n538), .ZN(new_n935));
  OR2_X1    g734(.A1(new_n935), .A2(KEYINPUT124), .ZN(new_n936));
  AOI21_X1  g735(.A(G155gat), .B1(new_n935), .B2(KEYINPUT124), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n934), .B1(new_n936), .B2(new_n937), .ZN(G1346gat));
  OAI21_X1  g737(.A(G162gat), .B1(new_n911), .B2(new_n613), .ZN(new_n939));
  OR2_X1    g738(.A1(new_n887), .A2(G162gat), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n939), .B1(new_n930), .B2(new_n940), .ZN(G1347gat));
  AND3_X1   g740(.A1(new_n697), .A2(new_n693), .A3(new_n476), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n871), .A2(new_n942), .ZN(new_n943));
  NOR3_X1   g742(.A1(new_n943), .A2(new_n314), .A3(new_n687), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n694), .B1(new_n868), .B2(new_n870), .ZN(new_n945));
  AND3_X1   g744(.A1(new_n945), .A2(new_n697), .A3(new_n435), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(new_n686), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n944), .B1(new_n314), .B2(new_n947), .ZN(G1348gat));
  NAND3_X1  g747(.A1(new_n946), .A2(new_n315), .A3(new_n645), .ZN(new_n949));
  OAI21_X1  g748(.A(G176gat), .B1(new_n943), .B2(new_n646), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(G1349gat));
  NAND2_X1  g750(.A1(new_n727), .A2(new_n297), .ZN(new_n952));
  INV_X1    g751(.A(new_n952), .ZN(new_n953));
  AOI22_X1  g752(.A1(new_n946), .A2(new_n953), .B1(KEYINPUT125), .B2(KEYINPUT60), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n310), .B1(new_n943), .B2(new_n538), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g755(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n957));
  INV_X1    g756(.A(new_n957), .ZN(new_n958));
  XNOR2_X1  g757(.A(new_n956), .B(new_n958), .ZN(G1350gat));
  NAND3_X1  g758(.A1(new_n946), .A2(new_n298), .A3(new_n614), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n871), .A2(new_n614), .A3(new_n942), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT61), .ZN(new_n962));
  AND3_X1   g761(.A1(new_n961), .A2(new_n962), .A3(G190gat), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n962), .B1(new_n961), .B2(G190gat), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n960), .B1(new_n963), .B2(new_n964), .ZN(G1351gat));
  NAND2_X1  g764(.A1(new_n907), .A2(KEYINPUT123), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n966), .A2(new_n538), .A3(new_n919), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n460), .B1(new_n967), .B2(new_n870), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n922), .B1(new_n968), .B2(KEYINPUT57), .ZN(new_n969));
  NOR3_X1   g768(.A1(new_n710), .A2(new_n694), .A3(new_n379), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n969), .A2(new_n686), .A3(new_n970), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT126), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND4_X1  g772(.A1(new_n969), .A2(KEYINPUT126), .A3(new_n686), .A4(new_n970), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n973), .A2(G197gat), .A3(new_n974), .ZN(new_n975));
  NOR3_X1   g774(.A1(new_n710), .A2(new_n379), .A3(new_n460), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n945), .A2(new_n976), .ZN(new_n977));
  OR3_X1    g776(.A1(new_n977), .A2(G197gat), .A3(new_n687), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n975), .A2(new_n978), .ZN(G1352gat));
  INV_X1    g778(.A(G204gat), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n645), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g780(.A(KEYINPUT62), .B1(new_n977), .B2(new_n981), .ZN(new_n982));
  OR3_X1    g781(.A1(new_n977), .A2(KEYINPUT62), .A3(new_n981), .ZN(new_n983));
  AND3_X1   g782(.A1(new_n969), .A2(new_n645), .A3(new_n970), .ZN(new_n984));
  OAI211_X1 g783(.A(new_n982), .B(new_n983), .C1(new_n984), .C2(new_n980), .ZN(G1353gat));
  INV_X1    g784(.A(new_n977), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n986), .A2(new_n288), .A3(new_n727), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n969), .A2(new_n727), .A3(new_n970), .ZN(new_n988));
  INV_X1    g787(.A(KEYINPUT63), .ZN(new_n989));
  AOI21_X1  g788(.A(new_n288), .B1(KEYINPUT127), .B2(new_n989), .ZN(new_n990));
  NOR2_X1   g789(.A1(new_n989), .A2(KEYINPUT127), .ZN(new_n991));
  AND3_X1   g790(.A1(new_n988), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  AOI21_X1  g791(.A(new_n991), .B1(new_n988), .B2(new_n990), .ZN(new_n993));
  OAI21_X1  g792(.A(new_n987), .B1(new_n992), .B2(new_n993), .ZN(G1354gat));
  NAND3_X1  g793(.A1(new_n986), .A2(new_n289), .A3(new_n614), .ZN(new_n995));
  AND3_X1   g794(.A1(new_n969), .A2(new_n614), .A3(new_n970), .ZN(new_n996));
  OAI21_X1  g795(.A(new_n995), .B1(new_n996), .B2(new_n289), .ZN(G1355gat));
endmodule


