

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U553 ( .A1(n574), .A2(n547), .ZN(n801) );
  XOR2_X1 U554 ( .A(KEYINPUT1), .B(n548), .Z(n798) );
  NOR2_X2 U555 ( .A1(n605), .A2(n604), .ZN(n928) );
  NOR2_X4 U556 ( .A1(n540), .A2(n539), .ZN(G160) );
  NOR2_X1 U557 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X2 U558 ( .A(n594), .B(n593), .ZN(n728) );
  NAND2_X2 U559 ( .A1(n729), .A2(n595), .ZN(n651) );
  XNOR2_X1 U560 ( .A(n522), .B(n521), .ZN(n534) );
  NOR2_X1 U561 ( .A1(G2105), .A2(G2104), .ZN(n521) );
  XNOR2_X1 U562 ( .A(n533), .B(n532), .ZN(n536) );
  XNOR2_X1 U563 ( .A(n531), .B(KEYINPUT66), .ZN(n532) );
  INV_X1 U564 ( .A(KEYINPUT23), .ZN(n531) );
  INV_X1 U565 ( .A(KEYINPUT29), .ZN(n642) );
  AND2_X1 U566 ( .A1(n708), .A2(n707), .ZN(n520) );
  INV_X1 U567 ( .A(KEYINPUT97), .ZN(n622) );
  NOR2_X1 U568 ( .A1(n635), .A2(n634), .ZN(n638) );
  INV_X1 U569 ( .A(n651), .ZN(n644) );
  XNOR2_X1 U570 ( .A(n654), .B(KEYINPUT100), .ZN(n655) );
  XNOR2_X1 U571 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U572 ( .A(n643), .B(n642), .ZN(n649) );
  XNOR2_X1 U573 ( .A(n652), .B(KEYINPUT92), .ZN(n663) );
  INV_X1 U574 ( .A(n752), .ZN(n741) );
  INV_X1 U575 ( .A(G2105), .ZN(n526) );
  NOR2_X1 U576 ( .A1(G651), .A2(n574), .ZN(n800) );
  NOR2_X2 U577 ( .A1(G2104), .A2(n526), .ZN(n896) );
  XNOR2_X1 U578 ( .A(KEYINPUT67), .B(KEYINPUT17), .ZN(n522) );
  BUF_X2 U579 ( .A(n534), .Z(n892) );
  NAND2_X1 U580 ( .A1(G138), .A2(n892), .ZN(n525) );
  INV_X1 U581 ( .A(G2105), .ZN(n523) );
  AND2_X4 U582 ( .A1(n523), .A2(G2104), .ZN(n893) );
  NAND2_X1 U583 ( .A1(G102), .A2(n893), .ZN(n524) );
  NAND2_X1 U584 ( .A1(n525), .A2(n524), .ZN(n530) );
  NAND2_X1 U585 ( .A1(G126), .A2(n896), .ZN(n528) );
  AND2_X1 U586 ( .A1(G2104), .A2(G2105), .ZN(n897) );
  NAND2_X1 U587 ( .A1(G114), .A2(n897), .ZN(n527) );
  NAND2_X1 U588 ( .A1(n528), .A2(n527), .ZN(n529) );
  NOR2_X1 U589 ( .A1(n530), .A2(n529), .ZN(G164) );
  NAND2_X1 U590 ( .A1(G101), .A2(n893), .ZN(n533) );
  NAND2_X1 U591 ( .A1(G137), .A2(n534), .ZN(n535) );
  NAND2_X1 U592 ( .A1(n536), .A2(n535), .ZN(n540) );
  NAND2_X1 U593 ( .A1(G125), .A2(n896), .ZN(n538) );
  NAND2_X1 U594 ( .A1(G113), .A2(n897), .ZN(n537) );
  NAND2_X1 U595 ( .A1(n538), .A2(n537), .ZN(n539) );
  NOR2_X1 U596 ( .A1(G543), .A2(G651), .ZN(n541) );
  XOR2_X2 U597 ( .A(KEYINPUT65), .B(n541), .Z(n804) );
  NAND2_X1 U598 ( .A1(G90), .A2(n804), .ZN(n543) );
  XOR2_X1 U599 ( .A(G543), .B(KEYINPUT0), .Z(n574) );
  INV_X1 U600 ( .A(G651), .ZN(n547) );
  NAND2_X1 U601 ( .A1(G77), .A2(n801), .ZN(n542) );
  NAND2_X1 U602 ( .A1(n543), .A2(n542), .ZN(n546) );
  XOR2_X1 U603 ( .A(KEYINPUT69), .B(KEYINPUT70), .Z(n544) );
  XNOR2_X1 U604 ( .A(KEYINPUT9), .B(n544), .ZN(n545) );
  XNOR2_X1 U605 ( .A(n546), .B(n545), .ZN(n552) );
  NAND2_X1 U606 ( .A1(G52), .A2(n800), .ZN(n550) );
  NOR2_X1 U607 ( .A1(G543), .A2(n547), .ZN(n548) );
  NAND2_X1 U608 ( .A1(G64), .A2(n798), .ZN(n549) );
  AND2_X1 U609 ( .A1(n550), .A2(n549), .ZN(n551) );
  NAND2_X1 U610 ( .A1(n552), .A2(n551), .ZN(G301) );
  INV_X1 U611 ( .A(G301), .ZN(G171) );
  NAND2_X1 U612 ( .A1(n804), .A2(G89), .ZN(n553) );
  XNOR2_X1 U613 ( .A(n553), .B(KEYINPUT4), .ZN(n555) );
  NAND2_X1 U614 ( .A1(G76), .A2(n801), .ZN(n554) );
  NAND2_X1 U615 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U616 ( .A(n556), .B(KEYINPUT5), .ZN(n561) );
  NAND2_X1 U617 ( .A1(G51), .A2(n800), .ZN(n558) );
  NAND2_X1 U618 ( .A1(G63), .A2(n798), .ZN(n557) );
  NAND2_X1 U619 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U620 ( .A(KEYINPUT6), .B(n559), .Z(n560) );
  NAND2_X1 U621 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U622 ( .A(n562), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U623 ( .A1(G50), .A2(n800), .ZN(n563) );
  XOR2_X1 U624 ( .A(KEYINPUT82), .B(n563), .Z(n568) );
  NAND2_X1 U625 ( .A1(G88), .A2(n804), .ZN(n565) );
  NAND2_X1 U626 ( .A1(G75), .A2(n801), .ZN(n564) );
  NAND2_X1 U627 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U628 ( .A(KEYINPUT83), .B(n566), .Z(n567) );
  NOR2_X1 U629 ( .A1(n568), .A2(n567), .ZN(n570) );
  NAND2_X1 U630 ( .A1(n798), .A2(G62), .ZN(n569) );
  NAND2_X1 U631 ( .A1(n570), .A2(n569), .ZN(G303) );
  XOR2_X1 U632 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U633 ( .A1(G49), .A2(n800), .ZN(n572) );
  NAND2_X1 U634 ( .A1(G74), .A2(G651), .ZN(n571) );
  NAND2_X1 U635 ( .A1(n572), .A2(n571), .ZN(n573) );
  NOR2_X1 U636 ( .A1(n798), .A2(n573), .ZN(n576) );
  NAND2_X1 U637 ( .A1(n574), .A2(G87), .ZN(n575) );
  NAND2_X1 U638 ( .A1(n576), .A2(n575), .ZN(G288) );
  NAND2_X1 U639 ( .A1(G73), .A2(n801), .ZN(n577) );
  XNOR2_X1 U640 ( .A(n577), .B(KEYINPUT2), .ZN(n584) );
  NAND2_X1 U641 ( .A1(G48), .A2(n800), .ZN(n579) );
  NAND2_X1 U642 ( .A1(G61), .A2(n798), .ZN(n578) );
  NAND2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n582) );
  NAND2_X1 U644 ( .A1(G86), .A2(n804), .ZN(n580) );
  XNOR2_X1 U645 ( .A(KEYINPUT81), .B(n580), .ZN(n581) );
  NOR2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n583) );
  NAND2_X1 U647 ( .A1(n584), .A2(n583), .ZN(G305) );
  NAND2_X1 U648 ( .A1(G85), .A2(n804), .ZN(n586) );
  NAND2_X1 U649 ( .A1(G72), .A2(n801), .ZN(n585) );
  NAND2_X1 U650 ( .A1(n586), .A2(n585), .ZN(n589) );
  NAND2_X1 U651 ( .A1(G47), .A2(n800), .ZN(n587) );
  XOR2_X1 U652 ( .A(KEYINPUT68), .B(n587), .Z(n588) );
  NOR2_X1 U653 ( .A1(n589), .A2(n588), .ZN(n591) );
  NAND2_X1 U654 ( .A1(n798), .A2(G60), .ZN(n590) );
  NAND2_X1 U655 ( .A1(n591), .A2(n590), .ZN(G290) );
  NOR2_X1 U656 ( .A1(G1384), .A2(G164), .ZN(n592) );
  XNOR2_X1 U657 ( .A(n592), .B(KEYINPUT64), .ZN(n729) );
  INV_X1 U658 ( .A(KEYINPUT85), .ZN(n594) );
  NAND2_X1 U659 ( .A1(G40), .A2(G160), .ZN(n593) );
  XNOR2_X1 U660 ( .A(n728), .B(KEYINPUT91), .ZN(n595) );
  NAND2_X1 U661 ( .A1(n651), .A2(G1341), .ZN(n596) );
  XNOR2_X1 U662 ( .A(n596), .B(KEYINPUT96), .ZN(n606) );
  NAND2_X1 U663 ( .A1(n804), .A2(G81), .ZN(n597) );
  XNOR2_X1 U664 ( .A(n597), .B(KEYINPUT12), .ZN(n599) );
  NAND2_X1 U665 ( .A1(G68), .A2(n801), .ZN(n598) );
  NAND2_X1 U666 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U667 ( .A(n600), .B(KEYINPUT13), .ZN(n602) );
  NAND2_X1 U668 ( .A1(G43), .A2(n800), .ZN(n601) );
  NAND2_X1 U669 ( .A1(n602), .A2(n601), .ZN(n605) );
  NAND2_X1 U670 ( .A1(n798), .A2(G56), .ZN(n603) );
  XOR2_X1 U671 ( .A(KEYINPUT14), .B(n603), .Z(n604) );
  NAND2_X1 U672 ( .A1(n606), .A2(n928), .ZN(n609) );
  XNOR2_X1 U673 ( .A(G1996), .B(KEYINPUT95), .ZN(n955) );
  NOR2_X1 U674 ( .A1(n651), .A2(n955), .ZN(n607) );
  XNOR2_X1 U675 ( .A(n607), .B(KEYINPUT26), .ZN(n608) );
  NOR2_X1 U676 ( .A1(n609), .A2(n608), .ZN(n624) );
  NAND2_X1 U677 ( .A1(G92), .A2(n804), .ZN(n611) );
  NAND2_X1 U678 ( .A1(G79), .A2(n801), .ZN(n610) );
  NAND2_X1 U679 ( .A1(n611), .A2(n610), .ZN(n615) );
  NAND2_X1 U680 ( .A1(G54), .A2(n800), .ZN(n613) );
  NAND2_X1 U681 ( .A1(G66), .A2(n798), .ZN(n612) );
  NAND2_X1 U682 ( .A1(n613), .A2(n612), .ZN(n614) );
  NOR2_X1 U683 ( .A1(n615), .A2(n614), .ZN(n617) );
  XNOR2_X1 U684 ( .A(KEYINPUT75), .B(KEYINPUT15), .ZN(n616) );
  XNOR2_X1 U685 ( .A(n617), .B(n616), .ZN(n912) );
  NAND2_X1 U686 ( .A1(n624), .A2(n912), .ZN(n621) );
  NOR2_X1 U687 ( .A1(n644), .A2(G1348), .ZN(n619) );
  NOR2_X1 U688 ( .A1(G2067), .A2(n651), .ZN(n618) );
  NOR2_X1 U689 ( .A1(n619), .A2(n618), .ZN(n620) );
  NAND2_X1 U690 ( .A1(n621), .A2(n620), .ZN(n623) );
  XNOR2_X1 U691 ( .A(n623), .B(n622), .ZN(n626) );
  OR2_X1 U692 ( .A1(n912), .A2(n624), .ZN(n625) );
  NAND2_X1 U693 ( .A1(n626), .A2(n625), .ZN(n637) );
  NAND2_X1 U694 ( .A1(G53), .A2(n800), .ZN(n628) );
  NAND2_X1 U695 ( .A1(G65), .A2(n798), .ZN(n627) );
  NAND2_X1 U696 ( .A1(n628), .A2(n627), .ZN(n632) );
  NAND2_X1 U697 ( .A1(G91), .A2(n804), .ZN(n630) );
  NAND2_X1 U698 ( .A1(G78), .A2(n801), .ZN(n629) );
  NAND2_X1 U699 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U700 ( .A1(n632), .A2(n631), .ZN(n936) );
  NAND2_X1 U701 ( .A1(n644), .A2(G2072), .ZN(n633) );
  XNOR2_X1 U702 ( .A(n633), .B(KEYINPUT27), .ZN(n635) );
  INV_X1 U703 ( .A(G1956), .ZN(n1004) );
  NOR2_X1 U704 ( .A1(n1004), .A2(n644), .ZN(n634) );
  NAND2_X1 U705 ( .A1(n936), .A2(n638), .ZN(n636) );
  NAND2_X1 U706 ( .A1(n637), .A2(n636), .ZN(n641) );
  NOR2_X1 U707 ( .A1(n936), .A2(n638), .ZN(n639) );
  XOR2_X1 U708 ( .A(n639), .B(KEYINPUT28), .Z(n640) );
  NAND2_X1 U709 ( .A1(n641), .A2(n640), .ZN(n643) );
  OR2_X1 U710 ( .A1(n644), .A2(G1961), .ZN(n646) );
  XNOR2_X1 U711 ( .A(KEYINPUT25), .B(G2078), .ZN(n956) );
  NAND2_X1 U712 ( .A1(n644), .A2(n956), .ZN(n645) );
  NAND2_X1 U713 ( .A1(n646), .A2(n645), .ZN(n658) );
  AND2_X1 U714 ( .A1(n658), .A2(G171), .ZN(n647) );
  XOR2_X1 U715 ( .A(KEYINPUT94), .B(n647), .Z(n648) );
  NAND2_X1 U716 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U717 ( .A(n650), .B(KEYINPUT98), .ZN(n676) );
  NAND2_X1 U718 ( .A1(n651), .A2(G8), .ZN(n652) );
  NOR2_X1 U719 ( .A1(n663), .A2(G1966), .ZN(n679) );
  NOR2_X1 U720 ( .A1(G2084), .A2(n651), .ZN(n680) );
  NOR2_X1 U721 ( .A1(n679), .A2(n680), .ZN(n653) );
  NAND2_X1 U722 ( .A1(G8), .A2(n653), .ZN(n656) );
  XOR2_X1 U723 ( .A(KEYINPUT30), .B(KEYINPUT99), .Z(n654) );
  NOR2_X1 U724 ( .A1(n657), .A2(G168), .ZN(n660) );
  NOR2_X1 U725 ( .A1(G171), .A2(n658), .ZN(n659) );
  NOR2_X1 U726 ( .A1(n660), .A2(n659), .ZN(n662) );
  INV_X1 U727 ( .A(KEYINPUT31), .ZN(n661) );
  XNOR2_X1 U728 ( .A(n662), .B(n661), .ZN(n677) );
  INV_X1 U729 ( .A(G8), .ZN(n668) );
  NOR2_X1 U730 ( .A1(n663), .A2(G1971), .ZN(n665) );
  NOR2_X1 U731 ( .A1(G2090), .A2(n651), .ZN(n664) );
  NOR2_X1 U732 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U733 ( .A1(n666), .A2(G303), .ZN(n667) );
  OR2_X1 U734 ( .A1(n668), .A2(n667), .ZN(n670) );
  AND2_X1 U735 ( .A1(n677), .A2(n670), .ZN(n669) );
  NAND2_X1 U736 ( .A1(n676), .A2(n669), .ZN(n674) );
  INV_X1 U737 ( .A(n670), .ZN(n672) );
  AND2_X1 U738 ( .A1(G286), .A2(G8), .ZN(n671) );
  OR2_X1 U739 ( .A1(n672), .A2(n671), .ZN(n673) );
  NAND2_X1 U740 ( .A1(n674), .A2(n673), .ZN(n675) );
  XNOR2_X1 U741 ( .A(n675), .B(KEYINPUT32), .ZN(n684) );
  AND2_X1 U742 ( .A1(n677), .A2(n676), .ZN(n678) );
  NOR2_X1 U743 ( .A1(n679), .A2(n678), .ZN(n682) );
  NAND2_X1 U744 ( .A1(G8), .A2(n680), .ZN(n681) );
  NAND2_X1 U745 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U746 ( .A1(n684), .A2(n683), .ZN(n703) );
  NOR2_X1 U747 ( .A1(G1976), .A2(G288), .ZN(n688) );
  NOR2_X1 U748 ( .A1(G1971), .A2(G303), .ZN(n685) );
  NOR2_X1 U749 ( .A1(n688), .A2(n685), .ZN(n926) );
  NAND2_X1 U750 ( .A1(n703), .A2(n926), .ZN(n686) );
  XNOR2_X1 U751 ( .A(KEYINPUT101), .B(n686), .ZN(n695) );
  NAND2_X1 U752 ( .A1(G1976), .A2(G288), .ZN(n937) );
  INV_X1 U753 ( .A(n663), .ZN(n687) );
  NAND2_X1 U754 ( .A1(n937), .A2(n687), .ZN(n693) );
  NAND2_X1 U755 ( .A1(n688), .A2(KEYINPUT33), .ZN(n689) );
  NOR2_X1 U756 ( .A1(n663), .A2(n689), .ZN(n691) );
  XOR2_X1 U757 ( .A(G1981), .B(G305), .Z(n929) );
  INV_X1 U758 ( .A(n929), .ZN(n690) );
  NOR2_X1 U759 ( .A1(n691), .A2(n690), .ZN(n696) );
  INV_X1 U760 ( .A(n696), .ZN(n692) );
  OR2_X1 U761 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U762 ( .A1(n695), .A2(n694), .ZN(n698) );
  AND2_X1 U763 ( .A1(n696), .A2(KEYINPUT33), .ZN(n697) );
  XNOR2_X1 U764 ( .A(n699), .B(KEYINPUT102), .ZN(n709) );
  NOR2_X1 U765 ( .A1(G1981), .A2(G305), .ZN(n700) );
  XOR2_X1 U766 ( .A(n700), .B(KEYINPUT24), .Z(n701) );
  NOR2_X1 U767 ( .A1(n663), .A2(n701), .ZN(n702) );
  XNOR2_X1 U768 ( .A(n702), .B(KEYINPUT93), .ZN(n708) );
  NOR2_X1 U769 ( .A1(G2090), .A2(G303), .ZN(n704) );
  NAND2_X1 U770 ( .A1(G8), .A2(n704), .ZN(n705) );
  NAND2_X1 U771 ( .A1(n703), .A2(n705), .ZN(n706) );
  NAND2_X1 U772 ( .A1(n663), .A2(n706), .ZN(n707) );
  NAND2_X1 U773 ( .A1(n709), .A2(n520), .ZN(n743) );
  NAND2_X1 U774 ( .A1(G141), .A2(n892), .ZN(n710) );
  XNOR2_X1 U775 ( .A(n710), .B(KEYINPUT88), .ZN(n717) );
  NAND2_X1 U776 ( .A1(G129), .A2(n896), .ZN(n712) );
  NAND2_X1 U777 ( .A1(G117), .A2(n897), .ZN(n711) );
  NAND2_X1 U778 ( .A1(n712), .A2(n711), .ZN(n715) );
  NAND2_X1 U779 ( .A1(n893), .A2(G105), .ZN(n713) );
  XOR2_X1 U780 ( .A(KEYINPUT38), .B(n713), .Z(n714) );
  NOR2_X1 U781 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U782 ( .A1(n717), .A2(n716), .ZN(n718) );
  XOR2_X1 U783 ( .A(KEYINPUT89), .B(n718), .Z(n883) );
  NAND2_X1 U784 ( .A1(G1996), .A2(n883), .ZN(n727) );
  NAND2_X1 U785 ( .A1(G119), .A2(n896), .ZN(n720) );
  NAND2_X1 U786 ( .A1(G107), .A2(n897), .ZN(n719) );
  NAND2_X1 U787 ( .A1(n720), .A2(n719), .ZN(n723) );
  NAND2_X1 U788 ( .A1(G131), .A2(n892), .ZN(n721) );
  XNOR2_X1 U789 ( .A(KEYINPUT87), .B(n721), .ZN(n722) );
  NOR2_X1 U790 ( .A1(n723), .A2(n722), .ZN(n725) );
  NAND2_X1 U791 ( .A1(n893), .A2(G95), .ZN(n724) );
  NAND2_X1 U792 ( .A1(n725), .A2(n724), .ZN(n888) );
  NAND2_X1 U793 ( .A1(G1991), .A2(n888), .ZN(n726) );
  NAND2_X1 U794 ( .A1(n727), .A2(n726), .ZN(n989) );
  NOR2_X1 U795 ( .A1(n729), .A2(n728), .ZN(n756) );
  NAND2_X1 U796 ( .A1(n989), .A2(n756), .ZN(n730) );
  XOR2_X1 U797 ( .A(KEYINPUT90), .B(n730), .Z(n749) );
  XNOR2_X1 U798 ( .A(G2067), .B(KEYINPUT37), .ZN(n754) );
  NAND2_X1 U799 ( .A1(n892), .A2(G140), .ZN(n731) );
  XNOR2_X1 U800 ( .A(n731), .B(KEYINPUT86), .ZN(n733) );
  NAND2_X1 U801 ( .A1(G104), .A2(n893), .ZN(n732) );
  NAND2_X1 U802 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U803 ( .A(KEYINPUT34), .B(n734), .ZN(n739) );
  NAND2_X1 U804 ( .A1(G128), .A2(n896), .ZN(n736) );
  NAND2_X1 U805 ( .A1(G116), .A2(n897), .ZN(n735) );
  NAND2_X1 U806 ( .A1(n736), .A2(n735), .ZN(n737) );
  XOR2_X1 U807 ( .A(KEYINPUT35), .B(n737), .Z(n738) );
  NOR2_X1 U808 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U809 ( .A(KEYINPUT36), .B(n740), .ZN(n905) );
  NOR2_X1 U810 ( .A1(n754), .A2(n905), .ZN(n981) );
  NAND2_X1 U811 ( .A1(n756), .A2(n981), .ZN(n752) );
  NOR2_X1 U812 ( .A1(n749), .A2(n741), .ZN(n742) );
  NAND2_X1 U813 ( .A1(n743), .A2(n742), .ZN(n744) );
  XNOR2_X1 U814 ( .A(n744), .B(KEYINPUT103), .ZN(n746) );
  XNOR2_X1 U815 ( .A(G1986), .B(G290), .ZN(n945) );
  NAND2_X1 U816 ( .A1(n945), .A2(n756), .ZN(n745) );
  NAND2_X1 U817 ( .A1(n746), .A2(n745), .ZN(n759) );
  NOR2_X1 U818 ( .A1(G1996), .A2(n883), .ZN(n975) );
  NOR2_X1 U819 ( .A1(G1986), .A2(G290), .ZN(n747) );
  NOR2_X1 U820 ( .A1(G1991), .A2(n888), .ZN(n992) );
  NOR2_X1 U821 ( .A1(n747), .A2(n992), .ZN(n748) );
  NOR2_X1 U822 ( .A1(n749), .A2(n748), .ZN(n750) );
  NOR2_X1 U823 ( .A1(n975), .A2(n750), .ZN(n751) );
  XNOR2_X1 U824 ( .A(KEYINPUT39), .B(n751), .ZN(n753) );
  NAND2_X1 U825 ( .A1(n753), .A2(n752), .ZN(n755) );
  NAND2_X1 U826 ( .A1(n754), .A2(n905), .ZN(n979) );
  NAND2_X1 U827 ( .A1(n755), .A2(n979), .ZN(n757) );
  NAND2_X1 U828 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U829 ( .A1(n759), .A2(n758), .ZN(n761) );
  XNOR2_X1 U830 ( .A(KEYINPUT40), .B(KEYINPUT104), .ZN(n760) );
  XNOR2_X1 U831 ( .A(n761), .B(n760), .ZN(G329) );
  XOR2_X1 U832 ( .A(G2438), .B(G2427), .Z(n763) );
  XNOR2_X1 U833 ( .A(G2446), .B(G2454), .ZN(n762) );
  XNOR2_X1 U834 ( .A(n763), .B(n762), .ZN(n769) );
  XOR2_X1 U835 ( .A(G2451), .B(G2430), .Z(n765) );
  XNOR2_X1 U836 ( .A(G1341), .B(G1348), .ZN(n764) );
  XNOR2_X1 U837 ( .A(n765), .B(n764), .ZN(n767) );
  XOR2_X1 U838 ( .A(G2435), .B(G2443), .Z(n766) );
  XNOR2_X1 U839 ( .A(n767), .B(n766), .ZN(n768) );
  XOR2_X1 U840 ( .A(n769), .B(n768), .Z(n770) );
  AND2_X1 U841 ( .A1(G14), .A2(n770), .ZN(G401) );
  INV_X1 U842 ( .A(G57), .ZN(G237) );
  INV_X1 U843 ( .A(G132), .ZN(G219) );
  INV_X1 U844 ( .A(G82), .ZN(G220) );
  NAND2_X1 U845 ( .A1(G94), .A2(G452), .ZN(n771) );
  XNOR2_X1 U846 ( .A(n771), .B(KEYINPUT71), .ZN(G173) );
  NAND2_X1 U847 ( .A1(G7), .A2(G661), .ZN(n772) );
  XNOR2_X1 U848 ( .A(n772), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U849 ( .A(G223), .ZN(n837) );
  NAND2_X1 U850 ( .A1(n837), .A2(G567), .ZN(n773) );
  XOR2_X1 U851 ( .A(KEYINPUT11), .B(n773), .Z(G234) );
  XOR2_X1 U852 ( .A(G860), .B(KEYINPUT73), .Z(n780) );
  NAND2_X1 U853 ( .A1(n780), .A2(n928), .ZN(n774) );
  XNOR2_X1 U854 ( .A(n774), .B(KEYINPUT74), .ZN(G153) );
  NAND2_X1 U855 ( .A1(G868), .A2(G301), .ZN(n776) );
  INV_X1 U856 ( .A(n912), .ZN(n939) );
  INV_X1 U857 ( .A(G868), .ZN(n820) );
  NAND2_X1 U858 ( .A1(n939), .A2(n820), .ZN(n775) );
  NAND2_X1 U859 ( .A1(n776), .A2(n775), .ZN(G284) );
  XOR2_X1 U860 ( .A(n936), .B(KEYINPUT72), .Z(G299) );
  NOR2_X1 U861 ( .A1(G299), .A2(G868), .ZN(n778) );
  NOR2_X1 U862 ( .A1(G286), .A2(n820), .ZN(n777) );
  NOR2_X1 U863 ( .A1(n778), .A2(n777), .ZN(G297) );
  INV_X1 U864 ( .A(G559), .ZN(n779) );
  NOR2_X1 U865 ( .A1(n780), .A2(n779), .ZN(n781) );
  NOR2_X1 U866 ( .A1(n939), .A2(n781), .ZN(n782) );
  XOR2_X1 U867 ( .A(n782), .B(KEYINPUT76), .Z(n783) );
  XNOR2_X1 U868 ( .A(KEYINPUT16), .B(n783), .ZN(G148) );
  NOR2_X1 U869 ( .A1(G559), .A2(n820), .ZN(n784) );
  NAND2_X1 U870 ( .A1(n912), .A2(n784), .ZN(n785) );
  XNOR2_X1 U871 ( .A(n785), .B(KEYINPUT77), .ZN(n787) );
  INV_X1 U872 ( .A(n928), .ZN(n810) );
  NOR2_X1 U873 ( .A1(n810), .A2(G868), .ZN(n786) );
  NOR2_X1 U874 ( .A1(n787), .A2(n786), .ZN(G282) );
  NAND2_X1 U875 ( .A1(G123), .A2(n896), .ZN(n788) );
  XNOR2_X1 U876 ( .A(n788), .B(KEYINPUT78), .ZN(n789) );
  XNOR2_X1 U877 ( .A(n789), .B(KEYINPUT18), .ZN(n791) );
  NAND2_X1 U878 ( .A1(G111), .A2(n897), .ZN(n790) );
  NAND2_X1 U879 ( .A1(n791), .A2(n790), .ZN(n795) );
  NAND2_X1 U880 ( .A1(G135), .A2(n892), .ZN(n793) );
  NAND2_X1 U881 ( .A1(G99), .A2(n893), .ZN(n792) );
  NAND2_X1 U882 ( .A1(n793), .A2(n792), .ZN(n794) );
  NOR2_X1 U883 ( .A1(n795), .A2(n794), .ZN(n983) );
  XNOR2_X1 U884 ( .A(n983), .B(G2096), .ZN(n797) );
  INV_X1 U885 ( .A(G2100), .ZN(n796) );
  NAND2_X1 U886 ( .A1(n797), .A2(n796), .ZN(G156) );
  NAND2_X1 U887 ( .A1(G67), .A2(n798), .ZN(n799) );
  XNOR2_X1 U888 ( .A(n799), .B(KEYINPUT80), .ZN(n809) );
  NAND2_X1 U889 ( .A1(G55), .A2(n800), .ZN(n803) );
  NAND2_X1 U890 ( .A1(G80), .A2(n801), .ZN(n802) );
  NAND2_X1 U891 ( .A1(n803), .A2(n802), .ZN(n807) );
  NAND2_X1 U892 ( .A1(G93), .A2(n804), .ZN(n805) );
  XNOR2_X1 U893 ( .A(KEYINPUT79), .B(n805), .ZN(n806) );
  NOR2_X1 U894 ( .A1(n807), .A2(n806), .ZN(n808) );
  NAND2_X1 U895 ( .A1(n809), .A2(n808), .ZN(n821) );
  NAND2_X1 U896 ( .A1(G559), .A2(n912), .ZN(n811) );
  XNOR2_X1 U897 ( .A(n811), .B(n810), .ZN(n818) );
  NOR2_X1 U898 ( .A1(G860), .A2(n818), .ZN(n812) );
  XOR2_X1 U899 ( .A(n821), .B(n812), .Z(G145) );
  XNOR2_X1 U900 ( .A(G299), .B(G303), .ZN(n813) );
  XNOR2_X1 U901 ( .A(n813), .B(n821), .ZN(n814) );
  XNOR2_X1 U902 ( .A(n814), .B(G290), .ZN(n815) );
  XNOR2_X1 U903 ( .A(n815), .B(G305), .ZN(n816) );
  XNOR2_X1 U904 ( .A(KEYINPUT19), .B(n816), .ZN(n817) );
  XNOR2_X1 U905 ( .A(n817), .B(G288), .ZN(n915) );
  XOR2_X1 U906 ( .A(n818), .B(n915), .Z(n819) );
  NOR2_X1 U907 ( .A1(n820), .A2(n819), .ZN(n823) );
  NOR2_X1 U908 ( .A1(G868), .A2(n821), .ZN(n822) );
  NOR2_X1 U909 ( .A1(n823), .A2(n822), .ZN(G295) );
  NAND2_X1 U910 ( .A1(G2084), .A2(G2078), .ZN(n824) );
  XOR2_X1 U911 ( .A(KEYINPUT20), .B(n824), .Z(n825) );
  NAND2_X1 U912 ( .A1(G2090), .A2(n825), .ZN(n826) );
  XNOR2_X1 U913 ( .A(KEYINPUT21), .B(n826), .ZN(n827) );
  NAND2_X1 U914 ( .A1(n827), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U915 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U916 ( .A1(G220), .A2(G219), .ZN(n828) );
  XOR2_X1 U917 ( .A(KEYINPUT22), .B(n828), .Z(n829) );
  NOR2_X1 U918 ( .A1(G218), .A2(n829), .ZN(n830) );
  XNOR2_X1 U919 ( .A(KEYINPUT84), .B(n830), .ZN(n831) );
  NAND2_X1 U920 ( .A1(n831), .A2(G96), .ZN(n842) );
  NAND2_X1 U921 ( .A1(n842), .A2(G2106), .ZN(n835) );
  NAND2_X1 U922 ( .A1(G69), .A2(G120), .ZN(n832) );
  NOR2_X1 U923 ( .A1(G237), .A2(n832), .ZN(n833) );
  NAND2_X1 U924 ( .A1(G108), .A2(n833), .ZN(n843) );
  NAND2_X1 U925 ( .A1(n843), .A2(G567), .ZN(n834) );
  NAND2_X1 U926 ( .A1(n835), .A2(n834), .ZN(n925) );
  NAND2_X1 U927 ( .A1(G661), .A2(G483), .ZN(n836) );
  NOR2_X1 U928 ( .A1(n925), .A2(n836), .ZN(n841) );
  NAND2_X1 U929 ( .A1(n841), .A2(G36), .ZN(G176) );
  NAND2_X1 U930 ( .A1(G2106), .A2(n837), .ZN(G217) );
  AND2_X1 U931 ( .A1(G15), .A2(G2), .ZN(n838) );
  NAND2_X1 U932 ( .A1(G661), .A2(n838), .ZN(G259) );
  NAND2_X1 U933 ( .A1(G3), .A2(G1), .ZN(n839) );
  XOR2_X1 U934 ( .A(KEYINPUT105), .B(n839), .Z(n840) );
  NAND2_X1 U935 ( .A1(n841), .A2(n840), .ZN(G188) );
  INV_X1 U937 ( .A(G120), .ZN(G236) );
  INV_X1 U938 ( .A(G96), .ZN(G221) );
  INV_X1 U939 ( .A(G69), .ZN(G235) );
  NOR2_X1 U940 ( .A1(n843), .A2(n842), .ZN(G325) );
  INV_X1 U941 ( .A(G325), .ZN(G261) );
  XOR2_X1 U942 ( .A(G2100), .B(KEYINPUT106), .Z(n845) );
  XNOR2_X1 U943 ( .A(KEYINPUT107), .B(KEYINPUT43), .ZN(n844) );
  XNOR2_X1 U944 ( .A(n845), .B(n844), .ZN(n849) );
  XOR2_X1 U945 ( .A(KEYINPUT42), .B(G2090), .Z(n847) );
  XNOR2_X1 U946 ( .A(G2067), .B(G2072), .ZN(n846) );
  XNOR2_X1 U947 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U948 ( .A(n849), .B(n848), .Z(n851) );
  XNOR2_X1 U949 ( .A(G2678), .B(G2096), .ZN(n850) );
  XNOR2_X1 U950 ( .A(n851), .B(n850), .ZN(n853) );
  XOR2_X1 U951 ( .A(G2084), .B(G2078), .Z(n852) );
  XNOR2_X1 U952 ( .A(n853), .B(n852), .ZN(G227) );
  XOR2_X1 U953 ( .A(G1981), .B(G1956), .Z(n855) );
  XNOR2_X1 U954 ( .A(G1986), .B(G1966), .ZN(n854) );
  XNOR2_X1 U955 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U956 ( .A(n856), .B(G2474), .Z(n858) );
  XNOR2_X1 U957 ( .A(G1971), .B(G1976), .ZN(n857) );
  XNOR2_X1 U958 ( .A(n858), .B(n857), .ZN(n862) );
  XOR2_X1 U959 ( .A(KEYINPUT41), .B(G1961), .Z(n860) );
  XNOR2_X1 U960 ( .A(G1996), .B(G1991), .ZN(n859) );
  XNOR2_X1 U961 ( .A(n860), .B(n859), .ZN(n861) );
  XNOR2_X1 U962 ( .A(n862), .B(n861), .ZN(G229) );
  NAND2_X1 U963 ( .A1(n896), .A2(G124), .ZN(n863) );
  XNOR2_X1 U964 ( .A(n863), .B(KEYINPUT44), .ZN(n865) );
  NAND2_X1 U965 ( .A1(G136), .A2(n892), .ZN(n864) );
  NAND2_X1 U966 ( .A1(n865), .A2(n864), .ZN(n866) );
  XNOR2_X1 U967 ( .A(KEYINPUT108), .B(n866), .ZN(n873) );
  NAND2_X1 U968 ( .A1(n897), .A2(G112), .ZN(n867) );
  XNOR2_X1 U969 ( .A(KEYINPUT109), .B(n867), .ZN(n870) );
  NAND2_X1 U970 ( .A1(n893), .A2(G100), .ZN(n868) );
  XOR2_X1 U971 ( .A(KEYINPUT110), .B(n868), .Z(n869) );
  NOR2_X1 U972 ( .A1(n870), .A2(n869), .ZN(n871) );
  XNOR2_X1 U973 ( .A(n871), .B(KEYINPUT111), .ZN(n872) );
  NOR2_X1 U974 ( .A1(n873), .A2(n872), .ZN(n874) );
  XNOR2_X1 U975 ( .A(KEYINPUT112), .B(n874), .ZN(G162) );
  NAND2_X1 U976 ( .A1(G130), .A2(n896), .ZN(n876) );
  NAND2_X1 U977 ( .A1(G118), .A2(n897), .ZN(n875) );
  NAND2_X1 U978 ( .A1(n876), .A2(n875), .ZN(n877) );
  XOR2_X1 U979 ( .A(KEYINPUT113), .B(n877), .Z(n882) );
  NAND2_X1 U980 ( .A1(G142), .A2(n892), .ZN(n879) );
  NAND2_X1 U981 ( .A1(G106), .A2(n893), .ZN(n878) );
  NAND2_X1 U982 ( .A1(n879), .A2(n878), .ZN(n880) );
  XOR2_X1 U983 ( .A(n880), .B(KEYINPUT45), .Z(n881) );
  NOR2_X1 U984 ( .A1(n882), .A2(n881), .ZN(n884) );
  XNOR2_X1 U985 ( .A(n884), .B(n883), .ZN(n909) );
  XOR2_X1 U986 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n886) );
  XNOR2_X1 U987 ( .A(G164), .B(KEYINPUT114), .ZN(n885) );
  XNOR2_X1 U988 ( .A(n886), .B(n885), .ZN(n887) );
  XNOR2_X1 U989 ( .A(KEYINPUT116), .B(n887), .ZN(n890) );
  XNOR2_X1 U990 ( .A(n888), .B(KEYINPUT115), .ZN(n889) );
  XNOR2_X1 U991 ( .A(n890), .B(n889), .ZN(n891) );
  XOR2_X1 U992 ( .A(n891), .B(n983), .Z(n904) );
  NAND2_X1 U993 ( .A1(G139), .A2(n892), .ZN(n895) );
  NAND2_X1 U994 ( .A1(G103), .A2(n893), .ZN(n894) );
  NAND2_X1 U995 ( .A1(n895), .A2(n894), .ZN(n902) );
  NAND2_X1 U996 ( .A1(G127), .A2(n896), .ZN(n899) );
  NAND2_X1 U997 ( .A1(G115), .A2(n897), .ZN(n898) );
  NAND2_X1 U998 ( .A1(n899), .A2(n898), .ZN(n900) );
  XOR2_X1 U999 ( .A(KEYINPUT47), .B(n900), .Z(n901) );
  NOR2_X1 U1000 ( .A1(n902), .A2(n901), .ZN(n984) );
  XNOR2_X1 U1001 ( .A(G160), .B(n984), .ZN(n903) );
  XNOR2_X1 U1002 ( .A(n904), .B(n903), .ZN(n906) );
  XNOR2_X1 U1003 ( .A(n906), .B(n905), .ZN(n907) );
  XNOR2_X1 U1004 ( .A(n907), .B(G162), .ZN(n908) );
  XOR2_X1 U1005 ( .A(n909), .B(n908), .Z(n910) );
  NOR2_X1 U1006 ( .A1(G37), .A2(n910), .ZN(n911) );
  XOR2_X1 U1007 ( .A(KEYINPUT117), .B(n911), .Z(G395) );
  XOR2_X1 U1008 ( .A(n928), .B(G286), .Z(n914) );
  XNOR2_X1 U1009 ( .A(G171), .B(n912), .ZN(n913) );
  XNOR2_X1 U1010 ( .A(n914), .B(n913), .ZN(n916) );
  XNOR2_X1 U1011 ( .A(n916), .B(n915), .ZN(n917) );
  NOR2_X1 U1012 ( .A1(G37), .A2(n917), .ZN(G397) );
  NOR2_X1 U1013 ( .A1(G227), .A2(G229), .ZN(n918) );
  XOR2_X1 U1014 ( .A(KEYINPUT49), .B(n918), .Z(n921) );
  NOR2_X1 U1015 ( .A1(G401), .A2(n925), .ZN(n919) );
  XNOR2_X1 U1016 ( .A(KEYINPUT118), .B(n919), .ZN(n920) );
  NAND2_X1 U1017 ( .A1(n921), .A2(n920), .ZN(n922) );
  XNOR2_X1 U1018 ( .A(KEYINPUT119), .B(n922), .ZN(n924) );
  NOR2_X1 U1019 ( .A1(G395), .A2(G397), .ZN(n923) );
  NAND2_X1 U1020 ( .A1(n924), .A2(n923), .ZN(G225) );
  INV_X1 U1021 ( .A(G225), .ZN(G308) );
  INV_X1 U1022 ( .A(n925), .ZN(G319) );
  INV_X1 U1023 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1024 ( .A(G16), .B(KEYINPUT56), .ZN(n949) );
  XNOR2_X1 U1025 ( .A(G171), .B(G1961), .ZN(n927) );
  NAND2_X1 U1026 ( .A1(n927), .A2(n926), .ZN(n935) );
  XNOR2_X1 U1027 ( .A(n928), .B(G1341), .ZN(n933) );
  XNOR2_X1 U1028 ( .A(G1966), .B(G168), .ZN(n930) );
  NAND2_X1 U1029 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1030 ( .A(n931), .B(KEYINPUT57), .ZN(n932) );
  NAND2_X1 U1031 ( .A1(n933), .A2(n932), .ZN(n934) );
  NOR2_X1 U1032 ( .A1(n935), .A2(n934), .ZN(n947) );
  XNOR2_X1 U1033 ( .A(n936), .B(G1956), .ZN(n938) );
  NAND2_X1 U1034 ( .A1(n938), .A2(n937), .ZN(n941) );
  XNOR2_X1 U1035 ( .A(G1348), .B(n939), .ZN(n940) );
  NOR2_X1 U1036 ( .A1(n941), .A2(n940), .ZN(n943) );
  NAND2_X1 U1037 ( .A1(G1971), .A2(G303), .ZN(n942) );
  NAND2_X1 U1038 ( .A1(n943), .A2(n942), .ZN(n944) );
  NOR2_X1 U1039 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1040 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1041 ( .A1(n949), .A2(n948), .ZN(n1031) );
  XNOR2_X1 U1042 ( .A(KEYINPUT54), .B(KEYINPUT124), .ZN(n950) );
  XNOR2_X1 U1043 ( .A(n950), .B(G34), .ZN(n951) );
  XNOR2_X1 U1044 ( .A(G2084), .B(n951), .ZN(n968) );
  XNOR2_X1 U1045 ( .A(G2090), .B(G35), .ZN(n965) );
  XOR2_X1 U1046 ( .A(G1991), .B(G25), .Z(n952) );
  NAND2_X1 U1047 ( .A1(n952), .A2(G28), .ZN(n962) );
  XNOR2_X1 U1048 ( .A(G2067), .B(G26), .ZN(n954) );
  XNOR2_X1 U1049 ( .A(G33), .B(G2072), .ZN(n953) );
  NOR2_X1 U1050 ( .A1(n954), .A2(n953), .ZN(n960) );
  XOR2_X1 U1051 ( .A(n955), .B(G32), .Z(n958) );
  XOR2_X1 U1052 ( .A(n956), .B(G27), .Z(n957) );
  NOR2_X1 U1053 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1054 ( .A1(n960), .A2(n959), .ZN(n961) );
  NOR2_X1 U1055 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1056 ( .A(KEYINPUT53), .B(n963), .ZN(n964) );
  NOR2_X1 U1057 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1058 ( .A(KEYINPUT123), .B(n966), .ZN(n967) );
  NOR2_X1 U1059 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1060 ( .A(KEYINPUT55), .B(n969), .ZN(n971) );
  INV_X1 U1061 ( .A(G29), .ZN(n970) );
  NAND2_X1 U1062 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1063 ( .A1(n972), .A2(G11), .ZN(n973) );
  XNOR2_X1 U1064 ( .A(n973), .B(KEYINPUT125), .ZN(n1003) );
  XNOR2_X1 U1065 ( .A(KEYINPUT52), .B(KEYINPUT121), .ZN(n998) );
  XOR2_X1 U1066 ( .A(G2090), .B(G162), .Z(n974) );
  NOR2_X1 U1067 ( .A1(n975), .A2(n974), .ZN(n976) );
  XOR2_X1 U1068 ( .A(n976), .B(KEYINPUT51), .Z(n977) );
  XNOR2_X1 U1069 ( .A(KEYINPUT120), .B(n977), .ZN(n978) );
  NAND2_X1 U1070 ( .A1(n979), .A2(n978), .ZN(n980) );
  NOR2_X1 U1071 ( .A1(n981), .A2(n980), .ZN(n995) );
  XOR2_X1 U1072 ( .A(G2084), .B(G160), .Z(n982) );
  NOR2_X1 U1073 ( .A1(n983), .A2(n982), .ZN(n991) );
  XOR2_X1 U1074 ( .A(G2072), .B(n984), .Z(n986) );
  XOR2_X1 U1075 ( .A(G164), .B(G2078), .Z(n985) );
  NOR2_X1 U1076 ( .A1(n986), .A2(n985), .ZN(n987) );
  XOR2_X1 U1077 ( .A(KEYINPUT50), .B(n987), .Z(n988) );
  NOR2_X1 U1078 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1079 ( .A1(n991), .A2(n990), .ZN(n993) );
  NOR2_X1 U1080 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1081 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1082 ( .A(KEYINPUT122), .B(n996), .ZN(n997) );
  XNOR2_X1 U1083 ( .A(n998), .B(n997), .ZN(n1000) );
  INV_X1 U1084 ( .A(KEYINPUT55), .ZN(n999) );
  NAND2_X1 U1085 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1086 ( .A1(G29), .A2(n1001), .ZN(n1002) );
  NAND2_X1 U1087 ( .A1(n1003), .A2(n1002), .ZN(n1029) );
  XOR2_X1 U1088 ( .A(KEYINPUT61), .B(KEYINPUT127), .Z(n1026) );
  XNOR2_X1 U1089 ( .A(G20), .B(n1004), .ZN(n1008) );
  XNOR2_X1 U1090 ( .A(G1341), .B(G19), .ZN(n1006) );
  XNOR2_X1 U1091 ( .A(G1981), .B(G6), .ZN(n1005) );
  NOR2_X1 U1092 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1093 ( .A1(n1008), .A2(n1007), .ZN(n1011) );
  XOR2_X1 U1094 ( .A(G4), .B(G1348), .Z(n1009) );
  XNOR2_X1 U1095 ( .A(KEYINPUT59), .B(n1009), .ZN(n1010) );
  NOR2_X1 U1096 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XOR2_X1 U1097 ( .A(KEYINPUT60), .B(n1012), .Z(n1014) );
  XNOR2_X1 U1098 ( .A(G1961), .B(G5), .ZN(n1013) );
  NOR2_X1 U1099 ( .A1(n1014), .A2(n1013), .ZN(n1024) );
  XNOR2_X1 U1100 ( .A(G1966), .B(KEYINPUT126), .ZN(n1015) );
  XNOR2_X1 U1101 ( .A(n1015), .B(G21), .ZN(n1022) );
  XNOR2_X1 U1102 ( .A(G1971), .B(G22), .ZN(n1017) );
  XNOR2_X1 U1103 ( .A(G23), .B(G1976), .ZN(n1016) );
  NOR2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1019) );
  XOR2_X1 U1105 ( .A(G1986), .B(G24), .Z(n1018) );
  NAND2_X1 U1106 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1107 ( .A(KEYINPUT58), .B(n1020), .ZN(n1021) );
  NOR2_X1 U1108 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1109 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1110 ( .A(n1026), .B(n1025), .ZN(n1027) );
  NOR2_X1 U1111 ( .A1(G16), .A2(n1027), .ZN(n1028) );
  NOR2_X1 U1112 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NAND2_X1 U1113 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XOR2_X1 U1114 ( .A(KEYINPUT62), .B(n1032), .Z(G311) );
  INV_X1 U1115 ( .A(G311), .ZN(G150) );
  INV_X1 U1116 ( .A(G303), .ZN(G166) );
endmodule

