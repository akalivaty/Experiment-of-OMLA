//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 0 0 1 0 0 1 0 1 1 1 1 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 0 1 0 0 1 0 1 0 0 0 0 0 1 1 1 1 1 1 0 1 1 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:44 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1304, new_n1305, new_n1306, new_n1307, new_n1308,
    new_n1309, new_n1310, new_n1311, new_n1312, new_n1313, new_n1314,
    new_n1315, new_n1316, new_n1317, new_n1318, new_n1319, new_n1320,
    new_n1321, new_n1322, new_n1323, new_n1324, new_n1325, new_n1326,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1394, new_n1395,
    new_n1396, new_n1397;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  INV_X1    g0014(.A(new_n201), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G50), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n218), .A2(new_n209), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT65), .Z(new_n222));
  XNOR2_X1  g0022(.A(KEYINPUT64), .B(G238), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n223), .A2(G68), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G116), .A2(G270), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G107), .B2(G264), .ZN(new_n227));
  NAND4_X1  g0027(.A1(new_n224), .A2(new_n225), .A3(new_n226), .A4(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n211), .B1(new_n222), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n214), .B(new_n220), .C1(KEYINPUT1), .C2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XOR2_X1   g0031(.A(G238), .B(G244), .Z(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G226), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n236), .B(new_n239), .Z(G358));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G58), .B(G77), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n241), .B(new_n242), .Z(new_n243));
  XOR2_X1   g0043(.A(G107), .B(G116), .Z(new_n244));
  XNOR2_X1  g0044(.A(G87), .B(G97), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  XNOR2_X1  g0047(.A(KEYINPUT67), .B(G1698), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(G222), .ZN(new_n249));
  XNOR2_X1  g0049(.A(KEYINPUT3), .B(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(G223), .A2(G1698), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n249), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n218), .B1(G33), .B2(G41), .ZN(new_n253));
  OAI211_X1 g0053(.A(new_n252), .B(new_n253), .C1(G77), .C2(new_n250), .ZN(new_n254));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  INV_X1    g0055(.A(G41), .ZN(new_n256));
  OAI211_X1 g0056(.A(G1), .B(G13), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G45), .ZN(new_n258));
  AOI21_X1  g0058(.A(G1), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  AND3_X1   g0059(.A1(new_n257), .A2(G274), .A3(new_n259), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n253), .A2(new_n259), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n260), .B1(G226), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n254), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G190), .ZN(new_n265));
  NAND3_X1  g0065(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(new_n218), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  XNOR2_X1  g0068(.A(KEYINPUT8), .B(G58), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n209), .A2(G33), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  NOR2_X1   g0072(.A1(G20), .A2(G33), .ZN(new_n273));
  AOI22_X1  g0073(.A1(new_n270), .A2(new_n272), .B1(G150), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n203), .A2(G20), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n268), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n278), .A2(new_n267), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n208), .A2(G20), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n279), .A2(G50), .A3(new_n280), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n281), .B1(G50), .B2(new_n277), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n276), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(KEYINPUT9), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT9), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n285), .B1(new_n276), .B2(new_n282), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n263), .A2(G200), .ZN(new_n287));
  NAND4_X1  g0087(.A1(new_n265), .A2(new_n284), .A3(new_n286), .A4(new_n287), .ZN(new_n288));
  XNOR2_X1  g0088(.A(new_n288), .B(KEYINPUT10), .ZN(new_n289));
  AND2_X1   g0089(.A1(KEYINPUT68), .A2(G179), .ZN(new_n290));
  NOR2_X1   g0090(.A1(KEYINPUT68), .A2(G179), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n264), .A2(new_n292), .ZN(new_n293));
  OAI221_X1 g0093(.A(new_n293), .B1(G169), .B2(new_n264), .C1(new_n276), .C2(new_n282), .ZN(new_n294));
  INV_X1    g0094(.A(new_n273), .ZN(new_n295));
  INV_X1    g0095(.A(G77), .ZN(new_n296));
  OAI22_X1  g0096(.A1(new_n269), .A2(new_n295), .B1(new_n209), .B2(new_n296), .ZN(new_n297));
  XNOR2_X1  g0097(.A(KEYINPUT15), .B(G87), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n298), .A2(new_n271), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n267), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n279), .A2(G77), .A3(new_n280), .ZN(new_n301));
  NOR3_X1   g0101(.A1(new_n277), .A2(KEYINPUT69), .A3(G77), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT69), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n303), .B1(new_n278), .B2(new_n296), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n300), .B(new_n301), .C1(new_n302), .C2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G232), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT3), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(new_n255), .ZN(new_n308));
  NAND2_X1  g0108(.A1(KEYINPUT3), .A2(G33), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n306), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  AND2_X1   g0110(.A1(KEYINPUT3), .A2(G33), .ZN(new_n311));
  NOR2_X1   g0111(.A1(KEYINPUT3), .A2(G33), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AOI22_X1  g0113(.A1(new_n310), .A2(new_n248), .B1(new_n313), .B2(G107), .ZN(new_n314));
  INV_X1    g0114(.A(G1698), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n315), .B1(new_n308), .B2(new_n309), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(new_n223), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n314), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(new_n253), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n260), .B1(G244), .B2(new_n261), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n305), .B1(new_n322), .B2(G190), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n321), .A2(G200), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(G169), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n321), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n319), .A2(new_n292), .A3(new_n320), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n328), .A2(new_n305), .A3(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n326), .A2(new_n331), .ZN(new_n332));
  AND3_X1   g0132(.A1(new_n289), .A2(new_n294), .A3(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n260), .B1(G232), .B2(new_n261), .ZN(new_n334));
  OAI211_X1 g0134(.A(G226), .B(G1698), .C1(new_n311), .C2(new_n312), .ZN(new_n335));
  INV_X1    g0135(.A(G87), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n335), .B1(new_n255), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n315), .A2(KEYINPUT67), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT67), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(G1698), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n338), .B(new_n340), .C1(new_n311), .C2(new_n312), .ZN(new_n341));
  INV_X1    g0141(.A(G223), .ZN(new_n342));
  OAI21_X1  g0142(.A(KEYINPUT78), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT78), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n250), .A2(new_n248), .A3(new_n344), .A4(G223), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n337), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n334), .B1(new_n346), .B2(new_n257), .ZN(new_n347));
  INV_X1    g0147(.A(G200), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(G190), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n350), .B(new_n334), .C1(new_n346), .C2(new_n257), .ZN(new_n351));
  AND2_X1   g0151(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT17), .ZN(new_n353));
  INV_X1    g0153(.A(G58), .ZN(new_n354));
  INV_X1    g0154(.A(G68), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  OAI21_X1  g0156(.A(G20), .B1(new_n356), .B2(new_n201), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n273), .A2(G159), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT7), .ZN(new_n361));
  NOR4_X1   g0161(.A1(new_n311), .A2(new_n312), .A3(new_n361), .A4(G20), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT76), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n363), .B1(new_n311), .B2(new_n312), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n308), .A2(KEYINPUT76), .A3(new_n309), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n364), .A2(new_n365), .A3(new_n209), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n362), .B1(new_n366), .B2(new_n361), .ZN(new_n367));
  OAI211_X1 g0167(.A(KEYINPUT16), .B(new_n360), .C1(new_n367), .C2(new_n355), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT16), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n361), .B1(new_n250), .B2(G20), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n313), .A2(KEYINPUT7), .A3(new_n209), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n355), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n369), .B1(new_n372), .B2(new_n359), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n368), .A2(new_n267), .A3(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n279), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n270), .A2(new_n280), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n375), .B1(new_n376), .B2(KEYINPUT77), .ZN(new_n377));
  OR2_X1    g0177(.A1(new_n376), .A2(KEYINPUT77), .ZN(new_n378));
  AOI22_X1  g0178(.A1(new_n377), .A2(new_n378), .B1(new_n278), .B2(new_n269), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n374), .A2(new_n379), .ZN(new_n380));
  NOR3_X1   g0180(.A1(new_n352), .A2(new_n353), .A3(new_n380), .ZN(new_n381));
  AND2_X1   g0181(.A1(new_n374), .A2(new_n379), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n349), .A2(new_n351), .ZN(new_n383));
  AOI21_X1  g0183(.A(KEYINPUT17), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n347), .A2(G169), .ZN(new_n386));
  INV_X1    g0186(.A(new_n292), .ZN(new_n387));
  OAI211_X1 g0187(.A(new_n387), .B(new_n334), .C1(new_n346), .C2(new_n257), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT18), .ZN(new_n390));
  AND3_X1   g0190(.A1(new_n380), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n390), .B1(new_n380), .B2(new_n389), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(KEYINPUT79), .B1(new_n385), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n380), .A2(new_n389), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(KEYINPUT18), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n353), .B1(new_n352), .B2(new_n380), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n380), .A2(new_n389), .A3(new_n390), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n382), .A2(KEYINPUT17), .A3(new_n383), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n396), .A2(new_n397), .A3(new_n398), .A4(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT79), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n333), .B1(new_n394), .B2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT75), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n278), .A2(new_n355), .ZN(new_n405));
  XNOR2_X1  g0205(.A(new_n405), .B(KEYINPUT12), .ZN(new_n406));
  AOI22_X1  g0206(.A1(new_n273), .A2(G50), .B1(G20), .B2(new_n355), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n407), .B1(new_n296), .B2(new_n271), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n408), .A2(KEYINPUT11), .A3(new_n267), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n279), .A2(G68), .A3(new_n280), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n406), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(KEYINPUT11), .B1(new_n408), .B2(new_n267), .ZN(new_n412));
  OR2_X1    g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT72), .ZN(new_n414));
  INV_X1    g0214(.A(new_n260), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n261), .A2(G238), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(G33), .A2(G97), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT71), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(KEYINPUT71), .A2(G33), .A3(G97), .ZN(new_n421));
  AOI22_X1  g0221(.A1(new_n310), .A2(G1698), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(G226), .ZN(new_n423));
  OAI21_X1  g0223(.A(KEYINPUT70), .B1(new_n341), .B2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT70), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n250), .A2(new_n248), .A3(new_n425), .A4(G226), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n422), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n417), .B1(new_n427), .B2(new_n253), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT13), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n414), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  AND2_X1   g0230(.A1(new_n427), .A2(new_n253), .ZN(new_n431));
  OAI21_X1  g0231(.A(KEYINPUT13), .B1(new_n431), .B2(new_n417), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n414), .B(KEYINPUT13), .C1(new_n431), .C2(new_n417), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n433), .A2(G169), .A3(new_n434), .ZN(new_n435));
  AND2_X1   g0235(.A1(new_n435), .A2(KEYINPUT14), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT14), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n433), .A2(new_n437), .A3(G169), .A4(new_n434), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n428), .A2(new_n429), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n432), .A2(G179), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(KEYINPUT74), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT74), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n432), .A2(new_n442), .A3(new_n439), .A4(G179), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n438), .A2(new_n441), .A3(new_n443), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n413), .B1(new_n436), .B2(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n433), .A2(G200), .A3(new_n434), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n350), .B1(new_n428), .B2(new_n429), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n413), .B1(new_n447), .B2(new_n432), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT73), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n446), .A2(KEYINPUT73), .A3(new_n448), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n404), .B1(new_n445), .B2(new_n453), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n403), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n445), .A2(new_n404), .A3(new_n453), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(G107), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n278), .A2(KEYINPUT25), .A3(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(KEYINPUT25), .B1(new_n278), .B2(new_n458), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n208), .A2(G33), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n277), .A2(new_n462), .A3(new_n218), .A4(new_n266), .ZN(new_n463));
  OAI22_X1  g0263(.A1(new_n460), .A2(new_n461), .B1(new_n458), .B2(new_n463), .ZN(new_n464));
  AND3_X1   g0264(.A1(new_n458), .A2(KEYINPUT23), .A3(G20), .ZN(new_n465));
  AOI21_X1  g0265(.A(KEYINPUT23), .B1(new_n458), .B2(G20), .ZN(new_n466));
  NAND2_X1  g0266(.A1(G33), .A2(G116), .ZN(new_n467));
  OAI22_X1  g0267(.A1(new_n465), .A2(new_n466), .B1(G20), .B2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT83), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(KEYINPUT22), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n250), .A2(new_n209), .A3(G87), .A4(new_n470), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n209), .B(G87), .C1(new_n311), .C2(new_n312), .ZN(new_n472));
  INV_X1    g0272(.A(new_n470), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AOI211_X1 g0274(.A(KEYINPUT24), .B(new_n468), .C1(new_n471), .C2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT24), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n474), .A2(new_n471), .ZN(new_n477));
  INV_X1    g0277(.A(new_n468), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n267), .B1(new_n475), .B2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT84), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  OAI211_X1 g0282(.A(KEYINPUT84), .B(new_n267), .C1(new_n475), .C2(new_n479), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n464), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n338), .A2(new_n340), .A3(G250), .ZN(new_n485));
  NAND2_X1  g0285(.A1(G257), .A2(G1698), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n313), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(G294), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n255), .A2(new_n488), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n253), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  OR2_X1    g0290(.A1(KEYINPUT5), .A2(G41), .ZN(new_n491));
  NAND2_X1  g0291(.A1(KEYINPUT5), .A2(G41), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n258), .A2(G1), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n493), .A2(new_n257), .A3(G274), .A4(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n253), .B1(new_n494), .B2(new_n493), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(G264), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n490), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n348), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(KEYINPUT85), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT85), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n498), .A2(new_n501), .A3(new_n348), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n500), .B(new_n502), .C1(G190), .C2(new_n498), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n484), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n498), .A2(new_n327), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n505), .B1(G179), .B2(new_n498), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n504), .B1(new_n484), .B2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT21), .ZN(new_n508));
  OAI211_X1 g0308(.A(G264), .B(G1698), .C1(new_n311), .C2(new_n312), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n308), .A2(G303), .A3(new_n309), .ZN(new_n510));
  AND2_X1   g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n250), .A2(new_n248), .A3(G257), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n257), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(new_n492), .ZN(new_n514));
  NOR2_X1   g0314(.A1(KEYINPUT5), .A2(G41), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n494), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n257), .ZN(new_n517));
  INV_X1    g0317(.A(G270), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n495), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g0319(.A(G169), .B1(new_n513), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n277), .A2(G116), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(G116), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n522), .B1(new_n463), .B2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT20), .ZN(new_n525));
  OR2_X1    g0325(.A1(KEYINPUT80), .A2(G97), .ZN(new_n526));
  NAND2_X1  g0326(.A1(KEYINPUT80), .A2(G97), .ZN(new_n527));
  AOI21_X1  g0327(.A(G33), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(G33), .A2(G283), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n209), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n266), .A2(new_n218), .B1(G20), .B2(new_n523), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n525), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  OAI211_X1 g0334(.A(KEYINPUT20), .B(new_n532), .C1(new_n528), .C2(new_n530), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n524), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n508), .B1(new_n520), .B2(new_n536), .ZN(new_n537));
  AND2_X1   g0337(.A1(new_n257), .A2(G274), .ZN(new_n538));
  INV_X1    g0338(.A(new_n516), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n496), .A2(G270), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(G257), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n341), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n509), .A2(new_n510), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n253), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n540), .A2(new_n544), .A3(G190), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n513), .A2(new_n519), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n536), .B(new_n545), .C1(new_n546), .C2(new_n348), .ZN(new_n547));
  INV_X1    g0347(.A(G179), .ZN(new_n548));
  NOR3_X1   g0348(.A1(new_n513), .A2(new_n548), .A3(new_n519), .ZN(new_n549));
  INV_X1    g0349(.A(new_n524), .ZN(new_n550));
  AND2_X1   g0350(.A1(KEYINPUT80), .A2(G97), .ZN(new_n551));
  NOR2_X1   g0351(.A1(KEYINPUT80), .A2(G97), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n209), .B(new_n529), .C1(new_n553), .C2(G33), .ZN(new_n554));
  AOI21_X1  g0354(.A(KEYINPUT20), .B1(new_n554), .B2(new_n532), .ZN(new_n555));
  INV_X1    g0355(.A(new_n535), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n550), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n549), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n540), .A2(new_n544), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n557), .A2(new_n559), .A3(KEYINPUT21), .A4(G169), .ZN(new_n560));
  AND4_X1   g0360(.A1(new_n537), .A2(new_n547), .A3(new_n558), .A4(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n298), .A2(new_n278), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n463), .A2(new_n336), .ZN(new_n564));
  AND3_X1   g0364(.A1(KEYINPUT71), .A2(G33), .A3(G97), .ZN(new_n565));
  AOI21_X1  g0365(.A(KEYINPUT71), .B1(G33), .B2(G97), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT19), .ZN(new_n567));
  NOR3_X1   g0367(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  OAI21_X1  g0368(.A(KEYINPUT82), .B1(new_n568), .B2(G20), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n420), .A2(KEYINPUT19), .A3(new_n421), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT82), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n570), .A2(new_n571), .A3(new_n209), .ZN(new_n572));
  NOR2_X1   g0372(.A1(G87), .A2(G107), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n553), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n569), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n250), .A2(new_n209), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n271), .B1(new_n526), .B2(new_n527), .ZN(new_n577));
  OAI22_X1  g0377(.A1(new_n576), .A2(new_n355), .B1(new_n577), .B2(KEYINPUT19), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n575), .A2(new_n579), .ZN(new_n580));
  AOI211_X1 g0380(.A(new_n563), .B(new_n564), .C1(new_n580), .C2(new_n267), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n257), .A2(G274), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n208), .A2(G45), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(G250), .ZN(new_n584));
  OAI22_X1  g0384(.A1(new_n582), .A2(new_n583), .B1(new_n253), .B2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(G244), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n586), .A2(new_n315), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n587), .B1(new_n248), .B2(G238), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n467), .B1(new_n588), .B2(new_n313), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n585), .B1(new_n589), .B2(new_n253), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n350), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n591), .B1(G200), .B2(new_n590), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n338), .A2(new_n340), .A3(G238), .ZN(new_n593));
  INV_X1    g0393(.A(new_n587), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n313), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(new_n467), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n253), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n253), .A2(new_n584), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n598), .B1(new_n538), .B2(new_n494), .ZN(new_n599));
  AOI21_X1  g0399(.A(G169), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n600), .B1(new_n292), .B2(new_n590), .ZN(new_n601));
  INV_X1    g0401(.A(new_n463), .ZN(new_n602));
  INV_X1    g0402(.A(new_n298), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n570), .A2(new_n209), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n605), .A2(KEYINPUT82), .B1(new_n553), .B2(new_n573), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n578), .B1(new_n606), .B2(new_n572), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n562), .B(new_n604), .C1(new_n607), .C2(new_n268), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n581), .A2(new_n592), .B1(new_n601), .B2(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n495), .B1(new_n517), .B2(new_n541), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT4), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n611), .B1(new_n341), .B2(new_n586), .ZN(new_n612));
  INV_X1    g0412(.A(new_n529), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n613), .B1(new_n316), .B2(G250), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n250), .A2(new_n248), .A3(KEYINPUT4), .A4(G244), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n612), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n610), .B1(new_n616), .B2(new_n253), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(G190), .ZN(new_n618));
  AOI21_X1  g0418(.A(KEYINPUT7), .B1(new_n313), .B2(new_n209), .ZN(new_n619));
  OAI21_X1  g0419(.A(G107), .B1(new_n619), .B2(new_n362), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n295), .A2(new_n296), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT6), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n622), .A2(G107), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n623), .B1(new_n551), .B2(new_n552), .ZN(new_n624));
  AND2_X1   g0424(.A1(G97), .A2(G107), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n622), .B1(new_n625), .B2(new_n205), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n621), .B1(new_n627), .B2(G20), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n268), .B1(new_n620), .B2(new_n628), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n277), .A2(G97), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n630), .B1(new_n602), .B2(G97), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n617), .A2(KEYINPUT81), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(G200), .B1(new_n617), .B2(KEYINPUT81), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n618), .B(new_n633), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n616), .A2(new_n253), .ZN(new_n638));
  INV_X1    g0438(.A(new_n610), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n327), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n620), .A2(new_n628), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n631), .B1(new_n642), .B2(new_n268), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n617), .A2(new_n292), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n641), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n561), .A2(new_n609), .A3(new_n637), .A4(new_n645), .ZN(new_n646));
  NOR3_X1   g0446(.A1(new_n457), .A2(new_n507), .A3(new_n646), .ZN(G372));
  INV_X1    g0447(.A(new_n294), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n435), .A2(KEYINPUT14), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n649), .A2(new_n438), .A3(new_n441), .A4(new_n443), .ZN(new_n650));
  AOI22_X1  g0450(.A1(new_n453), .A2(new_n331), .B1(new_n650), .B2(new_n413), .ZN(new_n651));
  INV_X1    g0451(.A(new_n385), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n393), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n648), .B1(new_n653), .B2(new_n289), .ZN(new_n654));
  OAI22_X1  g0454(.A1(new_n617), .A2(G169), .B1(new_n629), .B2(new_n632), .ZN(new_n655));
  AOI211_X1 g0455(.A(new_n387), .B(new_n610), .C1(new_n616), .C2(new_n253), .ZN(new_n656));
  OAI21_X1  g0456(.A(KEYINPUT89), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT89), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n641), .A2(new_n658), .A3(new_n643), .A4(new_n644), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT86), .ZN(new_n661));
  AOI21_X1  g0461(.A(G200), .B1(new_n597), .B2(new_n599), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n662), .B1(new_n350), .B2(new_n590), .ZN(new_n663));
  INV_X1    g0463(.A(new_n564), .ZN(new_n664));
  OAI211_X1 g0464(.A(new_n562), .B(new_n664), .C1(new_n607), .C2(new_n268), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n597), .A2(new_n599), .A3(new_n292), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n667), .B1(new_n590), .B2(G169), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n563), .B1(new_n580), .B2(new_n267), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n668), .B1(new_n669), .B2(new_n604), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n661), .B1(new_n666), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n601), .A2(new_n608), .ZN(new_n672));
  OAI211_X1 g0472(.A(new_n672), .B(KEYINPUT86), .C1(new_n665), .C2(new_n663), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT26), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n660), .A2(new_n671), .A3(new_n673), .A4(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT88), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n670), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n672), .A2(KEYINPUT88), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n655), .A2(new_n656), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n609), .A2(new_n680), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n679), .B1(KEYINPUT26), .B2(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n537), .A2(new_n558), .A3(new_n560), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n482), .A2(new_n483), .ZN(new_n684));
  INV_X1    g0484(.A(new_n464), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT87), .ZN(new_n687));
  INV_X1    g0487(.A(new_n506), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n686), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(KEYINPUT87), .B1(new_n484), .B2(new_n506), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n683), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n636), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(new_n634), .ZN(new_n693));
  AND2_X1   g0493(.A1(new_n618), .A2(new_n633), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n680), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n695), .A2(new_n671), .A3(new_n504), .A4(new_n673), .ZN(new_n696));
  OAI211_X1 g0496(.A(new_n675), .B(new_n682), .C1(new_n691), .C2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n654), .B1(new_n457), .B2(new_n698), .ZN(G369));
  OR2_X1    g0499(.A1(new_n561), .A2(KEYINPUT91), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n561), .A2(KEYINPUT91), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n702), .A2(KEYINPUT27), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(KEYINPUT27), .ZN(new_n704));
  AND3_X1   g0504(.A1(new_n703), .A2(G213), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(G343), .ZN(new_n706));
  XNOR2_X1  g0506(.A(new_n706), .B(KEYINPUT90), .ZN(new_n707));
  OAI211_X1 g0507(.A(new_n700), .B(new_n701), .C1(new_n536), .C2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n683), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n707), .A2(new_n536), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(G330), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n484), .A2(new_n707), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n506), .B1(new_n684), .B2(new_n685), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  OAI22_X1  g0517(.A1(new_n507), .A2(new_n715), .B1(new_n717), .B2(new_n707), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n714), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n689), .A2(new_n690), .A3(new_n707), .ZN(new_n720));
  INV_X1    g0520(.A(new_n707), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n709), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n717), .A2(new_n722), .A3(new_n504), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n719), .A2(new_n720), .A3(new_n723), .ZN(G399));
  INV_X1    g0524(.A(new_n212), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(G41), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n574), .A2(G116), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n727), .A2(G1), .A3(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n729), .B1(new_n216), .B2(new_n727), .ZN(new_n730));
  XNOR2_X1  g0530(.A(new_n730), .B(KEYINPUT28), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n697), .A2(new_n707), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT29), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n660), .A2(new_n671), .A3(new_n673), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(KEYINPUT26), .ZN(new_n736));
  NOR3_X1   g0536(.A1(new_n666), .A2(new_n670), .A3(new_n645), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n679), .B1(new_n737), .B2(new_n674), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT94), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n739), .B1(new_n716), .B2(new_n683), .ZN(new_n740));
  OAI211_X1 g0540(.A(new_n709), .B(KEYINPUT94), .C1(new_n484), .C2(new_n506), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  OAI211_X1 g0542(.A(new_n736), .B(new_n738), .C1(new_n742), .C2(new_n696), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n743), .A2(KEYINPUT29), .A3(new_n707), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n734), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g0545(.A(KEYINPUT92), .B(KEYINPUT31), .ZN(new_n746));
  AND4_X1   g0546(.A1(new_n497), .A2(new_n490), .A3(new_n597), .A4(new_n599), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n747), .A2(KEYINPUT30), .A3(new_n549), .A4(new_n617), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n387), .B1(new_n597), .B2(new_n599), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n640), .A2(new_n498), .A3(new_n559), .A4(new_n749), .ZN(new_n750));
  AND2_X1   g0550(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n747), .A2(new_n549), .A3(new_n617), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT30), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  AOI211_X1 g0554(.A(new_n707), .B(new_n746), .C1(new_n751), .C2(new_n754), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n490), .A2(new_n597), .A3(new_n497), .A4(new_n599), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n540), .A2(new_n544), .A3(G179), .ZN(new_n757));
  NOR3_X1   g0557(.A1(new_n640), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(KEYINPUT93), .B1(new_n758), .B2(KEYINPUT30), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT93), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n752), .A2(new_n760), .A3(new_n753), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n751), .A2(new_n759), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(new_n721), .ZN(new_n763));
  INV_X1    g0563(.A(KEYINPUT31), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n755), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n646), .ZN(new_n766));
  NAND4_X1  g0566(.A1(new_n766), .A2(new_n504), .A3(new_n717), .A4(new_n707), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n713), .B1(new_n765), .B2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n745), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(KEYINPUT95), .ZN(new_n771));
  INV_X1    g0571(.A(KEYINPUT95), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n745), .A2(new_n772), .A3(new_n769), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n731), .B1(new_n774), .B2(G1), .ZN(G364));
  XNOR2_X1  g0575(.A(new_n714), .B(KEYINPUT96), .ZN(new_n776));
  INV_X1    g0576(.A(G13), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(G20), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n208), .B1(new_n778), .B2(G45), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n726), .A2(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n781), .B1(new_n712), .B2(new_n713), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n776), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n212), .A2(new_n250), .ZN(new_n784));
  INV_X1    g0584(.A(G355), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n784), .A2(new_n785), .B1(G116), .B2(new_n212), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n364), .A2(new_n365), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n725), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n789), .B1(new_n258), .B2(new_n217), .ZN(new_n790));
  OR2_X1    g0590(.A1(new_n243), .A2(new_n258), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n786), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(G13), .A2(G33), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(G20), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n218), .B1(G20), .B2(new_n327), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n781), .B1(new_n792), .B2(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n209), .A2(G179), .ZN(new_n800));
  NOR2_X1   g0600(.A1(G190), .A2(G200), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(G159), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  XNOR2_X1  g0604(.A(KEYINPUT97), .B(KEYINPUT32), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n292), .A2(new_n209), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n350), .A2(G200), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n807), .A2(new_n801), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n806), .B1(new_n354), .B2(new_n809), .C1(new_n296), .C2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n808), .A2(new_n548), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(G20), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(G97), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n800), .A2(new_n350), .A3(G200), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n818), .A2(new_n458), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n800), .A2(G190), .A3(G200), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n820), .A2(new_n336), .ZN(new_n821));
  NOR4_X1   g0621(.A1(new_n817), .A2(new_n819), .A3(new_n821), .A4(new_n313), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n807), .A2(G190), .A3(G200), .ZN(new_n823));
  OAI211_X1 g0623(.A(new_n812), .B(new_n822), .C1(new_n202), .C2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n807), .A2(G200), .ZN(new_n825));
  OR3_X1    g0625(.A1(new_n825), .A2(KEYINPUT98), .A3(G190), .ZN(new_n826));
  OAI21_X1  g0626(.A(KEYINPUT98), .B1(new_n825), .B2(G190), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n829), .A2(new_n355), .ZN(new_n830));
  INV_X1    g0630(.A(G283), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n818), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n802), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n250), .B1(new_n833), .B2(G329), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n834), .B1(new_n488), .B2(new_n815), .ZN(new_n835));
  INV_X1    g0635(.A(new_n820), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n832), .B(new_n835), .C1(G303), .C2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n810), .ZN(new_n838));
  INV_X1    g0638(.A(new_n809), .ZN(new_n839));
  AOI22_X1  g0639(.A1(G311), .A2(new_n838), .B1(new_n839), .B2(G322), .ZN(new_n840));
  INV_X1    g0640(.A(G326), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n837), .B(new_n840), .C1(new_n841), .C2(new_n823), .ZN(new_n842));
  XOR2_X1   g0642(.A(KEYINPUT33), .B(G317), .Z(new_n843));
  NOR2_X1   g0643(.A1(new_n829), .A2(new_n843), .ZN(new_n844));
  OAI22_X1  g0644(.A1(new_n824), .A2(new_n830), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  OR2_X1    g0645(.A1(new_n845), .A2(KEYINPUT99), .ZN(new_n846));
  INV_X1    g0646(.A(new_n796), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n847), .B1(new_n845), .B2(KEYINPUT99), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n799), .B1(new_n846), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n712), .ZN(new_n850));
  INV_X1    g0650(.A(new_n795), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n849), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  AND3_X1   g0652(.A1(new_n783), .A2(KEYINPUT100), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(KEYINPUT100), .B1(new_n783), .B2(new_n852), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(G396));
  NAND2_X1  g0656(.A1(new_n330), .A2(KEYINPUT102), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n721), .A2(new_n305), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT102), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n328), .A2(new_n859), .A3(new_n305), .A4(new_n329), .ZN(new_n860));
  NAND4_X1  g0660(.A1(new_n857), .A2(new_n325), .A3(new_n858), .A4(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n331), .A2(new_n721), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n732), .A2(new_n864), .ZN(new_n865));
  AND2_X1   g0665(.A1(new_n857), .A2(new_n860), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n867), .A2(new_n326), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n697), .A2(new_n707), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n865), .A2(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n781), .B1(new_n870), .B2(new_n769), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n865), .A2(new_n768), .A3(new_n869), .ZN(new_n872));
  AND2_X1   g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n863), .A2(new_n794), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n796), .A2(new_n793), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n781), .B1(G77), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n828), .A2(G283), .ZN(new_n878));
  INV_X1    g0678(.A(new_n823), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(G303), .ZN(new_n880));
  INV_X1    g0680(.A(G311), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n313), .B1(new_n802), .B2(new_n881), .ZN(new_n882));
  OAI22_X1  g0682(.A1(new_n336), .A2(new_n818), .B1(new_n820), .B2(new_n458), .ZN(new_n883));
  NOR3_X1   g0683(.A1(new_n817), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  AOI22_X1  g0684(.A1(G116), .A2(new_n838), .B1(new_n839), .B2(G294), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n878), .A2(new_n880), .A3(new_n884), .A4(new_n885), .ZN(new_n886));
  AOI22_X1  g0686(.A1(G143), .A2(new_n839), .B1(new_n838), .B2(G159), .ZN(new_n887));
  INV_X1    g0687(.A(G137), .ZN(new_n888));
  INV_X1    g0688(.A(G150), .ZN(new_n889));
  OAI221_X1 g0689(.A(new_n887), .B1(new_n888), .B2(new_n823), .C1(new_n829), .C2(new_n889), .ZN(new_n890));
  XNOR2_X1  g0690(.A(new_n890), .B(KEYINPUT101), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT34), .ZN(new_n892));
  AND2_X1   g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n787), .ZN(new_n894));
  INV_X1    g0694(.A(new_n818), .ZN(new_n895));
  AOI22_X1  g0695(.A1(G68), .A2(new_n895), .B1(new_n814), .B2(G58), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n896), .B1(new_n202), .B2(new_n820), .ZN(new_n897));
  AOI211_X1 g0697(.A(new_n894), .B(new_n897), .C1(G132), .C2(new_n833), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n898), .B1(new_n891), .B2(new_n892), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n886), .B1(new_n893), .B2(new_n899), .ZN(new_n900));
  AOI211_X1 g0700(.A(new_n874), .B(new_n877), .C1(new_n900), .C2(new_n796), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n873), .A2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(G384));
  NOR2_X1   g0703(.A1(new_n778), .A2(new_n208), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT38), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n382), .A2(new_n383), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT37), .ZN(new_n907));
  INV_X1    g0707(.A(new_n705), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n386), .A2(new_n388), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n380), .ZN(new_n910));
  AND3_X1   g0710(.A1(new_n906), .A2(new_n907), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n366), .A2(new_n361), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n371), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(G68), .ZN(new_n914));
  AOI21_X1  g0714(.A(KEYINPUT16), .B1(new_n914), .B2(new_n360), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n368), .A2(new_n267), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n379), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(KEYINPUT103), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT103), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n919), .B(new_n379), .C1(new_n915), .C2(new_n916), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n918), .A2(new_n920), .A3(new_n909), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(new_n906), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n911), .B1(new_n922), .B2(KEYINPUT37), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n918), .A2(new_n705), .A3(new_n920), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n924), .B1(new_n385), .B2(new_n393), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n905), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n924), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n400), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n907), .B1(new_n921), .B2(new_n906), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n928), .B(KEYINPUT38), .C1(new_n929), .C2(new_n911), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n926), .A2(new_n930), .ZN(new_n931));
  AND3_X1   g0731(.A1(new_n446), .A2(KEYINPUT73), .A3(new_n448), .ZN(new_n932));
  AOI21_X1  g0732(.A(KEYINPUT73), .B1(new_n446), .B2(new_n448), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n413), .B(new_n721), .C1(new_n934), .C2(new_n650), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n721), .A2(new_n413), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n445), .A2(new_n453), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n746), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n939), .B1(new_n762), .B2(new_n721), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n760), .B1(new_n752), .B2(new_n753), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n748), .A2(new_n750), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n707), .B1(new_n943), .B2(new_n761), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n940), .B1(KEYINPUT31), .B2(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n864), .B1(new_n945), .B2(new_n767), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n931), .A2(new_n938), .A3(new_n946), .ZN(new_n947));
  XOR2_X1   g0747(.A(KEYINPUT106), .B(KEYINPUT40), .Z(new_n948));
  NAND3_X1  g0748(.A1(new_n762), .A2(KEYINPUT31), .A3(new_n721), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(new_n944), .B2(new_n939), .ZN(new_n950));
  NOR3_X1   g0750(.A1(new_n507), .A2(new_n646), .A3(new_n721), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n863), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n952), .B1(new_n937), .B2(new_n935), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT40), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n380), .A2(new_n705), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n955), .B1(new_n385), .B2(new_n393), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n906), .A2(new_n910), .ZN(new_n957));
  AOI21_X1  g0757(.A(KEYINPUT104), .B1(new_n909), .B2(new_n380), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n957), .B1(new_n907), .B2(new_n958), .ZN(new_n959));
  NAND4_X1  g0759(.A1(new_n906), .A2(KEYINPUT104), .A3(new_n910), .A4(KEYINPUT37), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n905), .B1(new_n956), .B2(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n954), .B1(new_n962), .B2(new_n930), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n947), .A2(new_n948), .B1(new_n953), .B2(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n950), .A2(new_n951), .ZN(new_n966));
  OR2_X1    g0766(.A1(new_n457), .A2(new_n966), .ZN(new_n967));
  AND2_X1   g0767(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n965), .A2(new_n967), .ZN(new_n969));
  NOR3_X1   g0769(.A1(new_n968), .A2(new_n969), .A3(new_n713), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n931), .A2(KEYINPUT39), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT105), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT39), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n962), .A2(new_n974), .A3(new_n930), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n972), .A2(new_n973), .A3(new_n975), .ZN(new_n976));
  AND3_X1   g0776(.A1(new_n962), .A2(new_n974), .A3(new_n930), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n974), .B1(new_n926), .B2(new_n930), .ZN(new_n978));
  OAI21_X1  g0778(.A(KEYINPUT105), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n650), .A2(new_n413), .A3(new_n707), .ZN(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n976), .A2(new_n979), .A3(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n393), .A2(new_n705), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n867), .A2(new_n707), .ZN(new_n984));
  AOI22_X1  g0784(.A1(new_n869), .A2(new_n984), .B1(new_n937), .B2(new_n935), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n983), .B1(new_n985), .B2(new_n931), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n982), .A2(new_n986), .ZN(new_n987));
  NAND4_X1  g0787(.A1(new_n734), .A2(new_n455), .A3(new_n456), .A4(new_n744), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(new_n654), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n987), .B(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n904), .B1(new_n971), .B2(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n991), .B1(new_n990), .B2(new_n971), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n219), .A2(G116), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n993), .B1(new_n627), .B2(KEYINPUT35), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(KEYINPUT35), .B2(new_n627), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT36), .ZN(new_n996));
  NOR3_X1   g0796(.A1(new_n216), .A2(new_n296), .A3(new_n356), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n355), .A2(G50), .ZN(new_n998));
  OAI211_X1 g0798(.A(G1), .B(new_n777), .C1(new_n997), .C2(new_n998), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n992), .A2(new_n996), .A3(new_n999), .ZN(G367));
  OAI221_X1 g0800(.A(new_n797), .B1(new_n212), .B2(new_n298), .C1(new_n789), .C2(new_n239), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(new_n781), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n836), .A2(G116), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT46), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(new_n823), .B2(new_n881), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(G283), .A2(new_n838), .B1(new_n839), .B2(G303), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n787), .B1(G317), .B2(new_n833), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n526), .A2(new_n527), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n1008), .A2(new_n895), .B1(new_n814), .B2(G107), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1006), .A2(new_n1007), .A3(new_n1009), .ZN(new_n1010));
  AOI211_X1 g0810(.A(new_n1005), .B(new_n1010), .C1(G294), .C2(new_n828), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT108), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n818), .A2(new_n296), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n1013), .A2(new_n313), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT109), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1015), .B1(G143), .B2(new_n879), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n814), .A2(G68), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n1017), .B1(new_n354), .B2(new_n820), .C1(new_n888), .C2(new_n802), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n202), .A2(new_n810), .B1(new_n809), .B2(new_n889), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n1016), .B(new_n1020), .C1(new_n803), .C2(new_n829), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1012), .A2(new_n1021), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT47), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1002), .B1(new_n1023), .B2(new_n796), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n671), .A2(new_n673), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n581), .A2(new_n707), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(new_n679), .B2(new_n1026), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1028), .A2(new_n795), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1024), .A2(new_n1029), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n637), .B(new_n645), .C1(new_n633), .C2(new_n707), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n680), .A2(new_n721), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n720), .A2(new_n723), .A3(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT107), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT45), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  OR2_X1    g0837(.A1(new_n1034), .A2(KEYINPUT107), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1034), .A2(KEYINPUT107), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1038), .A2(KEYINPUT45), .A3(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT44), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n720), .A2(new_n723), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n1042), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1041), .B1(new_n1043), .B2(new_n1033), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1033), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1042), .A2(KEYINPUT44), .A3(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1037), .A2(new_n1040), .A3(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n719), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n1035), .A2(new_n1036), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1051), .A2(new_n719), .A3(new_n1040), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1053));
  OR2_X1    g0853(.A1(new_n718), .A2(new_n722), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1054), .A2(new_n723), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n776), .A2(new_n1055), .ZN(new_n1056));
  NOR3_X1   g0856(.A1(new_n1055), .A2(new_n713), .A3(new_n712), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n774), .B1(new_n1053), .B2(new_n1059), .ZN(new_n1060));
  XOR2_X1   g0860(.A(new_n726), .B(KEYINPUT41), .Z(new_n1061));
  INV_X1    g0861(.A(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n780), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1063));
  OR2_X1    g0863(.A1(new_n1045), .A2(new_n723), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(KEYINPUT42), .ZN(new_n1065));
  AND2_X1   g0865(.A1(new_n716), .A2(new_n637), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n707), .B1(new_n1066), .B2(new_n680), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1065), .A2(new_n1067), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n1064), .A2(KEYINPUT42), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT43), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n1068), .A2(new_n1069), .B1(new_n1070), .B2(new_n1028), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1028), .A2(new_n1070), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1071), .B(new_n1072), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n719), .A2(new_n1045), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1073), .B(new_n1074), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1030), .B1(new_n1063), .B2(new_n1075), .ZN(G387));
  NAND3_X1  g0876(.A1(new_n1059), .A2(new_n773), .A3(new_n771), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1057), .B1(new_n776), .B2(new_n1055), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n774), .A2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1077), .A2(new_n1079), .A3(new_n726), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n781), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n789), .B1(new_n236), .B2(G45), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n728), .B(new_n258), .C1(new_n355), .C2(new_n296), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT110), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1086));
  OAI21_X1  g0886(.A(KEYINPUT50), .B1(new_n269), .B2(G50), .ZN(new_n1087));
  OR3_X1    g0887(.A1(new_n269), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1082), .B1(new_n1085), .B2(new_n1089), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n1090), .B1(G107), .B2(new_n212), .C1(new_n728), .C2(new_n784), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1081), .B1(new_n1091), .B2(new_n797), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1092), .B1(new_n718), .B2(new_n851), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n787), .B1(new_n816), .B2(new_n818), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n202), .A2(new_n809), .B1(new_n810), .B2(new_n355), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n1094), .B(new_n1095), .C1(new_n603), .C2(new_n814), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n836), .A2(G77), .B1(new_n833), .B2(G150), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n1097), .A2(KEYINPUT111), .B1(new_n823), .B2(new_n803), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(KEYINPUT111), .B2(new_n1097), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n1096), .B(new_n1099), .C1(new_n269), .C2(new_n829), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n815), .A2(new_n831), .B1(new_n820), .B2(new_n488), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n879), .A2(G322), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1102), .B1(new_n829), .B2(new_n881), .ZN(new_n1103));
  OR2_X1    g0903(.A1(new_n1103), .A2(KEYINPUT112), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1103), .A2(KEYINPUT112), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(G303), .A2(new_n838), .B1(new_n839), .B2(G317), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1104), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT48), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1101), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1109), .B1(new_n1108), .B2(new_n1107), .ZN(new_n1110));
  XOR2_X1   g0910(.A(new_n1110), .B(KEYINPUT49), .Z(new_n1111));
  OAI221_X1 g0911(.A(new_n894), .B1(new_n523), .B2(new_n818), .C1(new_n841), .C2(new_n802), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT113), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1100), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1093), .B1(new_n1114), .B2(new_n796), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1115), .B1(new_n780), .B2(new_n1078), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1080), .A2(new_n1116), .ZN(G393));
  INV_X1    g0917(.A(new_n1079), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1053), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n727), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT114), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1121), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n719), .B1(new_n1051), .B2(new_n1040), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1123), .A2(KEYINPUT114), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1079), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1120), .A2(new_n1125), .ZN(new_n1126));
  NOR3_X1   g0926(.A1(new_n1122), .A2(new_n1124), .A3(new_n779), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT116), .ZN(new_n1128));
  OAI221_X1 g0928(.A(new_n797), .B1(new_n212), .B2(new_n553), .C1(new_n789), .C2(new_n246), .ZN(new_n1129));
  AND2_X1   g0929(.A1(new_n1129), .A2(new_n781), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n250), .B(new_n819), .C1(G322), .C2(new_n833), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1131), .B1(new_n831), .B2(new_n820), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n879), .A2(G317), .B1(new_n839), .B2(G311), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(new_n1133), .B(KEYINPUT52), .ZN(new_n1134));
  AOI211_X1 g0934(.A(new_n1132), .B(new_n1134), .C1(G294), .C2(new_n838), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n828), .A2(G303), .B1(G116), .B2(new_n814), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(new_n1136), .B(KEYINPUT115), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n823), .A2(new_n889), .B1(new_n809), .B2(new_n803), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1138), .B(KEYINPUT51), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(G87), .A2(new_n895), .B1(new_n814), .B2(G77), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1140), .B1(new_n355), .B2(new_n820), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n894), .B1(G143), .B2(new_n833), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1142), .B1(new_n269), .B2(new_n810), .ZN(new_n1143));
  AOI211_X1 g0943(.A(new_n1141), .B(new_n1143), .C1(new_n828), .C2(G50), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n1135), .A2(new_n1137), .B1(new_n1139), .B2(new_n1144), .ZN(new_n1145));
  OAI221_X1 g0945(.A(new_n1130), .B1(new_n1033), .B2(new_n851), .C1(new_n1145), .C2(new_n847), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  NOR3_X1   g0947(.A1(new_n1127), .A2(new_n1128), .A3(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1052), .ZN(new_n1149));
  OAI21_X1  g0949(.A(KEYINPUT114), .B1(new_n1149), .B2(new_n1123), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1050), .A2(new_n1121), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1150), .A2(new_n780), .A3(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(KEYINPUT116), .B1(new_n1152), .B2(new_n1146), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1126), .B1(new_n1148), .B2(new_n1153), .ZN(G390));
  NOR2_X1   g0954(.A1(new_n966), .A2(new_n713), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n455), .A2(new_n1155), .A3(new_n456), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n988), .A2(new_n654), .A3(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n869), .A2(new_n984), .ZN(new_n1158));
  AOI211_X1 g0958(.A(new_n713), .B(new_n864), .C1(new_n765), .C2(new_n767), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1159), .A2(new_n938), .ZN(new_n1160));
  OAI211_X1 g0960(.A(G330), .B(new_n863), .C1(new_n950), .C2(new_n951), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(new_n937), .B2(new_n935), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1158), .B1(new_n1160), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1159), .A2(new_n938), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n743), .A2(new_n707), .A3(new_n868), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1161), .A2(new_n937), .A3(new_n935), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n1164), .A2(new_n984), .A3(new_n1165), .A4(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1157), .B1(new_n1163), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1158), .A2(new_n938), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(new_n980), .ZN(new_n1171));
  NOR3_X1   g0971(.A1(new_n977), .A2(new_n978), .A3(KEYINPUT105), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n973), .B1(new_n972), .B2(new_n975), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1171), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1165), .A2(new_n984), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1175), .A2(new_n938), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT117), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n981), .B1(new_n962), .B2(new_n930), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n1165), .A2(new_n984), .B1(new_n937), .B2(new_n935), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1178), .ZN(new_n1181));
  OAI21_X1  g0981(.A(KEYINPUT117), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1179), .A2(new_n1182), .ZN(new_n1183));
  AND3_X1   g0983(.A1(new_n1174), .A2(new_n1183), .A3(new_n1164), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1162), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(new_n1174), .B2(new_n1183), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1169), .B1(new_n1184), .B2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1174), .A2(new_n1183), .A3(new_n1164), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n976), .A2(new_n979), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n1189), .A2(new_n1171), .B1(new_n1179), .B2(new_n1182), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n1188), .B(new_n1168), .C1(new_n1190), .C2(new_n1185), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1187), .A2(new_n726), .A3(new_n1191), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1188), .B(new_n780), .C1(new_n1190), .C2(new_n1185), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1189), .A2(new_n793), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1081), .B1(new_n269), .B2(new_n875), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(KEYINPUT54), .B(G143), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n810), .A2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n313), .B1(new_n833), .B2(G125), .ZN(new_n1198));
  OAI221_X1 g0998(.A(new_n1198), .B1(new_n202), .B2(new_n818), .C1(new_n803), .C2(new_n815), .ZN(new_n1199));
  AOI211_X1 g0999(.A(new_n1197), .B(new_n1199), .C1(G132), .C2(new_n839), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT53), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1201), .B1(new_n820), .B2(new_n889), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n836), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n879), .A2(G128), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1200), .B(new_n1204), .C1(new_n888), .C2(new_n829), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n313), .B1(new_n802), .B2(new_n488), .C1(new_n336), .C2(new_n820), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n815), .A2(new_n296), .B1(new_n818), .B2(new_n355), .ZN(new_n1207));
  AOI211_X1 g1007(.A(new_n1206), .B(new_n1207), .C1(G116), .C2(new_n839), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n828), .A2(G107), .B1(new_n1008), .B2(new_n838), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n1208), .B1(new_n831), .B2(new_n823), .C1(new_n1209), .C2(KEYINPUT118), .ZN(new_n1210));
  AND2_X1   g1010(.A1(new_n1209), .A2(KEYINPUT118), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1205), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT119), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1215), .A2(new_n796), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n1194), .B(new_n1195), .C1(new_n1214), .C2(new_n1216), .ZN(new_n1217));
  AND2_X1   g1017(.A1(new_n1193), .A2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1192), .A2(new_n1218), .ZN(G378));
  NAND2_X1  g1019(.A1(new_n289), .A2(new_n294), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n283), .A2(new_n908), .ZN(new_n1221));
  XNOR2_X1  g1021(.A(new_n1220), .B(new_n1221), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  XNOR2_X1  g1024(.A(new_n1222), .B(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1226), .A2(new_n793), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n781), .B1(G50), .B2(new_n876), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n894), .A2(new_n256), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n809), .A2(new_n458), .ZN(new_n1230));
  AOI211_X1 g1030(.A(new_n1229), .B(new_n1230), .C1(new_n603), .C2(new_n838), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n836), .A2(G77), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n895), .A2(G58), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n833), .A2(G283), .ZN(new_n1234));
  NAND4_X1  g1034(.A1(new_n1232), .A2(new_n1233), .A3(new_n1017), .A4(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(new_n879), .B2(G116), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n1231), .B(new_n1236), .C1(new_n829), .C2(new_n816), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT58), .ZN(new_n1238));
  AOI21_X1  g1038(.A(G50), .B1(new_n255), .B2(new_n256), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(new_n1237), .A2(new_n1238), .B1(new_n1229), .B2(new_n1239), .ZN(new_n1240));
  OR2_X1    g1040(.A1(new_n820), .A2(new_n1196), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT120), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n1241), .A2(new_n1242), .B1(new_n815), .B2(new_n889), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(new_n879), .B2(G125), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n839), .A2(G128), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n838), .A2(G137), .B1(new_n1242), .B2(new_n1241), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1244), .A2(new_n1245), .A3(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1247), .B1(G132), .B2(new_n828), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(KEYINPUT59), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n895), .A2(G159), .ZN(new_n1251));
  AOI211_X1 g1051(.A(G33), .B(G41), .C1(new_n833), .C2(G124), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1250), .A2(new_n1251), .A3(new_n1252), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1249), .A2(KEYINPUT59), .ZN(new_n1254));
  OAI221_X1 g1054(.A(new_n1240), .B1(new_n1238), .B2(new_n1237), .C1(new_n1253), .C2(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1228), .B1(new_n1255), .B2(new_n796), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1227), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n947), .A2(new_n948), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n953), .A2(new_n963), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1259), .A2(G330), .A3(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(new_n1226), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n964), .A2(G330), .A3(new_n1225), .ZN(new_n1263));
  AND4_X1   g1063(.A1(KEYINPUT121), .A2(new_n987), .A3(new_n1262), .A4(new_n1263), .ZN(new_n1264));
  AOI22_X1  g1064(.A1(KEYINPUT121), .A2(new_n987), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1258), .B1(new_n1266), .B2(new_n780), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1157), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1191), .A2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT57), .ZN(new_n1270));
  AND4_X1   g1070(.A1(G330), .A2(new_n1259), .A3(new_n1260), .A4(new_n1225), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1225), .B1(new_n964), .B2(G330), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n987), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1262), .A2(new_n982), .A3(new_n1263), .A4(new_n986), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1270), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1269), .A2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(new_n726), .ZN(new_n1277));
  AOI21_X1  g1077(.A(KEYINPUT57), .B1(new_n1269), .B2(new_n1266), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1267), .B1(new_n1277), .B2(new_n1278), .ZN(G375));
  NAND2_X1  g1079(.A1(new_n1163), .A2(new_n1167), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1280), .A2(new_n780), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n781), .B1(G68), .B2(new_n876), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n894), .B1(G128), .B2(new_n833), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1283), .B1(new_n889), .B2(new_n810), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1284), .B1(G137), .B2(new_n839), .ZN(new_n1285));
  OAI221_X1 g1085(.A(new_n1233), .B1(new_n803), .B2(new_n820), .C1(new_n815), .C2(new_n202), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1286), .B1(new_n879), .B2(G132), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1285), .A2(new_n1287), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n829), .A2(new_n1196), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n829), .A2(new_n523), .ZN(new_n1290));
  AOI22_X1  g1090(.A1(G107), .A2(new_n838), .B1(new_n839), .B2(G283), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n879), .A2(G294), .ZN(new_n1292));
  AOI211_X1 g1092(.A(new_n250), .B(new_n1013), .C1(G303), .C2(new_n833), .ZN(new_n1293));
  AOI22_X1  g1093(.A1(G97), .A2(new_n836), .B1(new_n814), .B2(new_n603), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1291), .A2(new_n1292), .A3(new_n1293), .A4(new_n1294), .ZN(new_n1295));
  OAI22_X1  g1095(.A1(new_n1288), .A2(new_n1289), .B1(new_n1290), .B2(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1282), .B1(new_n1296), .B2(new_n796), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1297), .B1(new_n938), .B2(new_n794), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1281), .A2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1299), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1157), .A2(new_n1163), .A3(new_n1167), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1169), .A2(new_n1062), .A3(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1300), .A2(new_n1302), .ZN(G381));
  OAI21_X1  g1103(.A(new_n1128), .B1(new_n1127), .B2(new_n1147), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1152), .A2(KEYINPUT116), .A3(new_n1146), .ZN(new_n1305));
  AOI22_X1  g1105(.A1(new_n1304), .A2(new_n1305), .B1(new_n1120), .B2(new_n1125), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1307), .A2(new_n779), .ZN(new_n1308));
  XOR2_X1   g1108(.A(new_n1073), .B(new_n1074), .Z(new_n1309));
  AOI22_X1  g1109(.A1(new_n1308), .A2(new_n1309), .B1(new_n1029), .B2(new_n1024), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1306), .A2(new_n1310), .ZN(new_n1311));
  AND3_X1   g1111(.A1(new_n1080), .A2(new_n855), .A3(new_n1116), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1312), .ZN(new_n1313));
  NOR4_X1   g1113(.A1(new_n1311), .A2(G384), .A3(G381), .A4(new_n1313), .ZN(new_n1314));
  XNOR2_X1  g1114(.A(new_n1314), .B(KEYINPUT122), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n987), .A2(KEYINPUT121), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1317));
  XNOR2_X1  g1117(.A(new_n1316), .B(new_n1317), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1257), .B1(new_n1318), .B2(new_n779), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1269), .A2(new_n1266), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1320), .A2(new_n1270), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n727), .B1(new_n1269), .B2(new_n1275), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1319), .B1(new_n1321), .B2(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(G378), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1315), .A2(new_n1326), .ZN(G407));
  OAI211_X1 g1127(.A(G407), .B(G213), .C1(G343), .C2(new_n1325), .ZN(G409));
  AOI21_X1  g1128(.A(new_n855), .B1(new_n1080), .B2(new_n1116), .ZN(new_n1329));
  NOR2_X1   g1129(.A1(new_n1312), .A2(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1330), .A2(KEYINPUT124), .ZN(new_n1331));
  INV_X1    g1131(.A(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT124), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1333), .B1(new_n1312), .B2(new_n1329), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1334), .B1(G390), .B2(G387), .ZN(new_n1335));
  NOR2_X1   g1135(.A1(new_n1306), .A2(new_n1310), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1332), .B1(new_n1335), .B2(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT61), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(G390), .A2(G387), .ZN(new_n1339));
  NAND4_X1  g1139(.A1(new_n1339), .A2(new_n1311), .A3(new_n1331), .A4(new_n1334), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1337), .A2(new_n1338), .A3(new_n1340), .ZN(new_n1341));
  INV_X1    g1141(.A(KEYINPUT125), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1341), .A2(new_n1342), .ZN(new_n1343));
  NAND4_X1  g1143(.A1(new_n1337), .A2(KEYINPUT125), .A3(new_n1338), .A4(new_n1340), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1343), .A2(new_n1344), .ZN(new_n1345));
  INV_X1    g1145(.A(G213), .ZN(new_n1346));
  NOR2_X1   g1146(.A1(new_n1346), .A2(G343), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1348));
  AOI21_X1  g1148(.A(new_n1258), .B1(new_n1348), .B2(new_n780), .ZN(new_n1349));
  AND3_X1   g1149(.A1(new_n1192), .A2(new_n1218), .A3(new_n1349), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1269), .A2(new_n1266), .A3(new_n1062), .ZN(new_n1351));
  AOI21_X1  g1151(.A(new_n1347), .B1(new_n1350), .B2(new_n1351), .ZN(new_n1352));
  INV_X1    g1152(.A(KEYINPUT60), .ZN(new_n1353));
  OAI21_X1  g1153(.A(new_n1301), .B1(new_n1168), .B2(new_n1353), .ZN(new_n1354));
  NAND4_X1  g1154(.A1(new_n1157), .A2(new_n1163), .A3(KEYINPUT60), .A4(new_n1167), .ZN(new_n1355));
  AND2_X1   g1155(.A1(new_n1355), .A2(new_n726), .ZN(new_n1356));
  AOI211_X1 g1156(.A(new_n902), .B(new_n1299), .C1(new_n1354), .C2(new_n1356), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1354), .A2(new_n1356), .ZN(new_n1358));
  AOI21_X1  g1158(.A(G384), .B1(new_n1358), .B2(new_n1300), .ZN(new_n1359));
  NOR2_X1   g1159(.A1(new_n1357), .A2(new_n1359), .ZN(new_n1360));
  OAI211_X1 g1160(.A(new_n1352), .B(new_n1360), .C1(new_n1324), .C2(new_n1323), .ZN(new_n1361));
  INV_X1    g1161(.A(new_n1361), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1362), .A2(KEYINPUT63), .ZN(new_n1363));
  INV_X1    g1163(.A(KEYINPUT63), .ZN(new_n1364));
  OAI21_X1  g1164(.A(new_n1352), .B1(new_n1324), .B2(new_n1323), .ZN(new_n1365));
  NOR3_X1   g1165(.A1(new_n1357), .A2(new_n1359), .A3(KEYINPUT123), .ZN(new_n1366));
  OAI21_X1  g1166(.A(KEYINPUT123), .B1(new_n1357), .B2(new_n1359), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1347), .A2(G2897), .ZN(new_n1368));
  INV_X1    g1168(.A(new_n1368), .ZN(new_n1369));
  NAND2_X1  g1169(.A1(new_n1367), .A2(new_n1369), .ZN(new_n1370));
  OAI211_X1 g1170(.A(KEYINPUT123), .B(new_n1368), .C1(new_n1357), .C2(new_n1359), .ZN(new_n1371));
  AOI21_X1  g1171(.A(new_n1366), .B1(new_n1370), .B2(new_n1371), .ZN(new_n1372));
  AOI21_X1  g1172(.A(new_n1364), .B1(new_n1365), .B2(new_n1372), .ZN(new_n1373));
  OAI211_X1 g1173(.A(new_n1345), .B(new_n1363), .C1(new_n1362), .C2(new_n1373), .ZN(new_n1374));
  NOR2_X1   g1174(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1375));
  NAND2_X1  g1175(.A1(new_n1350), .A2(new_n1351), .ZN(new_n1376));
  INV_X1    g1176(.A(new_n1347), .ZN(new_n1377));
  NAND2_X1  g1177(.A1(new_n1376), .A2(new_n1377), .ZN(new_n1378));
  OAI21_X1  g1178(.A(new_n1372), .B1(new_n1375), .B2(new_n1378), .ZN(new_n1379));
  NAND2_X1  g1179(.A1(G375), .A2(G378), .ZN(new_n1380));
  INV_X1    g1180(.A(KEYINPUT62), .ZN(new_n1381));
  NAND4_X1  g1181(.A1(new_n1380), .A2(new_n1381), .A3(new_n1360), .A4(new_n1352), .ZN(new_n1382));
  AND3_X1   g1182(.A1(new_n1379), .A2(new_n1338), .A3(new_n1382), .ZN(new_n1383));
  NAND2_X1  g1183(.A1(new_n1361), .A2(KEYINPUT62), .ZN(new_n1384));
  AOI21_X1  g1184(.A(KEYINPUT126), .B1(new_n1383), .B2(new_n1384), .ZN(new_n1385));
  AOI21_X1  g1185(.A(KEYINPUT61), .B1(new_n1365), .B2(new_n1372), .ZN(new_n1386));
  NAND4_X1  g1186(.A1(new_n1386), .A2(new_n1384), .A3(KEYINPUT126), .A4(new_n1382), .ZN(new_n1387));
  INV_X1    g1187(.A(KEYINPUT127), .ZN(new_n1388));
  AND3_X1   g1188(.A1(new_n1337), .A2(new_n1388), .A3(new_n1340), .ZN(new_n1389));
  AOI21_X1  g1189(.A(new_n1388), .B1(new_n1337), .B2(new_n1340), .ZN(new_n1390));
  NOR2_X1   g1190(.A1(new_n1389), .A2(new_n1390), .ZN(new_n1391));
  NAND2_X1  g1191(.A1(new_n1387), .A2(new_n1391), .ZN(new_n1392));
  OAI21_X1  g1192(.A(new_n1374), .B1(new_n1385), .B2(new_n1392), .ZN(G405));
  OAI21_X1  g1193(.A(new_n1360), .B1(new_n1326), .B2(new_n1375), .ZN(new_n1394));
  OAI211_X1 g1194(.A(new_n1325), .B(new_n1380), .C1(new_n1359), .C2(new_n1357), .ZN(new_n1395));
  NAND2_X1  g1195(.A1(new_n1394), .A2(new_n1395), .ZN(new_n1396));
  NAND2_X1  g1196(.A1(new_n1337), .A2(new_n1340), .ZN(new_n1397));
  XOR2_X1   g1197(.A(new_n1396), .B(new_n1397), .Z(G402));
endmodule


