

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733;

  NOR2_X1 U370 ( .A1(n606), .A2(n707), .ZN(n367) );
  NOR2_X1 U371 ( .A1(n699), .A2(n707), .ZN(n701) );
  NOR2_X1 U372 ( .A1(n689), .A2(n707), .ZN(n371) );
  NAND2_X1 U373 ( .A1(n376), .A2(n416), .ZN(n722) );
  INV_X1 U374 ( .A(KEYINPUT35), .ZN(n347) );
  XNOR2_X1 U375 ( .A(n512), .B(KEYINPUT4), .ZN(n490) );
  XOR2_X1 U376 ( .A(KEYINPUT72), .B(KEYINPUT75), .Z(n487) );
  XNOR2_X1 U377 ( .A(KEYINPUT71), .B(KEYINPUT3), .ZN(n467) );
  XOR2_X1 U378 ( .A(G104), .B(G146), .Z(n352) );
  XNOR2_X2 U379 ( .A(n348), .B(n347), .ZN(n731) );
  NAND2_X1 U380 ( .A1(n359), .A2(n358), .ZN(n348) );
  XNOR2_X1 U381 ( .A(G116), .B(G119), .ZN(n469) );
  XNOR2_X1 U382 ( .A(n490), .B(n402), .ZN(n474) );
  XNOR2_X1 U383 ( .A(n361), .B(n418), .ZN(n376) );
  XOR2_X1 U384 ( .A(KEYINPUT90), .B(n474), .Z(n720) );
  XNOR2_X1 U385 ( .A(G125), .B(G146), .ZN(n362) );
  NAND2_X1 U386 ( .A1(n550), .A2(n350), .ZN(n361) );
  AND2_X1 U387 ( .A1(n414), .A2(n413), .ZN(n412) );
  OR2_X1 U388 ( .A1(n693), .A2(n410), .ZN(n409) );
  INV_X1 U389 ( .A(n362), .ZN(n489) );
  XNOR2_X1 U390 ( .A(n598), .B(KEYINPUT45), .ZN(n599) );
  INV_X2 U391 ( .A(G953), .ZN(n723) );
  BUF_X1 U392 ( .A(n644), .Z(n349) );
  XNOR2_X2 U393 ( .A(n591), .B(KEYINPUT89), .ZN(n585) );
  XNOR2_X1 U394 ( .A(n481), .B(n480), .ZN(n483) );
  XNOR2_X1 U395 ( .A(n429), .B(n428), .ZN(n550) );
  INV_X1 U396 ( .A(n632), .ZN(n380) );
  XOR2_X1 U397 ( .A(G122), .B(G104), .Z(n497) );
  XOR2_X1 U398 ( .A(G116), .B(G107), .Z(n513) );
  NAND2_X1 U399 ( .A1(n412), .A2(n409), .ZN(n406) );
  XNOR2_X1 U400 ( .A(n504), .B(n354), .ZN(n547) );
  XNOR2_X1 U401 ( .A(n489), .B(G140), .ZN(n450) );
  NAND2_X1 U402 ( .A1(n386), .A2(n385), .ZN(n360) );
  NOR2_X1 U403 ( .A1(n722), .A2(n639), .ZN(n385) );
  INV_X1 U404 ( .A(n638), .ZN(n386) );
  XNOR2_X1 U405 ( .A(n425), .B(n424), .ZN(n423) );
  INV_X1 U406 ( .A(n702), .ZN(n424) );
  NAND2_X1 U407 ( .A1(n703), .A2(G478), .ZN(n425) );
  INV_X1 U408 ( .A(KEYINPUT48), .ZN(n418) );
  XNOR2_X1 U409 ( .A(KEYINPUT9), .B(KEYINPUT104), .ZN(n506) );
  XNOR2_X1 U410 ( .A(n427), .B(n426), .ZN(n505) );
  INV_X1 U411 ( .A(KEYINPUT8), .ZN(n426) );
  NAND2_X1 U412 ( .A1(n723), .A2(G234), .ZN(n427) );
  XNOR2_X1 U413 ( .A(n366), .B(n431), .ZN(n603) );
  XNOR2_X1 U414 ( .A(n484), .B(n474), .ZN(n366) );
  XNOR2_X1 U415 ( .A(n401), .B(n400), .ZN(n708) );
  XNOR2_X1 U416 ( .A(n482), .B(n513), .ZN(n400) );
  XNOR2_X1 U417 ( .A(n483), .B(n484), .ZN(n401) );
  XNOR2_X1 U418 ( .A(n383), .B(n382), .ZN(n696) );
  XNOR2_X1 U419 ( .A(n500), .B(n503), .ZN(n382) );
  XNOR2_X1 U420 ( .A(n719), .B(n384), .ZN(n383) );
  XNOR2_X1 U421 ( .A(n708), .B(n394), .ZN(n684) );
  XNOR2_X1 U422 ( .A(n395), .B(n399), .ZN(n394) );
  XNOR2_X1 U423 ( .A(n490), .B(n488), .ZN(n399) );
  XNOR2_X1 U424 ( .A(n398), .B(n396), .ZN(n395) );
  NAND2_X1 U425 ( .A1(n407), .A2(n412), .ZN(n405) );
  NAND2_X1 U426 ( .A1(n406), .A2(n533), .ZN(n357) );
  AND2_X1 U427 ( .A1(n409), .A2(n408), .ZN(n407) );
  INV_X1 U428 ( .A(KEYINPUT0), .ZN(n562) );
  XNOR2_X1 U429 ( .A(n459), .B(n458), .ZN(n460) );
  AND2_X1 U430 ( .A1(n388), .A2(n356), .ZN(n387) );
  XNOR2_X1 U431 ( .A(n445), .B(n369), .ZN(n446) );
  XNOR2_X1 U432 ( .A(n487), .B(n352), .ZN(n369) );
  NOR2_X1 U433 ( .A1(G952), .A2(n723), .ZN(n707) );
  XNOR2_X1 U434 ( .A(n532), .B(KEYINPUT64), .ZN(n428) );
  OR2_X1 U435 ( .A1(n664), .A2(n622), .ZN(n379) );
  XOR2_X1 U436 ( .A(KEYINPUT103), .B(KEYINPUT101), .Z(n509) );
  XNOR2_X1 U437 ( .A(G122), .B(G134), .ZN(n508) );
  XOR2_X1 U438 ( .A(KEYINPUT102), .B(KEYINPUT7), .Z(n507) );
  NOR2_X1 U439 ( .A1(n626), .A2(n628), .ZN(n664) );
  OR2_X1 U440 ( .A1(G902), .A2(G237), .ZN(n492) );
  XNOR2_X1 U441 ( .A(n456), .B(n374), .ZN(n462) );
  XNOR2_X1 U442 ( .A(n457), .B(KEYINPUT94), .ZN(n374) );
  XOR2_X1 U443 ( .A(KEYINPUT95), .B(KEYINPUT20), .Z(n457) );
  NOR2_X1 U444 ( .A1(G237), .A2(G953), .ZN(n471) );
  XNOR2_X1 U445 ( .A(n365), .B(G146), .ZN(n470) );
  INV_X1 U446 ( .A(KEYINPUT5), .ZN(n365) );
  XOR2_X1 U447 ( .A(KEYINPUT99), .B(G131), .Z(n499) );
  XNOR2_X1 U448 ( .A(G143), .B(G113), .ZN(n498) );
  XNOR2_X1 U449 ( .A(n502), .B(n501), .ZN(n384) );
  XNOR2_X1 U450 ( .A(KEYINPUT15), .B(G902), .ZN(n601) );
  XNOR2_X1 U451 ( .A(n404), .B(n403), .ZN(n402) );
  XNOR2_X1 U452 ( .A(KEYINPUT70), .B(G131), .ZN(n404) );
  XNOR2_X1 U453 ( .A(G134), .B(G137), .ZN(n403) );
  XNOR2_X1 U454 ( .A(n489), .B(n487), .ZN(n398) );
  XNOR2_X1 U455 ( .A(n491), .B(n397), .ZN(n396) );
  INV_X1 U456 ( .A(KEYINPUT85), .ZN(n397) );
  NAND2_X1 U457 ( .A1(G237), .A2(G234), .ZN(n432) );
  NAND2_X1 U458 ( .A1(G469), .A2(n411), .ZN(n410) );
  INV_X1 U459 ( .A(G902), .ZN(n411) );
  NAND2_X1 U460 ( .A1(n415), .A2(G902), .ZN(n413) );
  NAND2_X1 U461 ( .A1(n650), .A2(n651), .ZN(n590) );
  NAND2_X1 U462 ( .A1(n373), .A2(n646), .ZN(n573) );
  INV_X1 U463 ( .A(n567), .ZN(n373) );
  AND2_X1 U464 ( .A1(n636), .A2(n417), .ZN(n416) );
  INV_X1 U465 ( .A(n635), .ZN(n417) );
  XOR2_X1 U466 ( .A(n518), .B(n517), .Z(n702) );
  NOR2_X1 U467 ( .A1(n638), .A2(n722), .ZN(n390) );
  INV_X1 U468 ( .A(n601), .ZN(n389) );
  XNOR2_X1 U469 ( .A(n442), .B(n441), .ZN(n443) );
  INV_X1 U470 ( .A(G140), .ZN(n441) );
  XNOR2_X1 U471 ( .A(n541), .B(n540), .ZN(n561) );
  XNOR2_X1 U472 ( .A(n547), .B(KEYINPUT100), .ZN(n529) );
  NOR2_X1 U473 ( .A1(G902), .A2(n603), .ZN(n475) );
  INV_X1 U474 ( .A(n649), .ZN(n589) );
  XNOR2_X1 U475 ( .A(n603), .B(n602), .ZN(n604) );
  XNOR2_X1 U476 ( .A(n453), .B(n452), .ZN(n454) );
  INV_X1 U477 ( .A(G137), .ZN(n452) );
  XNOR2_X1 U478 ( .A(n696), .B(n695), .ZN(n697) );
  XNOR2_X1 U479 ( .A(n686), .B(n685), .ZN(n687) );
  AND2_X1 U480 ( .A1(n381), .A2(n650), .ZN(n632) );
  INV_X1 U481 ( .A(n577), .ZN(n358) );
  XNOR2_X1 U482 ( .A(n392), .B(n391), .ZN(n732) );
  INV_X1 U483 ( .A(KEYINPUT32), .ZN(n391) );
  AND2_X1 U484 ( .A1(n572), .A2(n536), .ZN(n393) );
  OR2_X1 U485 ( .A1(n529), .A2(n524), .ZN(n623) );
  INV_X1 U486 ( .A(KEYINPUT124), .ZN(n421) );
  INV_X1 U487 ( .A(n707), .ZN(n422) );
  XNOR2_X1 U488 ( .A(n691), .B(n370), .ZN(n694) );
  AND2_X1 U489 ( .A1(n380), .A2(n351), .ZN(n350) );
  XOR2_X1 U490 ( .A(n535), .B(n649), .Z(n582) );
  AND2_X1 U491 ( .A1(n377), .A2(n621), .ZN(n351) );
  NAND2_X2 U492 ( .A1(n357), .A2(n405), .ZN(n650) );
  INV_X1 U493 ( .A(G469), .ZN(n415) );
  AND2_X1 U494 ( .A1(G210), .A2(n492), .ZN(n353) );
  XOR2_X1 U495 ( .A(KEYINPUT13), .B(G475), .Z(n354) );
  XOR2_X1 U496 ( .A(KEYINPUT80), .B(KEYINPUT34), .Z(n355) );
  XOR2_X1 U497 ( .A(n600), .B(KEYINPUT69), .Z(n356) );
  XNOR2_X1 U498 ( .A(n576), .B(n355), .ZN(n359) );
  NOR2_X1 U499 ( .A1(n705), .A2(G902), .ZN(n461) );
  XOR2_X2 U500 ( .A(n545), .B(KEYINPUT38), .Z(n660) );
  XNOR2_X2 U501 ( .A(n360), .B(KEYINPUT77), .ZN(n644) );
  INV_X1 U502 ( .A(n534), .ZN(n420) );
  XNOR2_X2 U503 ( .A(n531), .B(KEYINPUT40), .ZN(n733) );
  NAND2_X1 U504 ( .A1(n420), .A2(n372), .ZN(n465) );
  INV_X1 U505 ( .A(n573), .ZN(n372) );
  NOR2_X1 U506 ( .A1(n521), .A2(n465), .ZN(n466) );
  XNOR2_X2 U507 ( .A(n364), .B(n575), .ZN(n676) );
  NAND2_X1 U508 ( .A1(n574), .A2(n582), .ZN(n364) );
  XNOR2_X1 U509 ( .A(n367), .B(n607), .ZN(G57) );
  XNOR2_X1 U510 ( .A(n368), .B(n421), .ZN(G63) );
  NAND2_X1 U511 ( .A1(n423), .A2(n422), .ZN(n368) );
  XNOR2_X1 U512 ( .A(n693), .B(n692), .ZN(n370) );
  XNOR2_X1 U513 ( .A(n371), .B(n690), .ZN(G51) );
  NOR2_X2 U514 ( .A1(n733), .A2(n730), .ZN(n429) );
  XNOR2_X2 U515 ( .A(n375), .B(n599), .ZN(n638) );
  AND2_X2 U516 ( .A1(n419), .A2(n597), .ZN(n375) );
  XNOR2_X1 U517 ( .A(n379), .B(n378), .ZN(n377) );
  INV_X1 U518 ( .A(KEYINPUT47), .ZN(n378) );
  XNOR2_X1 U519 ( .A(n539), .B(KEYINPUT36), .ZN(n381) );
  NOR2_X4 U520 ( .A1(n644), .A2(n387), .ZN(n703) );
  NAND2_X1 U521 ( .A1(n390), .A2(n389), .ZN(n388) );
  NAND2_X1 U522 ( .A1(n571), .A2(n393), .ZN(n392) );
  XNOR2_X2 U523 ( .A(n565), .B(n566), .ZN(n571) );
  XOR2_X2 U524 ( .A(G101), .B(G113), .Z(n468) );
  XNOR2_X2 U525 ( .A(n468), .B(n467), .ZN(n484) );
  NOR2_X2 U526 ( .A1(n580), .A2(KEYINPUT73), .ZN(n579) );
  XNOR2_X2 U527 ( .A(G143), .B(G128), .ZN(n512) );
  NAND2_X1 U528 ( .A1(n412), .A2(n409), .ZN(n534) );
  INV_X1 U529 ( .A(n533), .ZN(n408) );
  NAND2_X1 U530 ( .A1(n693), .A2(n415), .ZN(n414) );
  XNOR2_X1 U531 ( .A(n579), .B(KEYINPUT44), .ZN(n419) );
  INV_X1 U532 ( .A(n567), .ZN(n645) );
  INV_X1 U533 ( .A(n465), .ZN(n586) );
  NAND2_X1 U534 ( .A1(n505), .A2(G221), .ZN(n449) );
  NOR2_X1 U535 ( .A1(n591), .A2(n662), .ZN(n564) );
  XNOR2_X1 U536 ( .A(n455), .B(n454), .ZN(n705) );
  NOR2_X1 U537 ( .A1(G902), .A2(n696), .ZN(n504) );
  XOR2_X2 U538 ( .A(G119), .B(G110), .Z(n481) );
  INV_X1 U539 ( .A(n512), .ZN(n514) );
  XNOR2_X1 U540 ( .A(n449), .B(n430), .ZN(n451) );
  XNOR2_X2 U541 ( .A(n450), .B(KEYINPUT10), .ZN(n719) );
  XOR2_X1 U542 ( .A(n448), .B(n447), .Z(n430) );
  XOR2_X1 U543 ( .A(n472), .B(n473), .Z(n431) );
  INV_X1 U544 ( .A(n497), .ZN(n482) );
  XNOR2_X1 U545 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U546 ( .A(n451), .B(n719), .ZN(n455) );
  XNOR2_X1 U547 ( .A(n605), .B(n604), .ZN(n606) );
  INV_X1 U548 ( .A(KEYINPUT63), .ZN(n607) );
  XOR2_X1 U549 ( .A(KEYINPUT14), .B(KEYINPUT87), .Z(n433) );
  XNOR2_X1 U550 ( .A(n433), .B(n432), .ZN(n434) );
  NAND2_X1 U551 ( .A1(G952), .A2(n434), .ZN(n673) );
  NOR2_X1 U552 ( .A1(G953), .A2(n673), .ZN(n559) );
  NAND2_X1 U553 ( .A1(G902), .A2(n434), .ZN(n435) );
  XOR2_X1 U554 ( .A(KEYINPUT88), .B(n435), .Z(n436) );
  NAND2_X1 U555 ( .A1(G953), .A2(n436), .ZN(n557) );
  NOR2_X1 U556 ( .A1(G900), .A2(n557), .ZN(n437) );
  XNOR2_X1 U557 ( .A(n437), .B(KEYINPUT108), .ZN(n438) );
  NOR2_X1 U558 ( .A1(n559), .A2(n438), .ZN(n521) );
  XOR2_X1 U559 ( .A(KEYINPUT91), .B(G110), .Z(n440) );
  XNOR2_X1 U560 ( .A(G107), .B(G101), .ZN(n439) );
  XNOR2_X1 U561 ( .A(n440), .B(n439), .ZN(n444) );
  NAND2_X1 U562 ( .A1(G227), .A2(n723), .ZN(n442) );
  XNOR2_X1 U563 ( .A(n446), .B(n720), .ZN(n693) );
  XOR2_X1 U564 ( .A(KEYINPUT93), .B(KEYINPUT92), .Z(n448) );
  XNOR2_X1 U565 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n447) );
  XNOR2_X1 U566 ( .A(G128), .B(n481), .ZN(n453) );
  NAND2_X1 U567 ( .A1(G234), .A2(n601), .ZN(n456) );
  NAND2_X1 U568 ( .A1(G217), .A2(n462), .ZN(n459) );
  INV_X1 U569 ( .A(KEYINPUT25), .ZN(n458) );
  XNOR2_X2 U570 ( .A(n461), .B(n460), .ZN(n567) );
  NAND2_X1 U571 ( .A1(G221), .A2(n462), .ZN(n464) );
  XNOR2_X1 U572 ( .A(KEYINPUT96), .B(KEYINPUT21), .ZN(n463) );
  XOR2_X1 U573 ( .A(n464), .B(n463), .Z(n646) );
  XNOR2_X1 U574 ( .A(n466), .B(KEYINPUT78), .ZN(n479) );
  XOR2_X1 U575 ( .A(KEYINPUT30), .B(KEYINPUT110), .Z(n477) );
  XNOR2_X1 U576 ( .A(n470), .B(n469), .ZN(n473) );
  XNOR2_X1 U577 ( .A(n471), .B(KEYINPUT76), .ZN(n496) );
  NAND2_X1 U578 ( .A1(G210), .A2(n496), .ZN(n472) );
  XNOR2_X2 U579 ( .A(n475), .B(G472), .ZN(n649) );
  NAND2_X1 U580 ( .A1(G214), .A2(n492), .ZN(n659) );
  NAND2_X1 U581 ( .A1(n589), .A2(n659), .ZN(n476) );
  XNOR2_X1 U582 ( .A(n477), .B(n476), .ZN(n478) );
  NAND2_X1 U583 ( .A1(n479), .A2(n478), .ZN(n548) );
  XNOR2_X1 U584 ( .A(KEYINPUT74), .B(KEYINPUT16), .ZN(n480) );
  XOR2_X1 U585 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n486) );
  XNOR2_X1 U586 ( .A(KEYINPUT79), .B(KEYINPUT86), .ZN(n485) );
  XNOR2_X1 U587 ( .A(n486), .B(n485), .ZN(n488) );
  NAND2_X1 U588 ( .A1(G224), .A2(n723), .ZN(n491) );
  NAND2_X1 U589 ( .A1(n684), .A2(n601), .ZN(n493) );
  XNOR2_X2 U590 ( .A(n493), .B(n353), .ZN(n544) );
  INV_X1 U591 ( .A(n660), .ZN(n494) );
  NOR2_X2 U592 ( .A1(n548), .A2(n494), .ZN(n495) );
  XNOR2_X1 U593 ( .A(n495), .B(KEYINPUT39), .ZN(n530) );
  NAND2_X1 U594 ( .A1(n496), .A2(G214), .ZN(n503) );
  XNOR2_X1 U595 ( .A(n497), .B(KEYINPUT11), .ZN(n502) );
  XOR2_X1 U596 ( .A(KEYINPUT12), .B(KEYINPUT98), .Z(n501) );
  XNOR2_X1 U597 ( .A(n499), .B(n498), .ZN(n500) );
  NAND2_X1 U598 ( .A1(n505), .A2(G217), .ZN(n518) );
  XNOR2_X1 U599 ( .A(n507), .B(n506), .ZN(n511) );
  XNOR2_X1 U600 ( .A(n509), .B(n508), .ZN(n510) );
  XOR2_X1 U601 ( .A(n511), .B(n510), .Z(n516) );
  XNOR2_X1 U602 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U603 ( .A(n516), .B(n515), .ZN(n517) );
  NOR2_X1 U604 ( .A1(G902), .A2(n702), .ZN(n519) );
  XOR2_X1 U605 ( .A(G478), .B(n519), .Z(n524) );
  NAND2_X1 U606 ( .A1(n529), .A2(n524), .ZN(n617) );
  NOR2_X1 U607 ( .A1(n530), .A2(n617), .ZN(n635) );
  XOR2_X1 U608 ( .A(KEYINPUT112), .B(KEYINPUT42), .Z(n528) );
  NAND2_X1 U609 ( .A1(n646), .A2(n567), .ZN(n520) );
  NOR2_X1 U610 ( .A1(n521), .A2(n520), .ZN(n538) );
  AND2_X1 U611 ( .A1(n538), .A2(n589), .ZN(n522) );
  XOR2_X1 U612 ( .A(KEYINPUT28), .B(n522), .Z(n523) );
  NOR2_X1 U613 ( .A1(n534), .A2(n523), .ZN(n543) );
  INV_X1 U614 ( .A(n524), .ZN(n546) );
  NAND2_X1 U615 ( .A1(n547), .A2(n546), .ZN(n662) );
  NAND2_X1 U616 ( .A1(n660), .A2(n659), .ZN(n663) );
  NOR2_X1 U617 ( .A1(n662), .A2(n663), .ZN(n526) );
  XNOR2_X1 U618 ( .A(KEYINPUT111), .B(KEYINPUT41), .ZN(n525) );
  XNOR2_X1 U619 ( .A(n526), .B(n525), .ZN(n675) );
  NAND2_X1 U620 ( .A1(n543), .A2(n675), .ZN(n527) );
  XNOR2_X1 U621 ( .A(n528), .B(n527), .ZN(n730) );
  NOR2_X1 U622 ( .A1(n530), .A2(n623), .ZN(n531) );
  XNOR2_X1 U623 ( .A(KEYINPUT46), .B(KEYINPUT84), .ZN(n532) );
  XNOR2_X1 U624 ( .A(KEYINPUT67), .B(KEYINPUT1), .ZN(n533) );
  INV_X1 U625 ( .A(n650), .ZN(n569) );
  XNOR2_X1 U626 ( .A(KEYINPUT6), .B(KEYINPUT105), .ZN(n535) );
  INV_X1 U627 ( .A(n582), .ZN(n536) );
  NOR2_X1 U628 ( .A1(n623), .A2(n536), .ZN(n537) );
  NAND2_X1 U629 ( .A1(n538), .A2(n537), .ZN(n551) );
  NAND2_X1 U630 ( .A1(n544), .A2(n659), .ZN(n541) );
  NOR2_X1 U631 ( .A1(n551), .A2(n541), .ZN(n539) );
  INV_X1 U632 ( .A(KEYINPUT19), .ZN(n540) );
  INV_X1 U633 ( .A(n561), .ZN(n542) );
  NAND2_X1 U634 ( .A1(n543), .A2(n542), .ZN(n622) );
  INV_X1 U635 ( .A(n623), .ZN(n626) );
  INV_X1 U636 ( .A(n617), .ZN(n628) );
  BUF_X1 U637 ( .A(n544), .Z(n545) );
  OR2_X1 U638 ( .A1(n547), .A2(n546), .ZN(n577) );
  NOR2_X1 U639 ( .A1(n548), .A2(n577), .ZN(n549) );
  NAND2_X1 U640 ( .A1(n545), .A2(n549), .ZN(n621) );
  XOR2_X1 U641 ( .A(KEYINPUT43), .B(KEYINPUT109), .Z(n554) );
  NOR2_X1 U642 ( .A1(n650), .A2(n551), .ZN(n552) );
  NAND2_X1 U643 ( .A1(n552), .A2(n659), .ZN(n553) );
  XNOR2_X1 U644 ( .A(n554), .B(n553), .ZN(n556) );
  INV_X1 U645 ( .A(n545), .ZN(n555) );
  NAND2_X1 U646 ( .A1(n556), .A2(n555), .ZN(n636) );
  XOR2_X1 U647 ( .A(KEYINPUT66), .B(KEYINPUT22), .Z(n566) );
  NOR2_X1 U648 ( .A1(G898), .A2(n557), .ZN(n558) );
  NOR2_X1 U649 ( .A1(n559), .A2(n558), .ZN(n560) );
  NOR2_X2 U650 ( .A1(n561), .A2(n560), .ZN(n563) );
  XNOR2_X2 U651 ( .A(n563), .B(n562), .ZN(n591) );
  NAND2_X1 U652 ( .A1(n564), .A2(n646), .ZN(n565) );
  NAND2_X1 U653 ( .A1(n569), .A2(n571), .ZN(n581) );
  NAND2_X1 U654 ( .A1(n567), .A2(n649), .ZN(n568) );
  NOR2_X1 U655 ( .A1(n581), .A2(n568), .ZN(n616) );
  NOR2_X1 U656 ( .A1(n569), .A2(n645), .ZN(n570) );
  XNOR2_X1 U657 ( .A(KEYINPUT106), .B(n570), .ZN(n572) );
  NOR2_X1 U658 ( .A1(n616), .A2(n732), .ZN(n578) );
  XOR2_X1 U659 ( .A(KEYINPUT107), .B(KEYINPUT33), .Z(n575) );
  INV_X1 U660 ( .A(n573), .ZN(n651) );
  INV_X1 U661 ( .A(n590), .ZN(n574) );
  NAND2_X1 U662 ( .A1(n585), .A2(n676), .ZN(n576) );
  NAND2_X1 U663 ( .A1(n578), .A2(n731), .ZN(n580) );
  NAND2_X1 U664 ( .A1(n580), .A2(KEYINPUT73), .ZN(n584) );
  NOR2_X1 U665 ( .A1(n582), .A2(n581), .ZN(n583) );
  NAND2_X1 U666 ( .A1(n583), .A2(n645), .ZN(n608) );
  NAND2_X1 U667 ( .A1(n584), .A2(n608), .ZN(n596) );
  NAND2_X1 U668 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U669 ( .A(KEYINPUT97), .B(n587), .Z(n588) );
  NOR2_X1 U670 ( .A1(n589), .A2(n588), .ZN(n613) );
  NOR2_X1 U671 ( .A1(n649), .A2(n590), .ZN(n656) );
  INV_X1 U672 ( .A(n591), .ZN(n592) );
  NAND2_X1 U673 ( .A1(n656), .A2(n592), .ZN(n593) );
  XNOR2_X1 U674 ( .A(KEYINPUT31), .B(n593), .ZN(n629) );
  NOR2_X1 U675 ( .A1(n613), .A2(n629), .ZN(n594) );
  NOR2_X1 U676 ( .A1(n664), .A2(n594), .ZN(n595) );
  NOR2_X1 U677 ( .A1(n596), .A2(n595), .ZN(n597) );
  INV_X1 U678 ( .A(KEYINPUT65), .ZN(n598) );
  INV_X1 U679 ( .A(KEYINPUT2), .ZN(n639) );
  OR2_X1 U680 ( .A1(n601), .A2(n639), .ZN(n600) );
  NAND2_X1 U681 ( .A1(n703), .A2(G472), .ZN(n605) );
  XOR2_X1 U682 ( .A(KEYINPUT113), .B(KEYINPUT62), .Z(n602) );
  XNOR2_X1 U683 ( .A(G101), .B(n608), .ZN(G3) );
  NAND2_X1 U684 ( .A1(n613), .A2(n626), .ZN(n609) );
  XNOR2_X1 U685 ( .A(n609), .B(G104), .ZN(G6) );
  XOR2_X1 U686 ( .A(KEYINPUT27), .B(KEYINPUT115), .Z(n611) );
  XNOR2_X1 U687 ( .A(G107), .B(KEYINPUT114), .ZN(n610) );
  XNOR2_X1 U688 ( .A(n611), .B(n610), .ZN(n612) );
  XOR2_X1 U689 ( .A(KEYINPUT26), .B(n612), .Z(n615) );
  NAND2_X1 U690 ( .A1(n613), .A2(n628), .ZN(n614) );
  XNOR2_X1 U691 ( .A(n615), .B(n614), .ZN(G9) );
  XOR2_X1 U692 ( .A(G110), .B(n616), .Z(G12) );
  NOR2_X1 U693 ( .A1(n617), .A2(n622), .ZN(n619) );
  XNOR2_X1 U694 ( .A(KEYINPUT116), .B(KEYINPUT29), .ZN(n618) );
  XNOR2_X1 U695 ( .A(n619), .B(n618), .ZN(n620) );
  XNOR2_X1 U696 ( .A(G128), .B(n620), .ZN(G30) );
  XNOR2_X1 U697 ( .A(G143), .B(n621), .ZN(G45) );
  NOR2_X1 U698 ( .A1(n623), .A2(n622), .ZN(n625) );
  XNOR2_X1 U699 ( .A(G146), .B(KEYINPUT117), .ZN(n624) );
  XNOR2_X1 U700 ( .A(n625), .B(n624), .ZN(G48) );
  NAND2_X1 U701 ( .A1(n629), .A2(n626), .ZN(n627) );
  XNOR2_X1 U702 ( .A(n627), .B(G113), .ZN(G15) );
  NAND2_X1 U703 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U704 ( .A(n630), .B(KEYINPUT118), .ZN(n631) );
  XNOR2_X1 U705 ( .A(G116), .B(n631), .ZN(G18) );
  XOR2_X1 U706 ( .A(KEYINPUT119), .B(KEYINPUT37), .Z(n634) );
  XNOR2_X1 U707 ( .A(G125), .B(n632), .ZN(n633) );
  XNOR2_X1 U708 ( .A(n634), .B(n633), .ZN(G27) );
  XOR2_X1 U709 ( .A(G134), .B(n635), .Z(G36) );
  XNOR2_X1 U710 ( .A(G140), .B(n636), .ZN(G42) );
  XOR2_X1 U711 ( .A(KEYINPUT53), .B(KEYINPUT122), .Z(n683) );
  NAND2_X1 U712 ( .A1(n722), .A2(n639), .ZN(n637) );
  XNOR2_X1 U713 ( .A(n637), .B(KEYINPUT82), .ZN(n641) );
  NAND2_X1 U714 ( .A1(n639), .A2(n638), .ZN(n640) );
  NAND2_X1 U715 ( .A1(n641), .A2(n640), .ZN(n642) );
  XOR2_X1 U716 ( .A(KEYINPUT81), .B(n642), .Z(n643) );
  NOR2_X1 U717 ( .A1(n349), .A2(n643), .ZN(n680) );
  NOR2_X1 U718 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U719 ( .A(n647), .B(KEYINPUT49), .ZN(n648) );
  NAND2_X1 U720 ( .A1(n649), .A2(n648), .ZN(n654) );
  NOR2_X1 U721 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U722 ( .A(n652), .B(KEYINPUT50), .ZN(n653) );
  NOR2_X1 U723 ( .A1(n654), .A2(n653), .ZN(n655) );
  NOR2_X1 U724 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U725 ( .A(n657), .B(KEYINPUT51), .ZN(n658) );
  NAND2_X1 U726 ( .A1(n658), .A2(n675), .ZN(n670) );
  NOR2_X1 U727 ( .A1(n660), .A2(n659), .ZN(n661) );
  NOR2_X1 U728 ( .A1(n662), .A2(n661), .ZN(n667) );
  NOR2_X1 U729 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U730 ( .A(KEYINPUT120), .B(n665), .ZN(n666) );
  OR2_X1 U731 ( .A1(n667), .A2(n666), .ZN(n668) );
  NAND2_X1 U732 ( .A1(n676), .A2(n668), .ZN(n669) );
  NAND2_X1 U733 ( .A1(n670), .A2(n669), .ZN(n671) );
  XOR2_X1 U734 ( .A(KEYINPUT52), .B(n671), .Z(n672) );
  NOR2_X1 U735 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U736 ( .A(n674), .B(KEYINPUT121), .ZN(n678) );
  NAND2_X1 U737 ( .A1(n676), .A2(n675), .ZN(n677) );
  NAND2_X1 U738 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U739 ( .A1(n680), .A2(n679), .ZN(n681) );
  NAND2_X1 U740 ( .A1(n681), .A2(n723), .ZN(n682) );
  XNOR2_X1 U741 ( .A(n683), .B(n682), .ZN(G75) );
  NAND2_X1 U742 ( .A1(n703), .A2(G210), .ZN(n688) );
  INV_X1 U743 ( .A(n684), .ZN(n686) );
  XOR2_X1 U744 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n685) );
  XNOR2_X1 U745 ( .A(n688), .B(n687), .ZN(n689) );
  XOR2_X1 U746 ( .A(KEYINPUT83), .B(KEYINPUT56), .Z(n690) );
  XOR2_X1 U747 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n692) );
  NAND2_X1 U748 ( .A1(n703), .A2(G469), .ZN(n691) );
  NOR2_X1 U749 ( .A1(n707), .A2(n694), .ZN(G54) );
  NAND2_X1 U750 ( .A1(n703), .A2(G475), .ZN(n698) );
  XOR2_X1 U751 ( .A(KEYINPUT59), .B(KEYINPUT68), .Z(n695) );
  XNOR2_X1 U752 ( .A(n698), .B(n697), .ZN(n699) );
  XOR2_X1 U753 ( .A(KEYINPUT60), .B(KEYINPUT123), .Z(n700) );
  XNOR2_X1 U754 ( .A(n701), .B(n700), .ZN(G60) );
  NAND2_X1 U755 ( .A1(G217), .A2(n703), .ZN(n704) );
  XNOR2_X1 U756 ( .A(n705), .B(n704), .ZN(n706) );
  NOR2_X1 U757 ( .A1(n707), .A2(n706), .ZN(G66) );
  XOR2_X1 U758 ( .A(n708), .B(KEYINPUT75), .Z(n709) );
  XNOR2_X1 U759 ( .A(KEYINPUT126), .B(n709), .ZN(n711) );
  NOR2_X1 U760 ( .A1(G898), .A2(n723), .ZN(n710) );
  NOR2_X1 U761 ( .A1(n711), .A2(n710), .ZN(n718) );
  NOR2_X1 U762 ( .A1(G953), .A2(n638), .ZN(n712) );
  XNOR2_X1 U763 ( .A(n712), .B(KEYINPUT125), .ZN(n716) );
  NAND2_X1 U764 ( .A1(G953), .A2(G224), .ZN(n713) );
  XNOR2_X1 U765 ( .A(KEYINPUT61), .B(n713), .ZN(n714) );
  NAND2_X1 U766 ( .A1(n714), .A2(G898), .ZN(n715) );
  NAND2_X1 U767 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U768 ( .A(n718), .B(n717), .ZN(G69) );
  XOR2_X1 U769 ( .A(n720), .B(n719), .Z(n725) );
  XOR2_X1 U770 ( .A(KEYINPUT127), .B(n725), .Z(n721) );
  XNOR2_X1 U771 ( .A(n722), .B(n721), .ZN(n724) );
  NAND2_X1 U772 ( .A1(n724), .A2(n723), .ZN(n729) );
  XNOR2_X1 U773 ( .A(G227), .B(n725), .ZN(n726) );
  NAND2_X1 U774 ( .A1(n726), .A2(G900), .ZN(n727) );
  NAND2_X1 U775 ( .A1(n727), .A2(G953), .ZN(n728) );
  NAND2_X1 U776 ( .A1(n729), .A2(n728), .ZN(G72) );
  XOR2_X1 U777 ( .A(n730), .B(G137), .Z(G39) );
  XNOR2_X1 U778 ( .A(n731), .B(G122), .ZN(G24) );
  XOR2_X1 U779 ( .A(n732), .B(G119), .Z(G21) );
  XOR2_X1 U780 ( .A(n733), .B(G131), .Z(G33) );
endmodule

