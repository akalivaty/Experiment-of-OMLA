//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 1 0 0 1 0 1 0 1 1 1 1 1 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 0 0 1 0 1 0 1 1 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:26 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n663, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n905,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968;
  INV_X1    g000(.A(G128), .ZN(new_n187));
  OAI21_X1  g001(.A(KEYINPUT23), .B1(new_n187), .B2(G119), .ZN(new_n188));
  INV_X1    g002(.A(G119), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(G128), .ZN(new_n190));
  MUX2_X1   g004(.A(new_n188), .B(KEYINPUT23), .S(new_n190), .Z(new_n191));
  XNOR2_X1  g005(.A(G119), .B(G128), .ZN(new_n192));
  XOR2_X1   g006(.A(KEYINPUT24), .B(G110), .Z(new_n193));
  OAI22_X1  g007(.A1(new_n191), .A2(G110), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G140), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G125), .ZN(new_n196));
  INV_X1    g010(.A(G125), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G140), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n196), .A2(new_n198), .A3(KEYINPUT16), .ZN(new_n199));
  OR3_X1    g013(.A1(new_n197), .A2(KEYINPUT16), .A3(G140), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n199), .A2(new_n200), .A3(G146), .ZN(new_n201));
  AND2_X1   g015(.A1(new_n196), .A2(new_n198), .ZN(new_n202));
  INV_X1    g016(.A(G146), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n194), .A2(new_n201), .A3(new_n204), .ZN(new_n205));
  AOI22_X1  g019(.A1(new_n191), .A2(G110), .B1(new_n192), .B2(new_n193), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n199), .A2(new_n200), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(new_n203), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(new_n201), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n206), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n205), .A2(new_n210), .ZN(new_n211));
  XNOR2_X1  g025(.A(KEYINPUT22), .B(G137), .ZN(new_n212));
  INV_X1    g026(.A(G221), .ZN(new_n213));
  INV_X1    g027(.A(G234), .ZN(new_n214));
  NOR3_X1   g028(.A1(new_n213), .A2(new_n214), .A3(G953), .ZN(new_n215));
  XOR2_X1   g029(.A(new_n212), .B(new_n215), .Z(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n211), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G902), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT72), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT25), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n205), .A2(new_n210), .A3(new_n216), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n218), .A2(new_n219), .A3(new_n222), .A4(new_n223), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n220), .A2(new_n221), .ZN(new_n225));
  OR2_X1    g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n224), .A2(new_n225), .ZN(new_n227));
  OAI21_X1  g041(.A(G217), .B1(new_n214), .B2(G902), .ZN(new_n228));
  XNOR2_X1  g042(.A(new_n228), .B(KEYINPUT71), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n226), .A2(new_n227), .A3(new_n229), .ZN(new_n230));
  AND2_X1   g044(.A1(new_n218), .A2(new_n223), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n228), .A2(new_n219), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n230), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT30), .ZN(new_n236));
  INV_X1    g050(.A(G137), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n237), .A2(G134), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(KEYINPUT65), .ZN(new_n239));
  INV_X1    g053(.A(G134), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G137), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT65), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  OAI211_X1 g057(.A(new_n239), .B(new_n243), .C1(new_n240), .C2(G137), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G131), .ZN(new_n245));
  OAI21_X1  g059(.A(KEYINPUT11), .B1(new_n240), .B2(G137), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT11), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n247), .A2(new_n237), .A3(G134), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(G131), .ZN(new_n250));
  AND4_X1   g064(.A1(KEYINPUT64), .A2(new_n249), .A3(new_n250), .A4(new_n241), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n238), .B1(new_n246), .B2(new_n248), .ZN(new_n252));
  AOI21_X1  g066(.A(KEYINPUT64), .B1(new_n252), .B2(new_n250), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n245), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n203), .A2(G143), .ZN(new_n255));
  INV_X1    g069(.A(G143), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G146), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT1), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n255), .A2(new_n257), .A3(new_n258), .A4(G128), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  OAI21_X1  g074(.A(KEYINPUT1), .B1(new_n256), .B2(G146), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(KEYINPUT66), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT66), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n255), .A2(new_n263), .A3(KEYINPUT1), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n262), .A2(G128), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n255), .A2(new_n257), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n260), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n254), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT0), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n269), .A2(new_n187), .ZN(new_n270));
  NOR2_X1   g084(.A1(KEYINPUT0), .A2(G128), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n266), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  XNOR2_X1  g086(.A(G143), .B(G146), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n273), .B1(new_n269), .B2(new_n187), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n249), .A2(new_n250), .A3(new_n241), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT64), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n252), .A2(KEYINPUT64), .A3(new_n250), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  OR2_X1    g095(.A1(new_n252), .A2(new_n250), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n276), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n236), .B1(new_n268), .B2(new_n283), .ZN(new_n284));
  XOR2_X1   g098(.A(G116), .B(G119), .Z(new_n285));
  XNOR2_X1  g099(.A(KEYINPUT2), .B(G113), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  XOR2_X1   g101(.A(KEYINPUT2), .B(G113), .Z(new_n288));
  XNOR2_X1  g102(.A(G116), .B(G119), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n287), .A2(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n282), .B1(new_n251), .B2(new_n253), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(new_n275), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n265), .A2(new_n266), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(new_n259), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n281), .A2(new_n295), .A3(new_n245), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n293), .A2(new_n296), .A3(KEYINPUT30), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n284), .A2(new_n291), .A3(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n291), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n293), .A2(new_n296), .A3(new_n299), .ZN(new_n300));
  XNOR2_X1  g114(.A(KEYINPUT67), .B(G237), .ZN(new_n301));
  INV_X1    g115(.A(G953), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n301), .A2(G210), .A3(new_n302), .ZN(new_n303));
  XNOR2_X1  g117(.A(KEYINPUT26), .B(G101), .ZN(new_n304));
  XOR2_X1   g118(.A(new_n303), .B(new_n304), .Z(new_n305));
  XNOR2_X1  g119(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n305), .B(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n298), .A2(new_n300), .A3(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT31), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n298), .A2(KEYINPUT31), .A3(new_n308), .A4(new_n300), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AND3_X1   g127(.A1(new_n293), .A2(new_n296), .A3(new_n299), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n299), .B1(new_n293), .B2(new_n296), .ZN(new_n315));
  OAI21_X1  g129(.A(KEYINPUT28), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT28), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n300), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n308), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  AOI21_X1  g134(.A(G902), .B1(new_n313), .B2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(G472), .ZN(new_n322));
  AOI21_X1  g136(.A(KEYINPUT32), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n319), .B1(new_n311), .B2(new_n312), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT32), .ZN(new_n325));
  NOR4_X1   g139(.A1(new_n324), .A2(new_n325), .A3(G472), .A4(G902), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n323), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n316), .A2(new_n308), .A3(new_n318), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT29), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(KEYINPUT69), .ZN(new_n330));
  XNOR2_X1  g144(.A(new_n328), .B(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT70), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n298), .A2(new_n300), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n332), .B1(new_n333), .B2(new_n307), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n333), .A2(new_n332), .A3(new_n307), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n331), .B1(new_n329), .B2(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(G472), .B1(new_n338), .B2(G902), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n235), .B1(new_n327), .B2(new_n339), .ZN(new_n340));
  OAI21_X1  g154(.A(G214), .B1(G237), .B2(G902), .ZN(new_n341));
  INV_X1    g155(.A(G101), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT3), .ZN(new_n343));
  INV_X1    g157(.A(G104), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n343), .B1(new_n344), .B2(G107), .ZN(new_n345));
  INV_X1    g159(.A(G107), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n346), .A2(KEYINPUT3), .A3(G104), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n344), .A2(G107), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n342), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT4), .ZN(new_n351));
  AOI22_X1  g165(.A1(new_n350), .A2(new_n351), .B1(new_n287), .B2(new_n290), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n348), .A2(new_n349), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(G101), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n348), .A2(new_n342), .A3(new_n349), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n354), .A2(KEYINPUT4), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n352), .A2(new_n356), .ZN(new_n357));
  XOR2_X1   g171(.A(G110), .B(G122), .Z(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n289), .A2(KEYINPUT5), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT5), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n361), .A2(new_n189), .A3(G116), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT76), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n361), .A2(new_n189), .A3(KEYINPUT76), .A4(G116), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n360), .A2(G113), .A3(new_n364), .A4(new_n365), .ZN(new_n366));
  OAI21_X1  g180(.A(KEYINPUT73), .B1(new_n344), .B2(G107), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT74), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n368), .B1(new_n346), .B2(G104), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT73), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n370), .A2(new_n346), .A3(G104), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n344), .A2(KEYINPUT74), .A3(G107), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n367), .A2(new_n369), .A3(new_n371), .A4(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(G101), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n366), .A2(new_n290), .A3(new_n374), .A4(new_n355), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n357), .A2(new_n359), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n366), .A2(new_n290), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n374), .A2(new_n355), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT80), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n378), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n364), .A2(G113), .A3(new_n365), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(KEYINPUT79), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT79), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n364), .A2(new_n385), .A3(G113), .A4(new_n365), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n384), .A2(new_n360), .A3(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n382), .A2(new_n387), .A3(new_n290), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n377), .A2(KEYINPUT80), .A3(new_n378), .ZN(new_n389));
  AND3_X1   g203(.A1(new_n381), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n358), .B(KEYINPUT8), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n376), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n275), .A2(G125), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n393), .B1(new_n267), .B2(G125), .ZN(new_n394));
  NAND2_X1  g208(.A1(KEYINPUT81), .A2(KEYINPUT7), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n302), .A2(G224), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(KEYINPUT7), .ZN(new_n398));
  XNOR2_X1  g212(.A(new_n396), .B(new_n398), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n219), .B1(new_n392), .B2(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(G210), .B1(G237), .B2(G902), .ZN(new_n401));
  XNOR2_X1  g215(.A(new_n401), .B(KEYINPUT82), .ZN(new_n402));
  AND3_X1   g216(.A1(new_n348), .A2(new_n342), .A3(new_n349), .ZN(new_n403));
  NOR3_X1   g217(.A1(new_n403), .A2(new_n350), .A3(new_n351), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n353), .A2(new_n351), .A3(G101), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n291), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n375), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(new_n358), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n408), .A2(KEYINPUT6), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT77), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n410), .B1(new_n408), .B2(new_n376), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n359), .B1(new_n357), .B2(new_n375), .ZN(new_n412));
  OAI21_X1  g226(.A(KEYINPUT6), .B1(new_n412), .B2(KEYINPUT77), .ZN(new_n413));
  OAI21_X1  g227(.A(KEYINPUT78), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n407), .A2(new_n358), .ZN(new_n415));
  OAI21_X1  g229(.A(KEYINPUT77), .B1(new_n415), .B2(new_n412), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT78), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT6), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n418), .B1(new_n408), .B2(new_n410), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n416), .A2(new_n417), .A3(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n409), .B1(new_n414), .B2(new_n420), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n394), .B(new_n397), .ZN(new_n422));
  AOI211_X1 g236(.A(new_n400), .B(new_n402), .C1(new_n421), .C2(new_n422), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n402), .B(KEYINPUT83), .ZN(new_n424));
  INV_X1    g238(.A(new_n409), .ZN(new_n425));
  NOR3_X1   g239(.A1(new_n411), .A2(new_n413), .A3(KEYINPUT78), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n417), .B1(new_n416), .B2(new_n419), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n425), .B(new_n422), .C1(new_n426), .C2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n400), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n424), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  OAI211_X1 g244(.A(KEYINPUT84), .B(new_n341), .C1(new_n423), .C2(new_n430), .ZN(new_n431));
  XNOR2_X1  g245(.A(G110), .B(G140), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n302), .A2(G227), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n432), .B(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n382), .A2(new_n295), .A3(KEYINPUT10), .ZN(new_n436));
  AOI22_X1  g250(.A1(new_n350), .A2(new_n351), .B1(new_n272), .B2(new_n274), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n356), .A2(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n187), .B1(new_n255), .B2(KEYINPUT1), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n259), .B1(new_n439), .B2(new_n273), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n374), .A2(new_n440), .A3(new_n355), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT10), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n436), .A2(new_n438), .A3(new_n443), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n444), .A2(new_n292), .ZN(new_n445));
  INV_X1    g259(.A(new_n292), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n442), .B1(new_n294), .B2(new_n259), .ZN(new_n447));
  AOI22_X1  g261(.A1(new_n447), .A2(new_n382), .B1(new_n356), .B2(new_n437), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n446), .B1(new_n448), .B2(new_n443), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n435), .B1(new_n445), .B2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(new_n441), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n451), .B1(new_n267), .B2(new_n378), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT75), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n292), .A2(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(KEYINPUT12), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n448), .A2(new_n446), .A3(new_n443), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n441), .B1(new_n382), .B2(new_n295), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT12), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n457), .A2(new_n453), .A3(new_n458), .A4(new_n292), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n455), .A2(new_n456), .A3(new_n459), .A4(new_n434), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n450), .A2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(G469), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n461), .A2(new_n462), .A3(new_n219), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n462), .A2(new_n219), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  AND3_X1   g279(.A1(new_n455), .A2(new_n456), .A3(new_n459), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n456), .A2(new_n434), .ZN(new_n467));
  OAI22_X1  g281(.A1(new_n466), .A2(new_n434), .B1(new_n449), .B2(new_n467), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n463), .B(new_n465), .C1(new_n462), .C2(new_n468), .ZN(new_n469));
  XOR2_X1   g283(.A(KEYINPUT9), .B(G234), .Z(new_n470));
  AOI21_X1  g284(.A(new_n213), .B1(new_n470), .B2(new_n219), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  AND2_X1   g286(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(G952), .ZN(new_n474));
  OR2_X1    g288(.A1(new_n474), .A2(KEYINPUT91), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(KEYINPUT91), .ZN(new_n476));
  AOI21_X1  g290(.A(G953), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(G234), .A2(G237), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  XOR2_X1   g294(.A(KEYINPUT21), .B(G898), .Z(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n478), .A2(G902), .A3(G953), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n480), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  AND3_X1   g300(.A1(new_n431), .A2(new_n473), .A3(new_n486), .ZN(new_n487));
  XNOR2_X1  g301(.A(G113), .B(G122), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n488), .B(new_n344), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  AND2_X1   g304(.A1(KEYINPUT67), .A2(G237), .ZN(new_n491));
  NOR2_X1   g305(.A1(KEYINPUT67), .A2(G237), .ZN(new_n492));
  OAI211_X1 g306(.A(G214), .B(new_n302), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(new_n256), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n301), .A2(G143), .A3(G214), .A4(new_n302), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n494), .A2(new_n495), .A3(new_n250), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(KEYINPUT86), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n494), .A2(new_n495), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(G131), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT86), .ZN(new_n500));
  NAND4_X1  g314(.A1(new_n494), .A2(new_n495), .A3(new_n500), .A4(new_n250), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n497), .A2(new_n499), .A3(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n201), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n202), .B(KEYINPUT19), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n503), .B1(new_n504), .B2(new_n203), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n494), .A2(new_n495), .A3(KEYINPUT85), .ZN(new_n507));
  NAND2_X1  g321(.A1(KEYINPUT18), .A2(G131), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n508), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n494), .A2(new_n495), .A3(KEYINPUT85), .A4(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n202), .B(new_n203), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n506), .A2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT17), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n497), .A2(new_n499), .A3(new_n516), .A4(new_n501), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n250), .B1(new_n494), .B2(new_n495), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n209), .B1(KEYINPUT17), .B2(new_n518), .ZN(new_n519));
  AOI22_X1  g333(.A1(new_n517), .A2(new_n519), .B1(new_n512), .B2(new_n513), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n489), .B(KEYINPUT87), .ZN(new_n521));
  AOI22_X1  g335(.A1(new_n490), .A2(new_n515), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g336(.A1(G475), .A2(G902), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  OAI21_X1  g338(.A(KEYINPUT88), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT88), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n517), .A2(new_n519), .ZN(new_n527));
  AND3_X1   g341(.A1(new_n527), .A2(new_n514), .A3(new_n521), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n489), .B1(new_n506), .B2(new_n514), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n526), .B(new_n523), .C1(new_n528), .C2(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n525), .A2(KEYINPUT20), .A3(new_n530), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n520), .A2(new_n489), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n219), .B1(new_n532), .B2(new_n528), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(G475), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT20), .ZN(new_n535));
  OAI211_X1 g349(.A(KEYINPUT88), .B(new_n535), .C1(new_n522), .C2(new_n524), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n531), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(KEYINPUT89), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT89), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n531), .A2(new_n539), .A3(new_n534), .A4(new_n536), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(G122), .ZN(new_n542));
  OAI21_X1  g356(.A(KEYINPUT14), .B1(new_n542), .B2(G116), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n543), .B(KEYINPUT90), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n542), .A2(G116), .ZN(new_n545));
  INV_X1    g359(.A(G116), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(G122), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n545), .B1(new_n547), .B2(KEYINPUT14), .ZN(new_n548));
  OAI21_X1  g362(.A(G107), .B1(new_n544), .B2(new_n548), .ZN(new_n549));
  AND2_X1   g363(.A1(new_n545), .A2(new_n547), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(new_n346), .ZN(new_n551));
  XNOR2_X1  g365(.A(G128), .B(G143), .ZN(new_n552));
  XNOR2_X1  g366(.A(new_n552), .B(new_n240), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n549), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n550), .B(new_n346), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n552), .A2(KEYINPUT13), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n256), .A2(G128), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n556), .B(G134), .C1(KEYINPUT13), .C2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n552), .A2(new_n240), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n555), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n554), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n470), .A2(G217), .A3(new_n302), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n562), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n554), .A2(new_n560), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(new_n219), .ZN(new_n567));
  INV_X1    g381(.A(G478), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n568), .A2(KEYINPUT15), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n567), .B(new_n569), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n541), .A2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT84), .ZN(new_n572));
  INV_X1    g386(.A(new_n402), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n428), .A2(new_n429), .A3(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n400), .B1(new_n421), .B2(new_n422), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n574), .B1(new_n575), .B2(new_n424), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n341), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n572), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n340), .A2(new_n487), .A3(new_n571), .A4(new_n579), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n580), .B(G101), .ZN(G3));
  XNOR2_X1  g395(.A(new_n566), .B(KEYINPUT33), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(G478), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n566), .A2(new_n568), .A3(new_n219), .ZN(new_n585));
  NAND2_X1  g399(.A1(G478), .A2(G902), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n541), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n422), .ZN(new_n590));
  AOI211_X1 g404(.A(new_n409), .B(new_n590), .C1(new_n414), .C2(new_n420), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n402), .B1(new_n591), .B2(new_n400), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(new_n574), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n593), .A2(new_n341), .A3(new_n486), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n589), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n313), .A2(new_n320), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n597), .A2(new_n322), .A3(new_n219), .ZN(new_n598));
  OAI21_X1  g412(.A(G472), .B1(new_n324), .B2(G902), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n600), .A2(new_n235), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(new_n473), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n596), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(KEYINPUT34), .B(G104), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n603), .B(new_n604), .ZN(G6));
  NAND4_X1  g419(.A1(new_n531), .A2(new_n570), .A3(new_n534), .A4(new_n536), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n594), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n608), .A2(new_n602), .ZN(new_n609));
  XNOR2_X1  g423(.A(KEYINPUT35), .B(G107), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n609), .B(new_n610), .ZN(G9));
  NOR2_X1   g425(.A1(new_n217), .A2(KEYINPUT36), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n211), .B(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(new_n233), .ZN(new_n614));
  AND2_X1   g428(.A1(new_n230), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n600), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n487), .A2(new_n571), .A3(new_n616), .A4(new_n579), .ZN(new_n617));
  XOR2_X1   g431(.A(KEYINPUT37), .B(G110), .Z(new_n618));
  XNOR2_X1  g432(.A(new_n617), .B(new_n618), .ZN(G12));
  AND3_X1   g433(.A1(new_n531), .A2(new_n534), .A3(new_n536), .ZN(new_n620));
  XOR2_X1   g434(.A(KEYINPUT92), .B(G900), .Z(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(new_n484), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n479), .A2(new_n622), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n620), .A2(KEYINPUT93), .A3(new_n570), .A4(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT93), .ZN(new_n625));
  INV_X1    g439(.A(new_n623), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n625), .B1(new_n606), .B2(new_n626), .ZN(new_n627));
  AND2_X1   g441(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n598), .A2(new_n325), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n321), .A2(KEYINPUT32), .A3(new_n322), .ZN(new_n630));
  INV_X1    g444(.A(new_n336), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n329), .B1(new_n631), .B2(new_n334), .ZN(new_n632));
  INV_X1    g446(.A(new_n330), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n328), .B(new_n633), .ZN(new_n634));
  AOI21_X1  g448(.A(G902), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  OAI211_X1 g449(.A(new_n629), .B(new_n630), .C1(new_n635), .C2(new_n322), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n230), .A2(new_n614), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n573), .B1(new_n428), .B2(new_n429), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n341), .B1(new_n423), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n469), .A2(new_n472), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n628), .A2(new_n636), .A3(new_n637), .A4(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(G128), .ZN(G30));
  XNOR2_X1  g457(.A(KEYINPUT94), .B(KEYINPUT38), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n577), .A2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n644), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n576), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n637), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n333), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n649), .A2(new_n307), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n314), .A2(new_n315), .ZN(new_n651));
  AOI21_X1  g465(.A(G902), .B1(new_n651), .B2(new_n307), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  OAI21_X1  g467(.A(G472), .B1(new_n650), .B2(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n629), .A2(new_n630), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n623), .B(KEYINPUT39), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n473), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(KEYINPUT40), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n648), .A2(new_n341), .A3(new_n655), .A4(new_n658), .ZN(new_n659));
  OAI211_X1 g473(.A(new_n570), .B(new_n541), .C1(new_n657), .C2(KEYINPUT40), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(new_n256), .ZN(G45));
  AOI211_X1 g476(.A(new_n626), .B(new_n587), .C1(new_n538), .C2(new_n540), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n636), .A2(new_n663), .A3(new_n637), .A4(new_n641), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G146), .ZN(G48));
  AOI21_X1  g479(.A(new_n462), .B1(new_n461), .B2(new_n219), .ZN(new_n666));
  AOI211_X1 g480(.A(G469), .B(G902), .C1(new_n450), .C2(new_n460), .ZN(new_n667));
  NOR3_X1   g481(.A1(new_n666), .A2(new_n667), .A3(new_n471), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT95), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n340), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n672), .A2(new_n596), .ZN(new_n673));
  XOR2_X1   g487(.A(KEYINPUT41), .B(G113), .Z(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G15));
  NOR2_X1   g489(.A1(new_n672), .A2(new_n608), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(new_n546), .ZN(G18));
  AOI21_X1  g491(.A(new_n615), .B1(new_n327), .B2(new_n339), .ZN(new_n678));
  OAI211_X1 g492(.A(new_n341), .B(new_n668), .C1(new_n423), .C2(new_n638), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(KEYINPUT96), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT96), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n593), .A2(new_n681), .A3(new_n341), .A4(new_n668), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n678), .A2(new_n683), .A3(new_n571), .A4(new_n486), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G119), .ZN(G21));
  NOR2_X1   g499(.A1(new_n670), .A2(new_n594), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n291), .B1(new_n268), .B2(new_n283), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n317), .B1(new_n687), .B2(new_n300), .ZN(new_n688));
  INV_X1    g502(.A(new_n318), .ZN(new_n689));
  OAI21_X1  g503(.A(KEYINPUT97), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT97), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n316), .A2(new_n691), .A3(new_n318), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n690), .A2(new_n692), .A3(new_n307), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n313), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g508(.A1(G472), .A2(G902), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AND2_X1   g510(.A1(new_n696), .A2(new_n599), .ZN(new_n697));
  INV_X1    g511(.A(new_n235), .ZN(new_n698));
  AND2_X1   g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT98), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n700), .B1(new_n541), .B2(new_n570), .ZN(new_n701));
  INV_X1    g515(.A(new_n570), .ZN(new_n702));
  AOI211_X1 g516(.A(KEYINPUT98), .B(new_n702), .C1(new_n538), .C2(new_n540), .ZN(new_n703));
  OAI211_X1 g517(.A(new_n686), .B(new_n699), .C1(new_n701), .C2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G122), .ZN(G24));
  AOI21_X1  g519(.A(new_n587), .B1(new_n538), .B2(new_n540), .ZN(new_n706));
  AND3_X1   g520(.A1(new_n696), .A2(new_n599), .A3(new_n637), .ZN(new_n707));
  AND3_X1   g521(.A1(new_n706), .A2(new_n707), .A3(new_n623), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n683), .ZN(new_n709));
  XOR2_X1   g523(.A(KEYINPUT99), .B(G125), .Z(new_n710));
  XNOR2_X1  g524(.A(new_n709), .B(new_n710), .ZN(G27));
  NOR2_X1   g525(.A1(KEYINPUT100), .A2(KEYINPUT42), .ZN(new_n712));
  OAI211_X1 g526(.A(new_n574), .B(new_n341), .C1(new_n575), .C2(new_n424), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n713), .A2(new_n640), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n629), .A2(new_n630), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n635), .A2(new_n322), .ZN(new_n716));
  OAI211_X1 g530(.A(new_n714), .B(new_n698), .C1(new_n715), .C2(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(new_n663), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n712), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(new_n712), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n340), .A2(new_n663), .A3(new_n714), .A4(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G131), .ZN(G33));
  INV_X1    g537(.A(new_n628), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n717), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(new_n240), .ZN(G36));
  NAND2_X1  g540(.A1(new_n600), .A2(new_n637), .ZN(new_n727));
  XOR2_X1   g541(.A(new_n727), .B(KEYINPUT103), .Z(new_n728));
  INV_X1    g542(.A(new_n541), .ZN(new_n729));
  OAI211_X1 g543(.A(new_n729), .B(new_n588), .C1(KEYINPUT102), .C2(KEYINPUT43), .ZN(new_n730));
  XNOR2_X1  g544(.A(KEYINPUT102), .B(KEYINPUT43), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n731), .B1(new_n541), .B2(new_n587), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  AND3_X1   g547(.A1(new_n728), .A2(KEYINPUT44), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g548(.A(KEYINPUT44), .B1(new_n728), .B2(new_n733), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n713), .B(KEYINPUT104), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  NOR3_X1   g551(.A1(new_n734), .A2(new_n735), .A3(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n468), .B(KEYINPUT45), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(G469), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(KEYINPUT101), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT101), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n739), .A2(new_n742), .A3(G469), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n464), .B1(new_n741), .B2(new_n743), .ZN(new_n744));
  OR2_X1    g558(.A1(new_n744), .A2(KEYINPUT46), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n667), .B1(new_n744), .B2(KEYINPUT46), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n471), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  AND2_X1   g561(.A1(new_n747), .A2(new_n656), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n738), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G137), .ZN(G39));
  NAND2_X1  g564(.A1(new_n744), .A2(KEYINPUT46), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(new_n463), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n744), .A2(KEYINPUT46), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n472), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(KEYINPUT47), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT47), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n747), .A2(new_n756), .ZN(new_n757));
  NOR3_X1   g571(.A1(new_n636), .A2(new_n698), .A3(new_n713), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n755), .A2(new_n757), .A3(new_n663), .A4(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G140), .ZN(G42));
  NAND2_X1  g574(.A1(new_n645), .A2(new_n647), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n698), .A2(new_n341), .A3(new_n472), .ZN(new_n762));
  OR2_X1    g576(.A1(new_n666), .A2(new_n667), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n762), .B1(KEYINPUT49), .B2(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n764), .A2(new_n729), .A3(new_n588), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT105), .ZN(new_n766));
  AOI211_X1 g580(.A(new_n655), .B(new_n761), .C1(new_n765), .C2(new_n766), .ZN(new_n767));
  OAI221_X1 g581(.A(new_n767), .B1(new_n766), .B2(new_n765), .C1(KEYINPUT49), .C2(new_n763), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n754), .A2(KEYINPUT47), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n747), .A2(new_n756), .ZN(new_n770));
  OAI22_X1  g584(.A1(new_n769), .A2(new_n770), .B1(new_n472), .B2(new_n763), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n699), .A2(new_n480), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n772), .B1(new_n730), .B2(new_n732), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT110), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n773), .A2(new_n774), .A3(new_n736), .ZN(new_n775));
  INV_X1    g589(.A(new_n775), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n774), .B1(new_n773), .B2(new_n736), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT111), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n771), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n763), .A2(new_n472), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n781), .B1(new_n755), .B2(new_n757), .ZN(new_n782));
  INV_X1    g596(.A(new_n777), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(new_n775), .ZN(new_n784));
  OAI21_X1  g598(.A(KEYINPUT111), .B1(new_n782), .B2(new_n784), .ZN(new_n785));
  NOR4_X1   g599(.A1(new_n713), .A2(new_n471), .A3(new_n479), .A4(new_n763), .ZN(new_n786));
  INV_X1    g600(.A(new_n655), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n786), .A2(new_n787), .A3(new_n698), .ZN(new_n788));
  NOR3_X1   g602(.A1(new_n788), .A2(new_n541), .A3(new_n588), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT113), .ZN(new_n790));
  AND3_X1   g604(.A1(new_n733), .A2(new_n790), .A3(new_n786), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n790), .B1(new_n733), .B2(new_n786), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n707), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT114), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  OAI211_X1 g609(.A(KEYINPUT114), .B(new_n707), .C1(new_n791), .C2(new_n792), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n789), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n645), .A2(new_n647), .A3(new_n578), .A4(new_n668), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n798), .A2(KEYINPUT112), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n798), .A2(KEYINPUT112), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n773), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT50), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n773), .B(KEYINPUT50), .C1(new_n799), .C2(new_n800), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n780), .A2(new_n785), .A3(new_n797), .A4(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(KEYINPUT109), .B(KEYINPUT51), .ZN(new_n807));
  AOI221_X4 g621(.A(new_n789), .B1(new_n803), .B2(new_n804), .C1(new_n795), .C2(new_n796), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT51), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n809), .B1(new_n771), .B2(new_n778), .ZN(new_n810));
  AOI22_X1  g624(.A1(new_n806), .A2(new_n807), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n340), .B1(new_n791), .B2(new_n792), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(KEYINPUT48), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n773), .A2(new_n683), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n477), .B(KEYINPUT115), .ZN(new_n815));
  OAI211_X1 g629(.A(new_n814), .B(new_n815), .C1(new_n589), .C2(new_n788), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT116), .ZN(new_n817));
  OR2_X1    g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n816), .A2(new_n817), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n811), .A2(new_n813), .A3(new_n818), .A4(new_n819), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n570), .B(KEYINPUT106), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n589), .B1(new_n541), .B2(new_n821), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n822), .A2(new_n579), .A3(new_n487), .A4(new_n601), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n704), .A2(new_n823), .A3(new_n580), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n340), .B(new_n671), .C1(new_n595), .C2(new_n607), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n825), .A2(new_n684), .A3(new_n617), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n725), .B1(new_n719), .B2(new_n721), .ZN(new_n827));
  OAI211_X1 g641(.A(new_n620), .B(new_n821), .C1(new_n715), .C2(new_n716), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n706), .A2(new_n697), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n830), .A2(new_n637), .A3(new_n623), .A4(new_n714), .ZN(new_n831));
  AND4_X1   g645(.A1(new_n824), .A2(new_n826), .A3(new_n827), .A4(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT52), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n709), .A2(new_n642), .A3(new_n664), .ZN(new_n834));
  INV_X1    g648(.A(new_n639), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n835), .B1(new_n701), .B2(new_n703), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT107), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n473), .A2(new_n837), .A3(new_n615), .A4(new_n623), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n615), .A2(new_n472), .A3(new_n469), .A4(new_n623), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(KEYINPUT107), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n838), .A2(new_n655), .A3(new_n840), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n836), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n833), .B1(new_n834), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n541), .A2(new_n570), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(KEYINPUT98), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n541), .A2(new_n700), .A3(new_n570), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n838), .A2(new_n655), .A3(new_n840), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n847), .A2(new_n848), .A3(new_n835), .ZN(new_n849));
  OAI211_X1 g663(.A(new_n678), .B(new_n641), .C1(new_n628), .C2(new_n663), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n849), .A2(KEYINPUT52), .A3(new_n850), .A4(new_n709), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n843), .A2(new_n851), .ZN(new_n852));
  AOI21_X1  g666(.A(KEYINPUT53), .B1(new_n832), .B2(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n825), .A2(new_n684), .A3(new_n617), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n704), .A2(new_n823), .A3(new_n580), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(new_n725), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n722), .A2(new_n831), .A3(new_n857), .ZN(new_n858));
  AND4_X1   g672(.A1(KEYINPUT53), .A2(new_n852), .A3(new_n856), .A4(new_n858), .ZN(new_n859));
  OAI21_X1  g673(.A(KEYINPUT54), .B1(new_n853), .B2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n852), .A2(new_n858), .A3(new_n856), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT53), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT54), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n852), .A2(new_n858), .A3(KEYINPUT53), .A4(new_n856), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n860), .A2(KEYINPUT108), .A3(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT108), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n864), .B1(new_n863), .B2(new_n865), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n868), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n820), .B1(new_n867), .B2(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(G952), .A2(G953), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n768), .B1(new_n872), .B2(new_n873), .ZN(G75));
  AOI21_X1  g688(.A(new_n219), .B1(new_n863), .B2(new_n865), .ZN(new_n875));
  INV_X1    g689(.A(new_n424), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT56), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n421), .A2(new_n422), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n879), .A2(new_n591), .ZN(new_n880));
  XOR2_X1   g694(.A(new_n880), .B(KEYINPUT55), .Z(new_n881));
  XOR2_X1   g695(.A(new_n881), .B(KEYINPUT117), .Z(new_n882));
  NAND3_X1  g696(.A1(new_n877), .A2(new_n878), .A3(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT118), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n877), .A2(KEYINPUT118), .A3(new_n878), .A4(new_n882), .ZN(new_n886));
  INV_X1    g700(.A(new_n875), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n878), .B1(new_n887), .B2(new_n573), .ZN(new_n888));
  AOI22_X1  g702(.A1(new_n885), .A2(new_n886), .B1(new_n881), .B2(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n302), .A2(G952), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(KEYINPUT119), .ZN(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n889), .A2(new_n892), .ZN(G51));
  NAND3_X1  g707(.A1(new_n860), .A2(KEYINPUT120), .A3(new_n866), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT120), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n870), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n465), .A2(KEYINPUT57), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n894), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n465), .A2(KEYINPUT57), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n461), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n875), .A2(new_n743), .A3(new_n741), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n890), .B1(new_n900), .B2(new_n901), .ZN(G54));
  NAND3_X1  g716(.A1(new_n875), .A2(KEYINPUT58), .A3(G475), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n903), .A2(new_n522), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n903), .A2(new_n522), .ZN(new_n905));
  NOR3_X1   g719(.A1(new_n904), .A2(new_n905), .A3(new_n890), .ZN(G60));
  XOR2_X1   g720(.A(new_n586), .B(KEYINPUT59), .Z(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n871), .A2(new_n867), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(new_n583), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(KEYINPUT122), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT122), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n909), .A2(new_n912), .A3(new_n583), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n583), .A2(new_n907), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n894), .A2(new_n896), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(new_n892), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT121), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n915), .A2(KEYINPUT121), .A3(new_n892), .ZN(new_n919));
  AOI22_X1  g733(.A1(new_n911), .A2(new_n913), .B1(new_n918), .B2(new_n919), .ZN(G63));
  NAND2_X1  g734(.A1(new_n863), .A2(new_n865), .ZN(new_n921));
  NAND2_X1  g735(.A1(G217), .A2(G902), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT123), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT60), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n921), .A2(new_n613), .A3(new_n924), .ZN(new_n925));
  AND2_X1   g739(.A1(new_n921), .A2(new_n924), .ZN(new_n926));
  OAI211_X1 g740(.A(new_n892), .B(new_n925), .C1(new_n926), .C2(new_n231), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT61), .Z(G66));
  INV_X1    g742(.A(new_n856), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(new_n302), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT124), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n302), .B1(new_n481), .B2(G224), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(G898), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n421), .B1(new_n934), .B2(G953), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n933), .B(new_n935), .ZN(G69));
  NOR2_X1   g750(.A1(new_n661), .A2(new_n834), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(KEYINPUT62), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n822), .A2(new_n340), .A3(new_n656), .A4(new_n714), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n938), .A2(new_n749), .A3(new_n759), .A4(new_n939), .ZN(new_n940));
  AND2_X1   g754(.A1(new_n940), .A2(new_n302), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n284), .A2(new_n297), .ZN(new_n942));
  XOR2_X1   g756(.A(KEYINPUT125), .B(KEYINPUT126), .Z(new_n943));
  XOR2_X1   g757(.A(new_n942), .B(new_n943), .Z(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(new_n504), .Z(new_n945));
  OR2_X1    g759(.A1(new_n941), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(G900), .A2(G953), .ZN(new_n947));
  INV_X1    g761(.A(new_n340), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n836), .A2(new_n948), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n748), .B1(new_n738), .B2(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(new_n834), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n950), .A2(new_n759), .A3(new_n827), .A4(new_n951), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n945), .B(new_n947), .C1(new_n952), .C2(G953), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n946), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n302), .B1(G227), .B2(G900), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT127), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n955), .B1(new_n953), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n954), .A2(new_n957), .ZN(new_n958));
  OAI211_X1 g772(.A(new_n946), .B(new_n953), .C1(new_n956), .C2(new_n955), .ZN(new_n959));
  AND2_X1   g773(.A1(new_n958), .A2(new_n959), .ZN(G72));
  NAND2_X1  g774(.A1(G472), .A2(G902), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n961), .B(KEYINPUT63), .Z(new_n962));
  OAI21_X1  g776(.A(new_n962), .B1(new_n940), .B2(new_n929), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n890), .B1(new_n963), .B2(new_n650), .ZN(new_n964));
  INV_X1    g778(.A(new_n309), .ZN(new_n965));
  OAI211_X1 g779(.A(new_n921), .B(new_n962), .C1(new_n337), .C2(new_n965), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n962), .B1(new_n952), .B2(new_n929), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n967), .A2(new_n649), .A3(new_n307), .ZN(new_n968));
  AND3_X1   g782(.A1(new_n964), .A2(new_n966), .A3(new_n968), .ZN(G57));
endmodule


