//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 1 0 1 1 0 0 0 1 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 0 0 1 0 0 1 1 1 0 0 0 0 1 0 1 0 1 0 0 0 0 0 0 1 1 0 0 0 0 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:45 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n773,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003;
  INV_X1    g000(.A(G128), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G119), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT75), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT23), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT23), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n188), .A2(new_n189), .A3(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G119), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G128), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n191), .A2(new_n193), .A3(new_n195), .ZN(new_n196));
  AND2_X1   g010(.A1(new_n188), .A2(new_n195), .ZN(new_n197));
  XNOR2_X1  g011(.A(KEYINPUT24), .B(G110), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  OAI22_X1  g013(.A1(new_n196), .A2(G110), .B1(new_n197), .B2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT80), .ZN(new_n201));
  OR2_X1    g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G140), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G125), .ZN(new_n204));
  INV_X1    g018(.A(G125), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G140), .ZN(new_n206));
  INV_X1    g020(.A(G146), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n204), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n200), .A2(new_n201), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT79), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n210), .B1(new_n204), .B2(KEYINPUT16), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n203), .A2(KEYINPUT78), .A3(G125), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT78), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n213), .B1(new_n205), .B2(G140), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n205), .A2(G140), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n212), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT16), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n211), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n206), .A2(KEYINPUT78), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(new_n204), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n220), .A2(new_n210), .A3(KEYINPUT16), .A4(new_n212), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n218), .A2(G146), .A3(new_n221), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n202), .A2(new_n208), .A3(new_n209), .A4(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G110), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT76), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n224), .B1(new_n196), .B2(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n226), .B1(new_n225), .B2(new_n196), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT77), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI211_X1 g043(.A(new_n226), .B(KEYINPUT77), .C1(new_n225), .C2(new_n196), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n218), .A2(new_n221), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(new_n207), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(new_n222), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n199), .A2(new_n197), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n223), .B1(new_n231), .B2(new_n236), .ZN(new_n237));
  XNOR2_X1  g051(.A(KEYINPUT22), .B(G137), .ZN(new_n238));
  INV_X1    g052(.A(G953), .ZN(new_n239));
  AND3_X1   g053(.A1(new_n239), .A2(G221), .A3(G234), .ZN(new_n240));
  XOR2_X1   g054(.A(new_n238), .B(new_n240), .Z(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  OR2_X1    g056(.A1(new_n237), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(G902), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n237), .A2(new_n242), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n243), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT81), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n247), .A2(KEYINPUT25), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n246), .A2(new_n249), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n243), .A2(new_n244), .A3(new_n245), .A4(new_n248), .ZN(new_n251));
  INV_X1    g065(.A(G217), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n252), .B1(G234), .B2(new_n244), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n250), .A2(new_n251), .A3(new_n253), .ZN(new_n254));
  AND2_X1   g068(.A1(new_n243), .A2(new_n245), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n253), .A2(G902), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n207), .A2(G143), .ZN(new_n260));
  INV_X1    g074(.A(G143), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G146), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  OAI211_X1 g077(.A(KEYINPUT84), .B(KEYINPUT1), .C1(new_n261), .C2(G146), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G128), .ZN(new_n265));
  AOI21_X1  g079(.A(KEYINPUT84), .B1(new_n260), .B2(KEYINPUT1), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n263), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(KEYINPUT85), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n187), .A2(KEYINPUT1), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n269), .A2(new_n260), .A3(new_n262), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(KEYINPUT67), .ZN(new_n271));
  XNOR2_X1  g085(.A(G143), .B(G146), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT67), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n272), .A2(new_n273), .A3(new_n269), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n271), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT85), .ZN(new_n276));
  OAI211_X1 g090(.A(new_n276), .B(new_n263), .C1(new_n265), .C2(new_n266), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n268), .A2(new_n275), .A3(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(G101), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT3), .ZN(new_n280));
  INV_X1    g094(.A(G107), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n280), .A2(new_n281), .A3(G104), .ZN(new_n282));
  INV_X1    g096(.A(G104), .ZN(new_n283));
  AOI21_X1  g097(.A(KEYINPUT3), .B1(new_n283), .B2(G107), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n283), .A2(G107), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n279), .B(new_n282), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n281), .A2(G104), .ZN(new_n287));
  OAI21_X1  g101(.A(G101), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  AND2_X1   g102(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(KEYINPUT10), .B1(new_n278), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT64), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n291), .B1(new_n207), .B2(G143), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n261), .A2(KEYINPUT64), .A3(G146), .ZN(new_n293));
  AOI22_X1  g107(.A1(new_n292), .A2(new_n293), .B1(G143), .B2(new_n207), .ZN(new_n294));
  XNOR2_X1  g108(.A(KEYINPUT0), .B(G128), .ZN(new_n295));
  NAND2_X1  g109(.A1(KEYINPUT0), .A2(G128), .ZN(new_n296));
  OAI22_X1  g110(.A1(new_n294), .A2(new_n295), .B1(new_n263), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n282), .B1(new_n284), .B2(new_n285), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT4), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n299), .A2(new_n300), .A3(G101), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n299), .A2(G101), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n302), .A2(KEYINPUT4), .A3(new_n286), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n298), .A2(new_n301), .A3(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n273), .B1(new_n272), .B2(new_n269), .ZN(new_n305));
  AND4_X1   g119(.A1(new_n273), .A2(new_n269), .A3(new_n260), .A4(new_n262), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n187), .B1(new_n260), .B2(KEYINPUT1), .ZN(new_n307));
  OAI22_X1  g121(.A1(new_n305), .A2(new_n306), .B1(new_n294), .B2(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n308), .A2(KEYINPUT10), .A3(new_n289), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n304), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT11), .ZN(new_n311));
  INV_X1    g125(.A(G134), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n311), .B1(new_n312), .B2(G137), .ZN(new_n313));
  INV_X1    g127(.A(G137), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n314), .A2(KEYINPUT11), .A3(G134), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n312), .A2(G137), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n313), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G131), .ZN(new_n318));
  INV_X1    g132(.A(G131), .ZN(new_n319));
  NAND4_X1  g133(.A1(new_n313), .A2(new_n315), .A3(new_n319), .A4(new_n316), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  NOR3_X1   g135(.A1(new_n290), .A2(new_n310), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n239), .A2(G227), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n323), .B(KEYINPUT82), .ZN(new_n324));
  XNOR2_X1  g138(.A(G110), .B(G140), .ZN(new_n325));
  XNOR2_X1  g139(.A(new_n324), .B(new_n325), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n322), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT86), .ZN(new_n328));
  AOI21_X1  g142(.A(KEYINPUT12), .B1(new_n321), .B2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n278), .A2(new_n289), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n308), .A2(new_n289), .ZN(new_n333));
  OAI211_X1 g147(.A(new_n321), .B(new_n330), .C1(new_n332), .C2(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n333), .B1(new_n289), .B2(new_n278), .ZN(new_n335));
  INV_X1    g149(.A(new_n321), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n329), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n334), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n327), .A2(new_n338), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n321), .B1(new_n290), .B2(new_n310), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n326), .B1(new_n341), .B2(new_n322), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  XNOR2_X1  g157(.A(KEYINPUT88), .B(G469), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n343), .A2(new_n244), .A3(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT89), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(G902), .B1(new_n339), .B2(new_n342), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n348), .A2(KEYINPUT89), .A3(new_n344), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT87), .ZN(new_n350));
  XOR2_X1   g164(.A(new_n326), .B(KEYINPUT83), .Z(new_n351));
  INV_X1    g165(.A(new_n322), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n351), .B1(new_n338), .B2(new_n352), .ZN(new_n353));
  NOR3_X1   g167(.A1(new_n341), .A2(new_n322), .A3(new_n326), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n350), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n327), .A2(new_n340), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n322), .B1(new_n334), .B2(new_n337), .ZN(new_n357));
  OAI211_X1 g171(.A(new_n356), .B(KEYINPUT87), .C1(new_n357), .C2(new_n351), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n355), .A2(new_n244), .A3(new_n358), .ZN(new_n359));
  AOI22_X1  g173(.A1(new_n347), .A2(new_n349), .B1(new_n359), .B2(G469), .ZN(new_n360));
  XOR2_X1   g174(.A(KEYINPUT9), .B(G234), .Z(new_n361));
  NAND3_X1  g175(.A1(new_n361), .A2(G217), .A3(new_n239), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  XNOR2_X1  g177(.A(G128), .B(G143), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(new_n312), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n261), .A2(KEYINPUT13), .A3(G128), .ZN(new_n366));
  AOI21_X1  g180(.A(KEYINPUT13), .B1(new_n261), .B2(G128), .ZN(new_n367));
  OAI221_X1 g181(.A(new_n366), .B1(G128), .B2(new_n261), .C1(new_n367), .C2(KEYINPUT97), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(KEYINPUT97), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(G134), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(G122), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT68), .ZN(new_n373));
  INV_X1    g187(.A(G116), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(KEYINPUT68), .A2(G116), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n372), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n374), .A2(G122), .ZN(new_n378));
  NOR3_X1   g192(.A1(new_n377), .A2(KEYINPUT96), .A3(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT96), .ZN(new_n380));
  INV_X1    g194(.A(new_n376), .ZN(new_n381));
  NOR2_X1   g195(.A1(KEYINPUT68), .A2(G116), .ZN(new_n382));
  OAI21_X1  g196(.A(G122), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n378), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n380), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NOR3_X1   g199(.A1(new_n379), .A2(new_n385), .A3(new_n281), .ZN(new_n386));
  OAI21_X1  g200(.A(KEYINPUT96), .B1(new_n377), .B2(new_n378), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n383), .A2(new_n380), .A3(new_n384), .ZN(new_n388));
  AOI21_X1  g202(.A(G107), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n365), .B(new_n371), .C1(new_n386), .C2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n389), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT14), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n377), .A2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n384), .B1(new_n377), .B2(new_n392), .ZN(new_n395));
  OAI21_X1  g209(.A(G107), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n364), .B(new_n312), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n391), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n363), .B1(new_n390), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n390), .A2(new_n398), .A3(new_n363), .ZN(new_n401));
  AOI21_X1  g215(.A(G902), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(G478), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n402), .B(KEYINPUT98), .C1(KEYINPUT15), .C2(new_n403), .ZN(new_n404));
  AND2_X1   g218(.A1(new_n239), .A2(G952), .ZN(new_n405));
  NAND2_X1  g219(.A1(G234), .A2(G237), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n407), .B(KEYINPUT99), .ZN(new_n408));
  AND3_X1   g222(.A1(new_n406), .A2(G902), .A3(G953), .ZN(new_n409));
  XNOR2_X1  g223(.A(KEYINPUT21), .B(G898), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  AND2_X1   g225(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n403), .A2(KEYINPUT15), .ZN(new_n414));
  INV_X1    g228(.A(new_n401), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n244), .B1(new_n415), .B2(new_n399), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT98), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n414), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n416), .A2(new_n417), .ZN(new_n419));
  OAI211_X1 g233(.A(new_n404), .B(new_n413), .C1(new_n418), .C2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  XNOR2_X1  g235(.A(KEYINPUT2), .B(G113), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n194), .B1(new_n375), .B2(new_n376), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n374), .A2(G119), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n422), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n422), .ZN(new_n426));
  OAI21_X1  g240(.A(G119), .B1(new_n381), .B2(new_n382), .ZN(new_n427));
  INV_X1    g241(.A(new_n424), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n425), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n303), .A2(new_n430), .A3(new_n301), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n427), .A2(KEYINPUT5), .A3(new_n428), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT5), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n424), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n432), .A2(G113), .A3(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n435), .A2(new_n429), .A3(new_n289), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n431), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(KEYINPUT90), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT90), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n431), .A2(new_n436), .A3(new_n439), .ZN(new_n440));
  XOR2_X1   g254(.A(G110), .B(G122), .Z(new_n441));
  NAND3_X1  g255(.A1(new_n438), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT6), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND4_X1  g258(.A1(new_n438), .A2(KEYINPUT6), .A3(new_n440), .A4(new_n441), .ZN(new_n445));
  INV_X1    g259(.A(new_n441), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n431), .A2(new_n436), .A3(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n444), .A2(new_n445), .A3(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(KEYINPUT91), .B1(new_n298), .B2(new_n205), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n292), .A2(new_n293), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(new_n260), .ZN(new_n451));
  INV_X1    g265(.A(new_n307), .ZN(new_n452));
  AOI22_X1  g266(.A1(new_n451), .A2(new_n452), .B1(new_n271), .B2(new_n274), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(new_n205), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT91), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n297), .A2(new_n455), .A3(G125), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n449), .A2(new_n454), .A3(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(G224), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n458), .A2(G953), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n459), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n449), .A2(new_n454), .A3(new_n461), .A4(new_n456), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n448), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(G210), .B1(G237), .B2(G902), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n454), .B1(new_n205), .B2(new_n298), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n461), .A2(KEYINPUT7), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g282(.A(KEYINPUT92), .B(KEYINPUT8), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n441), .B(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n436), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n289), .B1(new_n435), .B2(new_n429), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n468), .A2(new_n473), .A3(new_n447), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT7), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n462), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n244), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n464), .A2(new_n465), .A3(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n465), .ZN(new_n480));
  INV_X1    g294(.A(new_n463), .ZN(new_n481));
  INV_X1    g295(.A(new_n447), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n482), .B1(new_n442), .B2(new_n443), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n481), .B1(new_n483), .B2(new_n445), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n480), .B1(new_n484), .B2(new_n477), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n479), .A2(new_n485), .ZN(new_n486));
  OAI21_X1  g300(.A(G214), .B1(G237), .B2(G902), .ZN(new_n487));
  INV_X1    g301(.A(G475), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT72), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n489), .A2(G237), .ZN(new_n490));
  INV_X1    g304(.A(G237), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n491), .A2(KEYINPUT72), .ZN(new_n492));
  OAI211_X1 g306(.A(G214), .B(new_n239), .C1(new_n490), .C2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(new_n261), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n491), .A2(KEYINPUT72), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n489), .A2(G237), .ZN(new_n496));
  AOI21_X1  g310(.A(G953), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n497), .A2(G143), .A3(G214), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n319), .B1(new_n494), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(KEYINPUT18), .ZN(new_n500));
  NAND2_X1  g314(.A1(KEYINPUT18), .A2(G131), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n494), .A2(new_n498), .A3(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n216), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n208), .B1(new_n503), .B2(new_n207), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n500), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n493), .A2(new_n261), .ZN(new_n506));
  AOI21_X1  g320(.A(G143), .B1(new_n497), .B2(G214), .ZN(new_n507));
  OAI211_X1 g321(.A(KEYINPUT17), .B(G131), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n233), .A2(new_n222), .A3(new_n508), .ZN(new_n509));
  NOR3_X1   g323(.A1(new_n506), .A2(new_n507), .A3(G131), .ZN(new_n510));
  NOR3_X1   g324(.A1(new_n510), .A2(new_n499), .A3(KEYINPUT17), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n505), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  XNOR2_X1  g326(.A(G113), .B(G122), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n513), .B(new_n283), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n514), .B(new_n505), .C1(new_n509), .C2(new_n511), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n488), .B1(new_n518), .B2(new_n244), .ZN(new_n519));
  NOR2_X1   g333(.A1(G475), .A2(G902), .ZN(new_n520));
  OAI21_X1  g334(.A(KEYINPUT93), .B1(new_n510), .B2(new_n499), .ZN(new_n521));
  OAI21_X1  g335(.A(G131), .B1(new_n506), .B2(new_n507), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT93), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n494), .A2(new_n319), .A3(new_n498), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  OR2_X1    g339(.A1(KEYINPUT94), .A2(KEYINPUT19), .ZN(new_n526));
  NAND2_X1  g340(.A1(KEYINPUT94), .A2(KEYINPUT19), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n526), .A2(new_n204), .A3(new_n206), .A4(new_n527), .ZN(new_n528));
  OR2_X1    g342(.A1(new_n528), .A2(KEYINPUT95), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n216), .A2(KEYINPUT19), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n528), .A2(KEYINPUT95), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n529), .A2(new_n530), .A3(new_n207), .A4(new_n531), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n521), .A2(new_n222), .A3(new_n525), .A4(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n514), .B1(new_n533), .B2(new_n505), .ZN(new_n534));
  INV_X1    g348(.A(new_n517), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n520), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(KEYINPUT20), .ZN(new_n537));
  AND3_X1   g351(.A1(new_n500), .A2(new_n502), .A3(new_n504), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n523), .B1(new_n522), .B2(new_n524), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n222), .A2(new_n532), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n538), .B1(new_n541), .B2(new_n525), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n517), .B1(new_n542), .B2(new_n514), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT20), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n543), .A2(new_n544), .A3(new_n520), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n519), .B1(new_n537), .B2(new_n545), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n421), .A2(new_n486), .A3(new_n487), .A4(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(G221), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n548), .B1(new_n361), .B2(new_n244), .ZN(new_n549));
  NOR3_X1   g363(.A1(new_n360), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT74), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT28), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n298), .A2(new_n321), .ZN(new_n553));
  INV_X1    g367(.A(new_n430), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n312), .A2(G137), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n314), .A2(G134), .ZN(new_n557));
  OAI21_X1  g371(.A(G131), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n320), .A2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT69), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n320), .A2(new_n558), .A3(KEYINPUT69), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n451), .A2(new_n452), .ZN(new_n563));
  AOI22_X1  g377(.A1(new_n561), .A2(new_n562), .B1(new_n563), .B2(new_n275), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n552), .B1(new_n555), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n497), .A2(G210), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n566), .B(G101), .ZN(new_n567));
  XNOR2_X1  g381(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n567), .B(new_n568), .ZN(new_n569));
  AND2_X1   g383(.A1(new_n569), .A2(KEYINPUT29), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT70), .ZN(new_n571));
  AOI22_X1  g385(.A1(new_n564), .A2(new_n571), .B1(new_n321), .B2(new_n298), .ZN(new_n572));
  AND3_X1   g386(.A1(new_n320), .A2(new_n558), .A3(KEYINPUT69), .ZN(new_n573));
  AOI21_X1  g387(.A(KEYINPUT69), .B1(new_n320), .B2(new_n558), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  OAI21_X1  g389(.A(KEYINPUT70), .B1(new_n575), .B2(new_n453), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n554), .B1(new_n572), .B2(new_n576), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n308), .B(new_n571), .C1(new_n574), .C2(new_n573), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n576), .A2(new_n554), .A3(new_n578), .A4(new_n553), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(KEYINPUT71), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT71), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n572), .A2(new_n581), .A3(new_n554), .A4(new_n576), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n577), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n565), .B(new_n570), .C1(new_n583), .C2(new_n552), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n244), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n297), .A2(KEYINPUT65), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT65), .ZN(new_n587));
  OAI221_X1 g401(.A(new_n587), .B1(new_n263), .B2(new_n296), .C1(new_n294), .C2(new_n295), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n586), .A2(new_n321), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(KEYINPUT66), .ZN(new_n590));
  AOI22_X1  g404(.A1(new_n297), .A2(KEYINPUT65), .B1(new_n318), .B2(new_n320), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT66), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n591), .A2(new_n592), .A3(new_n588), .ZN(new_n593));
  OAI211_X1 g407(.A(new_n590), .B(new_n593), .C1(new_n453), .C2(new_n559), .ZN(new_n594));
  AOI22_X1  g408(.A1(new_n580), .A2(new_n582), .B1(new_n594), .B2(new_n430), .ZN(new_n595));
  OAI211_X1 g409(.A(new_n565), .B(new_n569), .C1(new_n595), .C2(new_n552), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT30), .ZN(new_n597));
  OAI22_X1  g411(.A1(new_n589), .A2(KEYINPUT66), .B1(new_n453), .B2(new_n559), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n592), .B1(new_n591), .B2(new_n588), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n597), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n572), .A2(KEYINPUT30), .A3(new_n576), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n600), .A2(new_n430), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n580), .A2(new_n582), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n569), .ZN(new_n605));
  AOI21_X1  g419(.A(KEYINPUT29), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n585), .B1(new_n596), .B2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(G472), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n551), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  AND2_X1   g423(.A1(new_n606), .A2(new_n596), .ZN(new_n610));
  OAI211_X1 g424(.A(KEYINPUT74), .B(G472), .C1(new_n610), .C2(new_n585), .ZN(new_n611));
  AND2_X1   g425(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n605), .B1(new_n580), .B2(new_n582), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n602), .B1(new_n613), .B2(KEYINPUT73), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT73), .ZN(new_n615));
  AOI211_X1 g429(.A(new_n615), .B(new_n605), .C1(new_n580), .C2(new_n582), .ZN(new_n616));
  OAI21_X1  g430(.A(KEYINPUT31), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n603), .A2(new_n569), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n615), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT31), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n613), .A2(KEYINPUT73), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n619), .A2(new_n620), .A3(new_n621), .A4(new_n602), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n565), .B1(new_n595), .B2(new_n552), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n605), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n617), .A2(new_n622), .A3(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(G472), .A2(G902), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT32), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n625), .A2(KEYINPUT32), .A3(new_n626), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  OAI211_X1 g445(.A(new_n259), .B(new_n550), .C1(new_n612), .C2(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(G101), .ZN(G3));
  NOR3_X1   g447(.A1(new_n360), .A2(new_n258), .A3(new_n549), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n464), .A2(KEYINPUT100), .A3(new_n465), .A4(new_n478), .ZN(new_n635));
  AND2_X1   g449(.A1(new_n635), .A2(new_n487), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT100), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n479), .A2(new_n485), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n537), .A2(new_n545), .ZN(new_n640));
  INV_X1    g454(.A(new_n519), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT33), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n643), .B1(new_n415), .B2(new_n399), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n400), .A2(KEYINPUT33), .A3(new_n401), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n644), .A2(new_n645), .A3(G478), .A4(new_n244), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n416), .A2(new_n403), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n642), .A2(new_n648), .ZN(new_n649));
  NOR3_X1   g463(.A1(new_n639), .A2(new_n412), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n625), .A2(new_n244), .ZN(new_n651));
  AOI22_X1  g465(.A1(new_n651), .A2(G472), .B1(new_n625), .B2(new_n626), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n634), .A2(new_n650), .A3(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT34), .B(G104), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G6));
  AOI21_X1  g469(.A(new_n544), .B1(new_n543), .B2(new_n520), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n519), .B1(new_n656), .B2(KEYINPUT101), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n404), .B1(new_n418), .B2(new_n419), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT101), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n537), .A2(new_n659), .A3(new_n545), .ZN(new_n660));
  AND3_X1   g474(.A1(new_n657), .A2(new_n658), .A3(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n662), .A2(new_n639), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n634), .A2(new_n652), .A3(new_n413), .A4(new_n663), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT35), .B(G107), .Z(new_n665));
  XNOR2_X1  g479(.A(KEYINPUT102), .B(KEYINPUT103), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n664), .B(new_n667), .ZN(G9));
  XNOR2_X1  g482(.A(new_n237), .B(KEYINPUT104), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n242), .A2(KEYINPUT36), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n669), .B1(KEYINPUT36), .B2(new_n242), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n672), .A2(new_n673), .A3(new_n256), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n254), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n550), .A2(new_n652), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(KEYINPUT37), .B(G110), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(KEYINPUT105), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n676), .B(new_n678), .ZN(G12));
  INV_X1    g493(.A(G900), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n409), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(KEYINPUT106), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n408), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n661), .A2(new_n638), .A3(new_n636), .A4(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT107), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AND3_X1   g500(.A1(new_n638), .A2(new_n487), .A3(new_n635), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n687), .A2(KEYINPUT107), .A3(new_n661), .A4(new_n683), .ZN(new_n688));
  AND2_X1   g502(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(new_n675), .ZN(new_n690));
  AND3_X1   g504(.A1(new_n625), .A2(KEYINPUT32), .A3(new_n626), .ZN(new_n691));
  AOI21_X1  g505(.A(KEYINPUT32), .B1(new_n625), .B2(new_n626), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n609), .A2(new_n611), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n690), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(new_n549), .ZN(new_n696));
  AND2_X1   g510(.A1(new_n359), .A2(G469), .ZN(new_n697));
  AND4_X1   g511(.A1(KEYINPUT89), .A2(new_n343), .A3(new_n244), .A4(new_n344), .ZN(new_n698));
  AOI21_X1  g512(.A(KEYINPUT89), .B1(new_n348), .B2(new_n344), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n696), .B1(new_n697), .B2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n689), .A2(new_n695), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G128), .ZN(G30));
  XOR2_X1   g518(.A(new_n683), .B(KEYINPUT39), .Z(new_n705));
  NOR2_X1   g519(.A1(new_n701), .A2(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  OR2_X1    g521(.A1(new_n707), .A2(KEYINPUT40), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n614), .A2(new_n616), .ZN(new_n709));
  INV_X1    g523(.A(new_n583), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n709), .B1(new_n605), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g525(.A(G472), .B1(new_n711), .B2(G902), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n693), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n707), .A2(KEYINPUT40), .ZN(new_n714));
  AND2_X1   g528(.A1(new_n479), .A2(new_n485), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(KEYINPUT38), .ZN(new_n716));
  INV_X1    g530(.A(new_n487), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n642), .A2(new_n658), .ZN(new_n718));
  NOR4_X1   g532(.A1(new_n716), .A2(new_n717), .A3(new_n675), .A4(new_n718), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n708), .A2(new_n713), .A3(new_n714), .A4(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G143), .ZN(G45));
  AOI22_X1  g535(.A1(new_n640), .A2(new_n641), .B1(new_n647), .B2(new_n646), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n636), .A2(new_n722), .A3(new_n638), .A4(new_n683), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT108), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n723), .B(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n694), .A2(new_n629), .A3(new_n630), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n725), .A2(new_n726), .A3(new_n702), .A4(new_n675), .ZN(new_n727));
  XOR2_X1   g541(.A(KEYINPUT109), .B(G146), .Z(new_n728));
  XNOR2_X1  g542(.A(new_n727), .B(new_n728), .ZN(G48));
  INV_X1    g543(.A(G469), .ZN(new_n730));
  OR2_X1    g544(.A1(new_n348), .A2(new_n730), .ZN(new_n731));
  OAI211_X1 g545(.A(new_n696), .B(new_n731), .C1(new_n698), .C2(new_n699), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(KEYINPUT110), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n726), .A2(new_n733), .A3(new_n259), .A4(new_n650), .ZN(new_n734));
  XNOR2_X1  g548(.A(KEYINPUT41), .B(G113), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n734), .B(new_n735), .ZN(G15));
  NOR3_X1   g550(.A1(new_n662), .A2(new_n639), .A3(new_n412), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n726), .A2(new_n733), .A3(new_n259), .A4(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G116), .ZN(G18));
  NAND2_X1  g553(.A1(new_n421), .A2(new_n546), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n639), .A2(new_n732), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n726), .A2(new_n741), .A3(new_n675), .A4(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G119), .ZN(G21));
  INV_X1    g558(.A(new_n565), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n745), .B1(new_n710), .B2(KEYINPUT28), .ZN(new_n746));
  OAI211_X1 g560(.A(new_n617), .B(new_n622), .C1(new_n569), .C2(new_n746), .ZN(new_n747));
  AOI22_X1  g561(.A1(new_n651), .A2(G472), .B1(new_n626), .B2(new_n747), .ZN(new_n748));
  NOR3_X1   g562(.A1(new_n639), .A2(new_n412), .A3(new_n718), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n733), .A2(new_n259), .A3(new_n748), .A4(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G122), .ZN(G24));
  INV_X1    g565(.A(new_n683), .ZN(new_n752));
  OAI21_X1  g566(.A(KEYINPUT111), .B1(new_n649), .B2(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT111), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n722), .A2(new_n754), .A3(new_n683), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  AND4_X1   g570(.A1(new_n675), .A2(new_n756), .A3(new_n748), .A4(new_n742), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(new_n205), .ZN(G27));
  NAND2_X1  g572(.A1(new_n347), .A2(new_n349), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n353), .A2(new_n354), .ZN(new_n760));
  OAI21_X1  g574(.A(G469), .B1(new_n760), .B2(G902), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n549), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n486), .A2(new_n717), .ZN(new_n763));
  AND2_X1   g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n726), .A2(new_n259), .A3(new_n756), .A4(new_n764), .ZN(new_n765));
  NOR2_X1   g579(.A1(KEYINPUT112), .A2(KEYINPUT42), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n258), .B1(new_n693), .B2(new_n694), .ZN(new_n768));
  INV_X1    g582(.A(new_n766), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n768), .A2(new_n756), .A3(new_n764), .A4(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n767), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G131), .ZN(G33));
  NOR2_X1   g586(.A1(new_n662), .A2(new_n752), .ZN(new_n773));
  AND4_X1   g587(.A1(new_n259), .A2(new_n726), .A3(new_n764), .A4(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(new_n312), .ZN(G36));
  INV_X1    g589(.A(new_n652), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n546), .A2(new_n648), .ZN(new_n777));
  NAND2_X1  g591(.A1(KEYINPUT113), .A2(KEYINPUT43), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g593(.A1(KEYINPUT113), .A2(KEYINPUT43), .ZN(new_n780));
  MUX2_X1   g594(.A(new_n779), .B(new_n777), .S(new_n780), .Z(new_n781));
  NAND3_X1  g595(.A1(new_n776), .A2(new_n781), .A3(new_n675), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT44), .ZN(new_n783));
  OR2_X1    g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT45), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n355), .A2(new_n785), .A3(new_n358), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n730), .B1(new_n760), .B2(KEYINPUT45), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(G469), .A2(G902), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n790), .A2(KEYINPUT46), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n788), .A2(new_n789), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT46), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n791), .A2(new_n759), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(new_n696), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n796), .A2(new_n705), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n763), .B(KEYINPUT114), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n782), .A2(new_n783), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n784), .A2(new_n797), .A3(new_n799), .A4(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(KEYINPUT115), .B(G137), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n801), .B(new_n802), .ZN(G39));
  NAND2_X1  g617(.A1(new_n796), .A2(KEYINPUT47), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT47), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n795), .A2(new_n805), .A3(new_n696), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(new_n763), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n722), .A2(new_n258), .A3(new_n683), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n726), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n808), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(G140), .ZN(G42));
  INV_X1    g627(.A(new_n408), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n781), .A2(new_n814), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n748), .A2(new_n259), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(new_n716), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n818), .A2(new_n487), .A3(new_n732), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT50), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n820), .B(new_n821), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n809), .A2(new_n732), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n815), .A2(new_n823), .ZN(new_n824));
  AND2_X1   g638(.A1(new_n748), .A2(new_n675), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n823), .A2(new_n259), .A3(new_n814), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n713), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n642), .A2(new_n648), .ZN(new_n828));
  AOI22_X1  g642(.A1(new_n824), .A2(new_n825), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n822), .A2(new_n829), .ZN(new_n830));
  OR2_X1    g644(.A1(new_n808), .A2(KEYINPUT116), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n808), .A2(KEYINPUT116), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n759), .A2(new_n549), .A3(new_n731), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n831), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n817), .A2(new_n799), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n830), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  OR2_X1    g650(.A1(new_n836), .A2(KEYINPUT51), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n824), .A2(new_n768), .ZN(new_n838));
  XNOR2_X1  g652(.A(new_n838), .B(KEYINPUT48), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n817), .A2(new_n742), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n827), .A2(new_n722), .ZN(new_n841));
  AND4_X1   g655(.A1(new_n405), .A2(new_n839), .A3(new_n840), .A4(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n822), .A2(KEYINPUT51), .A3(new_n829), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT117), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n807), .A2(new_n844), .A3(new_n833), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(new_n835), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n844), .B1(new_n807), .B2(new_n833), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  OAI21_X1  g662(.A(KEYINPUT118), .B1(new_n843), .B2(new_n848), .ZN(new_n849));
  OR3_X1    g663(.A1(new_n843), .A2(new_n848), .A3(KEYINPUT118), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n837), .A2(new_n842), .A3(new_n849), .A4(new_n850), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n774), .B1(new_n767), .B2(new_n770), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n657), .A2(new_n660), .ZN(new_n853));
  NOR4_X1   g667(.A1(new_n809), .A2(new_n853), .A3(new_n658), .A4(new_n752), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n726), .A2(new_n702), .A3(new_n854), .A4(new_n675), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n764), .A2(new_n675), .A3(new_n748), .A4(new_n756), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n546), .A2(new_n658), .ZN(new_n858));
  AOI211_X1 g672(.A(new_n717), .B(new_n715), .C1(new_n649), .C2(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n634), .A2(new_n859), .A3(new_n413), .A4(new_n652), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n632), .A2(new_n676), .A3(new_n860), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n857), .A2(new_n861), .ZN(new_n862));
  AND4_X1   g676(.A1(new_n734), .A2(new_n738), .A3(new_n743), .A4(new_n750), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n852), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n825), .A2(new_n742), .A3(new_n756), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n639), .A2(new_n718), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n675), .A2(new_n752), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n713), .A2(new_n866), .A3(new_n762), .A4(new_n867), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n703), .A2(new_n727), .A3(new_n865), .A4(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT52), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  AOI211_X1 g685(.A(new_n701), .B(new_n690), .C1(new_n693), .C2(new_n694), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n757), .B1(new_n872), .B2(new_n689), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n873), .A2(KEYINPUT52), .A3(new_n727), .A4(new_n868), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n864), .A2(new_n875), .A3(KEYINPUT53), .ZN(new_n876));
  AOI21_X1  g690(.A(KEYINPUT53), .B1(new_n864), .B2(new_n875), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n876), .A2(new_n877), .A3(KEYINPUT54), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT54), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT53), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n871), .A2(new_n874), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n852), .A2(new_n862), .A3(new_n863), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n880), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n864), .A2(new_n875), .A3(KEYINPUT53), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n879), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  OR2_X1    g699(.A1(new_n878), .A2(new_n885), .ZN(new_n886));
  OAI22_X1  g700(.A1(new_n851), .A2(new_n886), .B1(G952), .B2(G953), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n759), .A2(new_n731), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(KEYINPUT49), .ZN(new_n889));
  OR4_X1    g703(.A1(new_n258), .A2(new_n777), .A3(new_n549), .A4(new_n717), .ZN(new_n890));
  OR4_X1    g704(.A1(new_n713), .A2(new_n889), .A3(new_n818), .A4(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n887), .A2(new_n891), .ZN(G75));
  NOR2_X1   g706(.A1(new_n239), .A2(G952), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n883), .A2(new_n884), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(G902), .ZN(new_n896));
  INV_X1    g710(.A(new_n896), .ZN(new_n897));
  AOI21_X1  g711(.A(KEYINPUT56), .B1(new_n897), .B2(G210), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n448), .A2(new_n463), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n899), .A2(new_n484), .ZN(new_n900));
  XOR2_X1   g714(.A(KEYINPUT119), .B(KEYINPUT55), .Z(new_n901));
  XNOR2_X1  g715(.A(new_n900), .B(new_n901), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n894), .B1(new_n898), .B2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT56), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n896), .A2(KEYINPUT120), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT120), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n895), .A2(new_n907), .A3(G902), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n905), .B1(new_n909), .B2(new_n480), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n903), .A2(new_n910), .ZN(G51));
  XOR2_X1   g725(.A(new_n789), .B(KEYINPUT57), .Z(new_n912));
  OAI21_X1  g726(.A(new_n912), .B1(new_n878), .B2(new_n885), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT121), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  OAI211_X1 g729(.A(KEYINPUT121), .B(new_n912), .C1(new_n878), .C2(new_n885), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n915), .A2(new_n343), .A3(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n909), .A2(new_n786), .A3(new_n787), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n893), .B1(new_n917), .B2(new_n918), .ZN(G54));
  NAND2_X1  g733(.A1(KEYINPUT58), .A2(G475), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n920), .B1(new_n906), .B2(new_n908), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n894), .B1(new_n921), .B2(new_n543), .ZN(new_n922));
  INV_X1    g736(.A(new_n543), .ZN(new_n923));
  AOI211_X1 g737(.A(new_n923), .B(new_n920), .C1(new_n906), .C2(new_n908), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n922), .A2(new_n924), .ZN(G60));
  NAND2_X1  g739(.A1(G478), .A2(G902), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(KEYINPUT122), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT59), .ZN(new_n928));
  AND4_X1   g742(.A1(new_n644), .A2(new_n886), .A3(new_n645), .A4(new_n928), .ZN(new_n929));
  AOI22_X1  g743(.A1(new_n886), .A2(new_n928), .B1(new_n644), .B2(new_n645), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n929), .A2(new_n893), .A3(new_n930), .ZN(G63));
  NAND2_X1  g745(.A1(new_n672), .A2(new_n673), .ZN(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(G217), .A2(G902), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT60), .ZN(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(KEYINPUT123), .B1(new_n895), .B2(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT123), .ZN(new_n938));
  AOI211_X1 g752(.A(new_n938), .B(new_n935), .C1(new_n883), .C2(new_n884), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n933), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n936), .B1(new_n876), .B2(new_n877), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(new_n938), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n895), .A2(KEYINPUT123), .A3(new_n936), .ZN(new_n943));
  INV_X1    g757(.A(new_n255), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n940), .A2(new_n894), .A3(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT61), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n940), .A2(KEYINPUT61), .A3(new_n945), .A4(new_n894), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n949), .ZN(G66));
  OAI21_X1  g764(.A(G953), .B1(new_n410), .B2(new_n458), .ZN(new_n951));
  INV_X1    g765(.A(new_n861), .ZN(new_n952));
  AND2_X1   g766(.A1(new_n863), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n951), .B1(new_n953), .B2(G953), .ZN(new_n954));
  OAI211_X1 g768(.A(new_n483), .B(new_n445), .C1(G898), .C2(new_n239), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n954), .B(new_n955), .ZN(G69));
  NAND2_X1  g770(.A1(new_n600), .A2(new_n601), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n957), .B(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n873), .A2(new_n727), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n720), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT62), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n961), .A2(KEYINPUT62), .A3(new_n720), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n649), .A2(new_n858), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n768), .A2(new_n706), .A3(new_n763), .A4(new_n967), .ZN(new_n968));
  AND3_X1   g782(.A1(new_n812), .A2(new_n968), .A3(new_n801), .ZN(new_n969));
  AND2_X1   g783(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n960), .B1(new_n970), .B2(G953), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT124), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n961), .A2(new_n801), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(KEYINPUT125), .ZN(new_n975));
  INV_X1    g789(.A(new_n852), .ZN(new_n976));
  OR2_X1    g790(.A1(new_n976), .A2(KEYINPUT126), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n797), .A2(new_n768), .A3(new_n866), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n812), .A2(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n979), .B1(KEYINPUT126), .B2(new_n976), .ZN(new_n980));
  NAND4_X1  g794(.A1(new_n975), .A2(new_n239), .A3(new_n977), .A4(new_n980), .ZN(new_n981));
  OAI211_X1 g795(.A(new_n981), .B(new_n959), .C1(new_n680), .C2(new_n239), .ZN(new_n982));
  OAI211_X1 g796(.A(KEYINPUT124), .B(new_n960), .C1(new_n970), .C2(G953), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n973), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n239), .B1(G227), .B2(G900), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g800(.A(new_n985), .ZN(new_n987));
  NAND4_X1  g801(.A1(new_n973), .A2(new_n982), .A3(new_n987), .A4(new_n983), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n986), .A2(new_n988), .ZN(G72));
  NAND3_X1  g803(.A1(new_n966), .A2(new_n953), .A3(new_n969), .ZN(new_n990));
  NAND2_X1  g804(.A1(G472), .A2(G902), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n991), .B(KEYINPUT63), .Z(new_n992));
  NAND2_X1  g806(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  INV_X1    g807(.A(new_n604), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n994), .A2(new_n605), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n996), .A2(new_n894), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n975), .A2(new_n953), .A3(new_n977), .A4(new_n980), .ZN(new_n998));
  AOI211_X1 g812(.A(new_n569), .B(new_n604), .C1(new_n998), .C2(new_n992), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n994), .A2(new_n569), .ZN(new_n1000));
  OAI211_X1 g814(.A(new_n895), .B(new_n992), .C1(new_n709), .C2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1001), .A2(KEYINPUT127), .ZN(new_n1002));
  OR2_X1    g816(.A1(new_n1001), .A2(KEYINPUT127), .ZN(new_n1003));
  AOI211_X1 g817(.A(new_n997), .B(new_n999), .C1(new_n1002), .C2(new_n1003), .ZN(G57));
endmodule


