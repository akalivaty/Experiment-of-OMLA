//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 0 1 0 0 0 1 1 1 0 0 0 0 0 1 0 0 0 1 1 1 0 1 0 1 1 0 0 1 1 0 0 0 0 0 1 0 0 0 1 0 1 1 0 1 0 0 1 1 1 0 1 1 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:33 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  NOR2_X1   g001(.A1(G237), .A2(G953), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G210), .ZN(new_n189));
  INV_X1    g003(.A(G101), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n192));
  XOR2_X1   g006(.A(new_n191), .B(new_n192), .Z(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT71), .ZN(new_n195));
  AND2_X1   g009(.A1(KEYINPUT64), .A2(G146), .ZN(new_n196));
  NOR2_X1   g010(.A1(KEYINPUT64), .A2(G146), .ZN(new_n197));
  OAI21_X1  g011(.A(G143), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G143), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G146), .ZN(new_n200));
  XNOR2_X1  g014(.A(KEYINPUT68), .B(KEYINPUT1), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n198), .A2(G128), .A3(new_n200), .A4(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G128), .ZN(new_n203));
  XOR2_X1   g017(.A(KEYINPUT68), .B(KEYINPUT1), .Z(new_n204));
  AOI21_X1  g018(.A(new_n203), .B1(new_n204), .B2(new_n198), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n199), .A2(G146), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n196), .A2(new_n197), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n206), .B1(new_n207), .B2(new_n199), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n202), .B1(new_n205), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G137), .ZN(new_n210));
  AND3_X1   g024(.A1(new_n210), .A2(KEYINPUT11), .A3(G134), .ZN(new_n211));
  INV_X1    g025(.A(G134), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(KEYINPUT66), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT66), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G134), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n211), .B1(new_n216), .B2(G137), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n213), .A2(new_n215), .A3(new_n210), .ZN(new_n218));
  AND2_X1   g032(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n219));
  NOR2_X1   g033(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n218), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G131), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n217), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n212), .A2(G137), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n218), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G131), .ZN(new_n227));
  AND3_X1   g041(.A1(new_n209), .A2(new_n224), .A3(new_n227), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n198), .A2(KEYINPUT0), .A3(G128), .A4(new_n200), .ZN(new_n229));
  XOR2_X1   g043(.A(KEYINPUT0), .B(G128), .Z(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n229), .B1(new_n208), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n217), .A2(new_n222), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G131), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n232), .B1(new_n234), .B2(new_n224), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n195), .B1(new_n228), .B2(new_n235), .ZN(new_n236));
  XNOR2_X1  g050(.A(KEYINPUT2), .B(G113), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  XNOR2_X1  g052(.A(G116), .B(G119), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n239), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(new_n237), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  AND3_X1   g058(.A1(new_n198), .A2(G128), .A3(new_n200), .ZN(new_n245));
  INV_X1    g059(.A(new_n206), .ZN(new_n246));
  OR2_X1    g060(.A1(KEYINPUT64), .A2(G146), .ZN(new_n247));
  NAND2_X1  g061(.A1(KEYINPUT64), .A2(G146), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n246), .B1(new_n249), .B2(G143), .ZN(new_n250));
  AOI22_X1  g064(.A1(new_n245), .A2(KEYINPUT0), .B1(new_n250), .B2(new_n230), .ZN(new_n251));
  INV_X1    g065(.A(new_n224), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n223), .B1(new_n217), .B2(new_n222), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n251), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n209), .A2(new_n224), .A3(new_n227), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n254), .A2(KEYINPUT71), .A3(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n236), .A2(new_n244), .A3(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT28), .ZN(new_n258));
  AND2_X1   g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n224), .A2(KEYINPUT67), .A3(new_n227), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(new_n209), .ZN(new_n261));
  AOI21_X1  g075(.A(KEYINPUT67), .B1(new_n224), .B2(new_n227), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n254), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(new_n243), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n255), .A2(KEYINPUT69), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT69), .ZN(new_n266));
  NAND4_X1  g080(.A1(new_n209), .A2(new_n266), .A3(new_n224), .A4(new_n227), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n265), .A2(new_n244), .A3(new_n254), .A4(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n258), .B1(new_n264), .B2(new_n268), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n194), .B1(new_n259), .B2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT72), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n264), .A2(new_n268), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(KEYINPUT28), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n257), .A2(new_n258), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n276), .A2(KEYINPUT72), .A3(new_n194), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT30), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n263), .A2(new_n278), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n265), .A2(KEYINPUT30), .A3(new_n254), .A4(new_n267), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n279), .A2(new_n243), .A3(new_n280), .ZN(new_n281));
  AND2_X1   g095(.A1(new_n281), .A2(new_n268), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n282), .A2(KEYINPUT70), .A3(KEYINPUT31), .A4(new_n193), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n281), .A2(KEYINPUT70), .A3(new_n268), .A4(new_n193), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT31), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AOI22_X1  g100(.A1(new_n272), .A2(new_n277), .B1(new_n283), .B2(new_n286), .ZN(new_n287));
  NOR2_X1   g101(.A1(G472), .A2(G902), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n187), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(KEYINPUT72), .B1(new_n276), .B2(new_n194), .ZN(new_n291));
  AOI211_X1 g105(.A(new_n271), .B(new_n193), .C1(new_n274), .C2(new_n275), .ZN(new_n292));
  AND2_X1   g106(.A1(new_n284), .A2(new_n285), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n284), .A2(new_n285), .ZN(new_n294));
  OAI22_X1  g108(.A1(new_n291), .A2(new_n292), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n295), .A2(KEYINPUT32), .A3(new_n288), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n276), .A2(new_n194), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n282), .A2(new_n193), .ZN(new_n298));
  NOR3_X1   g112(.A1(new_n297), .A2(new_n298), .A3(KEYINPUT29), .ZN(new_n299));
  INV_X1    g113(.A(G902), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n265), .A2(new_n254), .A3(new_n267), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(new_n243), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(new_n268), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(KEYINPUT28), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(new_n275), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n193), .A2(KEYINPUT29), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n300), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  OAI21_X1  g121(.A(G472), .B1(new_n299), .B2(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n290), .A2(new_n296), .A3(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(G234), .ZN(new_n310));
  OAI21_X1  g124(.A(G217), .B1(new_n310), .B2(G902), .ZN(new_n311));
  XNOR2_X1  g125(.A(new_n311), .B(KEYINPUT73), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G146), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT16), .ZN(new_n315));
  INV_X1    g129(.A(G140), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n315), .A2(new_n316), .A3(G125), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(KEYINPUT75), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n316), .A2(G125), .ZN(new_n319));
  INV_X1    g133(.A(G125), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(G140), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n318), .B1(new_n322), .B2(new_n315), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT75), .ZN(new_n325));
  NOR3_X1   g139(.A1(new_n322), .A2(new_n325), .A3(new_n315), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n314), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n322), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n328), .A2(KEYINPUT75), .A3(KEYINPUT16), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n329), .A2(G146), .A3(new_n323), .ZN(new_n330));
  AND2_X1   g144(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  XOR2_X1   g145(.A(KEYINPUT24), .B(G110), .Z(new_n332));
  XNOR2_X1  g146(.A(new_n332), .B(KEYINPUT74), .ZN(new_n333));
  XNOR2_X1  g147(.A(G119), .B(G128), .ZN(new_n334));
  AND2_X1   g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT23), .ZN(new_n336));
  INV_X1    g150(.A(G119), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n336), .B1(new_n337), .B2(G128), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n203), .A2(G119), .ZN(new_n339));
  MUX2_X1   g153(.A(new_n336), .B(new_n338), .S(new_n339), .Z(new_n340));
  INV_X1    g154(.A(G110), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NOR3_X1   g156(.A1(new_n331), .A2(new_n335), .A3(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n340), .A2(new_n341), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n345), .B1(new_n333), .B2(new_n334), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n328), .A2(new_n249), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n346), .A2(new_n330), .A3(new_n347), .ZN(new_n348));
  XNOR2_X1  g162(.A(KEYINPUT22), .B(G137), .ZN(new_n349));
  INV_X1    g163(.A(G221), .ZN(new_n350));
  NOR3_X1   g164(.A1(new_n350), .A2(new_n310), .A3(G953), .ZN(new_n351));
  XOR2_X1   g165(.A(new_n349), .B(new_n351), .Z(new_n352));
  NAND3_X1  g166(.A1(new_n344), .A2(new_n348), .A3(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n352), .ZN(new_n354));
  INV_X1    g168(.A(new_n348), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n354), .B1(new_n343), .B2(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n353), .A2(new_n356), .A3(new_n300), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT25), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n353), .A2(new_n356), .A3(KEYINPUT25), .A4(new_n300), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n313), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n353), .A2(new_n356), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n312), .A2(G902), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n361), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n309), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(KEYINPUT76), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n347), .B1(new_n314), .B2(new_n328), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n188), .A2(G214), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n199), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n188), .A2(G143), .A3(G214), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT18), .ZN(new_n373));
  OAI211_X1 g187(.A(new_n371), .B(new_n372), .C1(new_n373), .C2(new_n223), .ZN(new_n374));
  INV_X1    g188(.A(new_n372), .ZN(new_n375));
  AOI21_X1  g189(.A(G143), .B1(new_n188), .B2(G214), .ZN(new_n376));
  OAI21_X1  g190(.A(G131), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  OAI211_X1 g191(.A(new_n369), .B(new_n374), .C1(new_n373), .C2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT17), .ZN(new_n379));
  OAI211_X1 g193(.A(new_n327), .B(new_n330), .C1(new_n379), .C2(new_n377), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n371), .A2(new_n223), .A3(new_n372), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n377), .A2(new_n381), .A3(new_n379), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT88), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n377), .A2(new_n381), .A3(KEYINPUT88), .A4(new_n379), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n378), .B1(new_n380), .B2(new_n386), .ZN(new_n387));
  XNOR2_X1  g201(.A(G113), .B(G122), .ZN(new_n388));
  XNOR2_X1  g202(.A(new_n388), .B(G104), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  OR2_X1    g204(.A1(new_n390), .A2(KEYINPUT89), .ZN(new_n391));
  AOI21_X1  g205(.A(G902), .B1(new_n387), .B2(new_n391), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n392), .B1(new_n387), .B2(new_n391), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(G475), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT20), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n377), .A2(new_n381), .ZN(new_n396));
  OR2_X1    g210(.A1(new_n322), .A2(KEYINPUT19), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n322), .A2(KEYINPUT19), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n397), .A2(new_n249), .A3(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n330), .A2(new_n396), .A3(new_n399), .ZN(new_n400));
  AND3_X1   g214(.A1(new_n378), .A2(new_n389), .A3(new_n400), .ZN(new_n401));
  AOI211_X1 g215(.A(G475), .B(new_n401), .C1(new_n387), .C2(new_n390), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n395), .B1(new_n402), .B2(new_n300), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n401), .B1(new_n387), .B2(new_n390), .ZN(new_n404));
  INV_X1    g218(.A(G475), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n404), .A2(new_n395), .A3(new_n405), .A4(new_n300), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n394), .B1(new_n403), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  XNOR2_X1  g223(.A(G128), .B(G143), .ZN(new_n410));
  AND2_X1   g224(.A1(new_n216), .A2(new_n410), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n216), .A2(new_n410), .ZN(new_n412));
  OR3_X1    g226(.A1(new_n411), .A2(new_n412), .A3(KEYINPUT91), .ZN(new_n413));
  XNOR2_X1  g227(.A(G116), .B(G122), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT14), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(G107), .ZN(new_n417));
  INV_X1    g231(.A(G122), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n418), .A2(G116), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n417), .B1(new_n419), .B2(KEYINPUT14), .ZN(new_n420));
  AOI22_X1  g234(.A1(new_n416), .A2(new_n420), .B1(new_n417), .B2(new_n414), .ZN(new_n421));
  OAI21_X1  g235(.A(KEYINPUT91), .B1(new_n411), .B2(new_n412), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n413), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  OR2_X1    g237(.A1(new_n411), .A2(KEYINPUT90), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT13), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n425), .A2(new_n199), .A3(G128), .ZN(new_n426));
  INV_X1    g240(.A(new_n410), .ZN(new_n427));
  OAI211_X1 g241(.A(G134), .B(new_n426), .C1(new_n427), .C2(new_n425), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n414), .B(new_n417), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n411), .A2(KEYINPUT90), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n424), .A2(new_n428), .A3(new_n429), .A4(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n423), .A2(new_n431), .ZN(new_n432));
  XOR2_X1   g246(.A(KEYINPUT9), .B(G234), .Z(new_n433));
  INV_X1    g247(.A(G953), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n433), .A2(G217), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n432), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n435), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n423), .A2(new_n437), .A3(new_n431), .ZN(new_n438));
  AOI21_X1  g252(.A(G902), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(G478), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n440), .A2(KEYINPUT15), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n439), .B(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n409), .A2(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(G214), .B1(G237), .B2(G902), .ZN(new_n444));
  XOR2_X1   g258(.A(new_n444), .B(KEYINPUT82), .Z(new_n445));
  XOR2_X1   g259(.A(new_n445), .B(KEYINPUT83), .Z(new_n446));
  INV_X1    g260(.A(G104), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(G107), .ZN(new_n448));
  AND3_X1   g262(.A1(new_n417), .A2(KEYINPUT3), .A3(G104), .ZN(new_n449));
  AOI21_X1  g263(.A(KEYINPUT3), .B1(new_n417), .B2(G104), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n448), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(G101), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n190), .B(new_n448), .C1(new_n449), .C2(new_n450), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n452), .A2(KEYINPUT4), .A3(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT4), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n451), .A2(new_n455), .A3(G101), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n454), .A2(new_n243), .A3(new_n456), .ZN(new_n457));
  XOR2_X1   g271(.A(G110), .B(G122), .Z(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(KEYINPUT78), .B1(new_n417), .B2(G104), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT78), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n461), .A2(new_n447), .A3(G107), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n417), .A2(G104), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n460), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(G101), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT79), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n465), .A2(new_n466), .A3(new_n453), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n466), .B1(new_n465), .B2(new_n453), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(G113), .ZN(new_n471));
  XNOR2_X1  g285(.A(KEYINPUT84), .B(KEYINPUT5), .ZN(new_n472));
  AND2_X1   g286(.A1(new_n337), .A2(G116), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n474), .B1(new_n241), .B2(new_n472), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(new_n240), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n457), .B(new_n459), .C1(new_n470), .C2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n232), .A2(G125), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n434), .A2(G224), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(KEYINPUT7), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n478), .B(new_n481), .C1(G125), .C2(new_n209), .ZN(new_n482));
  AND2_X1   g296(.A1(new_n477), .A2(new_n482), .ZN(new_n483));
  XOR2_X1   g297(.A(new_n458), .B(KEYINPUT8), .Z(new_n484));
  INV_X1    g298(.A(KEYINPUT5), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n474), .B1(new_n485), .B2(new_n241), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(new_n240), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n465), .A2(new_n453), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(KEYINPUT79), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n487), .B1(new_n489), .B2(new_n467), .ZN(new_n490));
  AND2_X1   g304(.A1(new_n476), .A2(new_n488), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n484), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT86), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n478), .B1(G125), .B2(new_n209), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n480), .ZN(new_n496));
  OAI211_X1 g310(.A(KEYINPUT86), .B(new_n484), .C1(new_n490), .C2(new_n491), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n483), .A2(new_n494), .A3(new_n496), .A4(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n476), .B1(new_n489), .B2(new_n467), .ZN(new_n499));
  INV_X1    g313(.A(new_n457), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n458), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n501), .A2(KEYINPUT6), .A3(new_n477), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT6), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n503), .B(new_n458), .C1(new_n499), .C2(new_n500), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n479), .B(KEYINPUT85), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n495), .B(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n502), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n498), .A2(new_n507), .A3(new_n300), .ZN(new_n508));
  OAI21_X1  g322(.A(G210), .B1(G237), .B2(G902), .ZN(new_n509));
  XOR2_X1   g323(.A(new_n509), .B(KEYINPUT87), .Z(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n498), .A2(new_n507), .A3(new_n300), .A4(new_n510), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(G234), .A2(G237), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n515), .A2(G952), .A3(new_n434), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n516), .B(KEYINPUT92), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  XOR2_X1   g332(.A(KEYINPUT21), .B(G898), .Z(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n515), .A2(G902), .A3(G953), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n518), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  NOR4_X1   g337(.A1(new_n443), .A2(new_n446), .A3(new_n514), .A4(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n350), .B1(new_n433), .B2(new_n300), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  AND2_X1   g340(.A1(new_n198), .A2(new_n200), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n203), .B1(new_n246), .B2(KEYINPUT1), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n202), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n529), .A2(new_n453), .A3(new_n465), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT10), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  OAI211_X1 g346(.A(KEYINPUT10), .B(new_n209), .C1(new_n468), .C2(new_n469), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n251), .A2(new_n456), .A3(new_n454), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n252), .A2(new_n253), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n532), .A2(new_n533), .A3(new_n536), .A4(new_n534), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n434), .A2(G227), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n541), .B(new_n316), .ZN(new_n542));
  XNOR2_X1  g356(.A(KEYINPUT77), .B(G110), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n542), .B(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n540), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n199), .B1(new_n247), .B2(new_n248), .ZN(new_n547));
  OAI21_X1  g361(.A(G128), .B1(new_n547), .B2(new_n201), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(new_n250), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n489), .A2(new_n549), .A3(new_n202), .A4(new_n467), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(KEYINPUT80), .ZN(new_n551));
  AOI22_X1  g365(.A1(new_n245), .A2(new_n201), .B1(new_n548), .B2(new_n250), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT80), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n552), .A2(new_n553), .A3(new_n489), .A4(new_n467), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n551), .A2(new_n530), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(new_n537), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(KEYINPUT12), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT12), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n555), .A2(new_n558), .A3(new_n537), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n557), .A2(new_n539), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n546), .B1(new_n560), .B2(new_n545), .ZN(new_n561));
  OAI21_X1  g375(.A(G469), .B1(new_n561), .B2(G902), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(KEYINPUT81), .ZN(new_n563));
  NAND4_X1  g377(.A1(new_n557), .A2(new_n539), .A3(new_n544), .A4(new_n559), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n540), .A2(new_n545), .ZN(new_n565));
  AOI21_X1  g379(.A(G902), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(G469), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT81), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n569), .B(G469), .C1(new_n561), .C2(G902), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n563), .A2(new_n568), .A3(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n524), .A2(new_n526), .A3(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT76), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n309), .A2(new_n574), .A3(new_n366), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n368), .A2(new_n573), .A3(new_n575), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n576), .B(G101), .ZN(G3));
  INV_X1    g391(.A(G472), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n578), .B1(new_n295), .B2(new_n300), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n287), .A2(new_n289), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n366), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n582), .A2(new_n525), .ZN(new_n583));
  AND3_X1   g397(.A1(new_n581), .A2(new_n583), .A3(new_n571), .ZN(new_n584));
  INV_X1    g398(.A(new_n445), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n514), .A2(new_n523), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n404), .A2(new_n405), .A3(new_n300), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(KEYINPUT20), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(new_n406), .ZN(new_n590));
  INV_X1    g404(.A(new_n439), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n591), .A2(KEYINPUT94), .A3(new_n440), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT94), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n593), .B1(new_n439), .B2(G478), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n436), .A2(new_n438), .ZN(new_n596));
  OAI21_X1  g410(.A(KEYINPUT33), .B1(new_n437), .B2(KEYINPUT93), .ZN(new_n597));
  OR2_X1    g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n596), .A2(new_n597), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n440), .A2(G902), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  AOI22_X1  g415(.A1(new_n590), .A2(new_n394), .B1(new_n595), .B2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n587), .A2(new_n603), .ZN(new_n604));
  XOR2_X1   g418(.A(KEYINPUT34), .B(G104), .Z(new_n605));
  XNOR2_X1  g419(.A(new_n605), .B(KEYINPUT95), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n604), .B(new_n606), .ZN(G6));
  XNOR2_X1  g421(.A(new_n406), .B(KEYINPUT96), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n589), .ZN(new_n609));
  INV_X1    g423(.A(new_n442), .ZN(new_n610));
  AND3_X1   g424(.A1(new_n609), .A2(new_n394), .A3(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n587), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(KEYINPUT35), .B(G107), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(G9));
  NAND2_X1  g429(.A1(new_n344), .A2(new_n348), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n354), .A2(KEYINPUT36), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n361), .B1(new_n363), .B2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n581), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n572), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(KEYINPUT37), .B(G110), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(G12));
  AND2_X1   g438(.A1(new_n571), .A2(new_n526), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n512), .A2(new_n585), .A3(new_n513), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(G900), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n518), .B1(new_n628), .B2(new_n522), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  AND3_X1   g444(.A1(new_n611), .A2(new_n627), .A3(new_n630), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n625), .A2(new_n631), .A3(new_n309), .A4(new_n620), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(G128), .ZN(G30));
  NAND2_X1  g447(.A1(new_n282), .A2(new_n193), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n303), .A2(new_n194), .ZN(new_n635));
  AND2_X1   g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  OAI21_X1  g450(.A(G472), .B1(new_n636), .B2(G902), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n290), .A2(new_n296), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(KEYINPUT97), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT97), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n290), .A2(new_n640), .A3(new_n296), .A4(new_n637), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(KEYINPUT98), .ZN(new_n643));
  XOR2_X1   g457(.A(new_n629), .B(KEYINPUT39), .Z(new_n644));
  NAND2_X1  g458(.A1(new_n625), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n643), .B1(KEYINPUT40), .B2(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n645), .A2(KEYINPUT40), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n408), .A2(new_n610), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n514), .B(KEYINPUT38), .ZN(new_n651));
  NOR4_X1   g465(.A1(new_n650), .A2(new_n445), .A3(new_n620), .A4(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(new_n199), .ZN(G45));
  NAND4_X1  g467(.A1(new_n309), .A2(new_n526), .A3(new_n571), .A4(new_n620), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n602), .A2(new_n630), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT99), .ZN(new_n656));
  NOR3_X1   g470(.A1(new_n655), .A2(new_n656), .A3(new_n626), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n656), .B1(new_n655), .B2(new_n626), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  OR3_X1    g473(.A1(new_n654), .A2(new_n657), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G146), .ZN(G48));
  NAND2_X1  g475(.A1(new_n564), .A2(new_n565), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n300), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(G469), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n664), .A2(new_n602), .A3(new_n526), .A4(new_n568), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n586), .A2(new_n585), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n667), .A2(new_n309), .A3(new_n366), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT100), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n667), .A2(new_n309), .A3(KEYINPUT100), .A4(new_n366), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(KEYINPUT41), .B(G113), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G15));
  NAND3_X1  g488(.A1(new_n664), .A2(new_n526), .A3(new_n568), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n675), .A2(new_n626), .ZN(new_n676));
  INV_X1    g490(.A(new_n523), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n609), .A2(new_n394), .A3(new_n610), .A4(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n678), .A2(new_n582), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n309), .A2(new_n676), .A3(new_n679), .ZN(new_n680));
  XOR2_X1   g494(.A(KEYINPUT101), .B(G116), .Z(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G18));
  NOR3_X1   g496(.A1(new_n619), .A2(new_n443), .A3(new_n523), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n309), .A2(new_n676), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G119), .ZN(G21));
  AOI21_X1  g499(.A(new_n442), .B1(new_n590), .B2(new_n394), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n686), .A2(new_n585), .A3(new_n513), .A4(new_n512), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n675), .A2(new_n687), .A3(new_n523), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n283), .A2(new_n286), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n305), .A2(new_n194), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n289), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n579), .A2(new_n691), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n688), .A2(KEYINPUT102), .A3(new_n366), .A4(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT102), .ZN(new_n694));
  INV_X1    g508(.A(new_n691), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n272), .A2(new_n277), .ZN(new_n696));
  AOI21_X1  g510(.A(G902), .B1(new_n696), .B2(new_n689), .ZN(new_n697));
  OAI211_X1 g511(.A(new_n695), .B(new_n366), .C1(new_n697), .C2(new_n578), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n566), .B(G469), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n648), .A2(new_n626), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n699), .A2(new_n700), .A3(new_n526), .A4(new_n677), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n694), .B1(new_n698), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n693), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G122), .ZN(G24));
  INV_X1    g518(.A(new_n655), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n692), .A2(new_n676), .A3(new_n620), .A4(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G125), .ZN(G27));
  INV_X1    g521(.A(KEYINPUT103), .ZN(new_n708));
  AND3_X1   g522(.A1(new_n555), .A2(new_n558), .A3(new_n537), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n558), .B1(new_n555), .B2(new_n537), .ZN(new_n710));
  INV_X1    g524(.A(new_n539), .ZN(new_n711));
  NOR3_X1   g525(.A1(new_n709), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n708), .B1(new_n712), .B2(new_n544), .ZN(new_n713));
  INV_X1    g527(.A(new_n546), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n560), .A2(KEYINPUT103), .A3(new_n545), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n713), .A2(G469), .A3(new_n714), .A4(new_n715), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n567), .A2(new_n300), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n717), .B1(new_n566), .B2(new_n567), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n526), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT104), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n445), .B1(new_n512), .B2(new_n513), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n525), .B1(new_n716), .B2(new_n718), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(KEYINPUT104), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n722), .A2(new_n723), .A3(new_n725), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n726), .A2(new_n367), .ZN(new_n727));
  NOR2_X1   g541(.A1(KEYINPUT105), .A2(KEYINPUT42), .ZN(new_n728));
  INV_X1    g542(.A(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n727), .A2(new_n705), .A3(new_n729), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n724), .A2(KEYINPUT104), .ZN(new_n731));
  AOI211_X1 g545(.A(new_n721), .B(new_n525), .C1(new_n716), .C2(new_n718), .ZN(new_n732));
  INV_X1    g546(.A(new_n723), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n731), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  AND2_X1   g548(.A1(new_n309), .A2(new_n366), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n734), .A2(new_n735), .A3(new_n705), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(new_n728), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n730), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G131), .ZN(G33));
  NOR2_X1   g553(.A1(new_n612), .A2(new_n629), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n734), .A2(new_n735), .A3(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G134), .ZN(G36));
  OR2_X1    g556(.A1(new_n561), .A2(KEYINPUT45), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n713), .A2(new_n714), .A3(new_n715), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT45), .ZN(new_n745));
  OAI211_X1 g559(.A(new_n743), .B(G469), .C1(new_n744), .C2(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(new_n717), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n746), .A2(KEYINPUT46), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(new_n568), .ZN(new_n749));
  AOI21_X1  g563(.A(KEYINPUT46), .B1(new_n746), .B2(new_n747), .ZN(new_n750));
  OR2_X1    g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  AND2_X1   g565(.A1(new_n751), .A2(new_n526), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(new_n644), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n595), .A2(new_n601), .ZN(new_n755));
  AOI21_X1  g569(.A(KEYINPUT106), .B1(new_n409), .B2(new_n755), .ZN(new_n756));
  XOR2_X1   g570(.A(new_n756), .B(KEYINPUT43), .Z(new_n757));
  OAI211_X1 g571(.A(new_n757), .B(new_n620), .C1(new_n580), .C2(new_n579), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT44), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n733), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  OAI211_X1 g574(.A(new_n754), .B(new_n760), .C1(new_n759), .C2(new_n758), .ZN(new_n761));
  XNOR2_X1  g575(.A(KEYINPUT107), .B(G137), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n761), .B(new_n762), .ZN(G39));
  NAND2_X1  g577(.A1(new_n751), .A2(new_n526), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT47), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n764), .B(new_n765), .ZN(new_n766));
  NOR3_X1   g580(.A1(new_n309), .A2(new_n366), .A3(new_n733), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n766), .A2(new_n705), .A3(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G140), .ZN(G42));
  INV_X1    g583(.A(new_n643), .ZN(new_n770));
  INV_X1    g584(.A(new_n699), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n770), .B1(KEYINPUT49), .B2(new_n771), .ZN(new_n772));
  OR2_X1    g586(.A1(new_n771), .A2(KEYINPUT49), .ZN(new_n773));
  INV_X1    g587(.A(new_n446), .ZN(new_n774));
  AND4_X1   g588(.A1(new_n409), .A2(new_n651), .A3(new_n774), .A4(new_n755), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n772), .A2(new_n583), .A3(new_n773), .A4(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n757), .A2(new_n518), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(KEYINPUT111), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT111), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n757), .A2(new_n779), .A3(new_n518), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n698), .B1(new_n778), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n771), .A2(new_n526), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n723), .B(new_n781), .C1(new_n766), .C2(new_n782), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n675), .A2(new_n733), .ZN(new_n784));
  AND4_X1   g598(.A1(new_n366), .A2(new_n643), .A3(new_n518), .A4(new_n784), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n785), .A2(new_n409), .A3(new_n595), .A4(new_n601), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n699), .A2(new_n526), .A3(new_n445), .ZN(new_n787));
  OR2_X1    g601(.A1(new_n787), .A2(KEYINPUT112), .ZN(new_n788));
  INV_X1    g602(.A(new_n651), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n789), .B1(new_n787), .B2(KEYINPUT112), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n781), .A2(new_n788), .A3(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT50), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n781), .A2(KEYINPUT50), .A3(new_n788), .A4(new_n790), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  AOI211_X1 g609(.A(new_n675), .B(new_n733), .C1(new_n778), .C2(new_n780), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n796), .A2(new_n620), .A3(new_n692), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n783), .A2(new_n786), .A3(new_n795), .A4(new_n797), .ZN(new_n798));
  AOI21_X1  g612(.A(KEYINPUT51), .B1(new_n783), .B2(KEYINPUT113), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n798), .B(new_n799), .ZN(new_n800));
  OAI211_X1 g614(.A(new_n309), .B(new_n676), .C1(new_n683), .C2(new_n679), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n672), .A2(new_n703), .A3(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT108), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n602), .A2(new_n803), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n803), .B1(new_n408), .B2(new_n442), .ZN(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n804), .B1(new_n806), .B2(new_n602), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n584), .A2(new_n774), .A3(new_n586), .A4(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(new_n622), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n576), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n802), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n610), .A2(new_n629), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n620), .A2(new_n394), .A3(new_n609), .A4(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n813), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n814), .A2(new_n625), .A3(new_n309), .A4(new_n723), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n741), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n692), .A2(new_n620), .A3(new_n705), .ZN(new_n817));
  OAI21_X1  g631(.A(KEYINPUT109), .B1(new_n726), .B2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(new_n817), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT109), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n734), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n816), .B1(new_n818), .B2(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n811), .A2(new_n822), .A3(new_n738), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT53), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n625), .A2(new_n309), .A3(new_n620), .A4(new_n658), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n632), .B(new_n706), .C1(new_n825), .C2(new_n657), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n620), .A2(new_n629), .A3(new_n687), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n642), .A2(new_n724), .A3(new_n827), .ZN(new_n828));
  OAI21_X1  g642(.A(KEYINPUT52), .B1(new_n826), .B2(new_n828), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n632), .A2(new_n706), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n642), .A2(new_n724), .A3(new_n827), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT52), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n830), .A2(new_n660), .A3(new_n831), .A4(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n829), .A2(new_n833), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n823), .A2(new_n824), .A3(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n309), .A2(new_n526), .A3(new_n571), .A4(new_n723), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n836), .A2(new_n813), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n837), .B1(new_n727), .B2(new_n740), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n821), .A2(new_n818), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n729), .B1(new_n727), .B2(new_n705), .ZN(new_n840));
  NOR4_X1   g654(.A1(new_n726), .A2(new_n367), .A3(new_n655), .A4(new_n728), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n838), .B(new_n839), .C1(new_n840), .C2(new_n841), .ZN(new_n842));
  AND3_X1   g656(.A1(new_n309), .A2(new_n574), .A3(new_n366), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n574), .B1(new_n309), .B2(new_n366), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n622), .B1(new_n845), .B2(new_n573), .ZN(new_n846));
  INV_X1    g660(.A(new_n801), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n847), .B1(new_n702), .B2(new_n693), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n846), .A2(new_n672), .A3(new_n848), .A4(new_n808), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n842), .A2(new_n849), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n829), .A2(new_n833), .ZN(new_n851));
  AOI21_X1  g665(.A(KEYINPUT53), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g666(.A(KEYINPUT54), .B1(new_n835), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n781), .A2(new_n676), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n824), .B1(new_n823), .B2(new_n834), .ZN(new_n855));
  INV_X1    g669(.A(new_n842), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n810), .B1(new_n802), .B2(KEYINPUT110), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT110), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n672), .A2(new_n858), .A3(new_n703), .A4(new_n801), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n859), .A2(KEYINPUT53), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n851), .A2(new_n856), .A3(new_n857), .A4(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT54), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n855), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n434), .A2(G952), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n864), .B1(new_n785), .B2(new_n602), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n853), .A2(new_n854), .A3(new_n863), .A4(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n796), .A2(new_n735), .ZN(new_n867));
  XOR2_X1   g681(.A(new_n867), .B(KEYINPUT48), .Z(new_n868));
  NOR3_X1   g682(.A1(new_n800), .A2(new_n866), .A3(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(G952), .A2(G953), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n776), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT114), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OAI211_X1 g687(.A(KEYINPUT114), .B(new_n776), .C1(new_n869), .C2(new_n870), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(G75));
  XNOR2_X1  g689(.A(KEYINPUT115), .B(KEYINPUT55), .ZN(new_n876));
  INV_X1    g690(.A(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n300), .B1(new_n855), .B2(new_n861), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n878), .A2(new_n510), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT56), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n877), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  AOI211_X1 g695(.A(KEYINPUT56), .B(new_n876), .C1(new_n878), .C2(new_n510), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n502), .A2(new_n504), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n884), .B(new_n506), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n434), .A2(G952), .ZN(new_n887));
  INV_X1    g701(.A(new_n885), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n881), .A2(new_n882), .A3(new_n888), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n886), .A2(new_n887), .A3(new_n889), .ZN(G51));
  XOR2_X1   g704(.A(new_n746), .B(KEYINPUT117), .Z(new_n891));
  AND2_X1   g705(.A1(new_n878), .A2(new_n891), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n670), .A2(new_n671), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n703), .A2(new_n801), .ZN(new_n894));
  OAI21_X1  g708(.A(KEYINPUT110), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  AND3_X1   g709(.A1(new_n576), .A2(new_n808), .A3(new_n809), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n895), .A2(KEYINPUT53), .A3(new_n896), .A4(new_n859), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n897), .A2(new_n834), .A3(new_n842), .ZN(new_n898));
  OAI21_X1  g712(.A(KEYINPUT54), .B1(new_n852), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(new_n863), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n717), .B(KEYINPUT57), .Z(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(KEYINPUT116), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT116), .ZN(new_n904));
  AOI211_X1 g718(.A(new_n904), .B(new_n901), .C1(new_n899), .C2(new_n863), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n892), .B1(new_n906), .B2(new_n662), .ZN(new_n907));
  OAI21_X1  g721(.A(KEYINPUT118), .B1(new_n907), .B2(new_n887), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT118), .ZN(new_n909));
  INV_X1    g723(.A(new_n887), .ZN(new_n910));
  INV_X1    g724(.A(new_n662), .ZN(new_n911));
  NOR3_X1   g725(.A1(new_n903), .A2(new_n905), .A3(new_n911), .ZN(new_n912));
  OAI211_X1 g726(.A(new_n909), .B(new_n910), .C1(new_n912), .C2(new_n892), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n908), .A2(new_n913), .ZN(G54));
  NAND3_X1  g728(.A1(new_n878), .A2(KEYINPUT58), .A3(G475), .ZN(new_n915));
  INV_X1    g729(.A(new_n404), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n917), .B(KEYINPUT119), .Z(new_n918));
  OAI21_X1  g732(.A(new_n910), .B1(new_n915), .B2(new_n916), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n918), .A2(new_n919), .ZN(G60));
  INV_X1    g734(.A(new_n900), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n598), .A2(new_n599), .ZN(new_n922));
  NAND2_X1  g736(.A1(G478), .A2(G902), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n923), .B(KEYINPUT59), .Z(new_n924));
  OR3_X1    g738(.A1(new_n921), .A2(new_n922), .A3(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(new_n922), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n924), .B1(new_n853), .B2(new_n863), .ZN(new_n927));
  OAI211_X1 g741(.A(new_n925), .B(new_n910), .C1(new_n926), .C2(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(G63));
  NAND2_X1  g743(.A1(G217), .A2(G902), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n930), .B(KEYINPUT60), .Z(new_n931));
  OAI21_X1  g745(.A(new_n931), .B1(new_n852), .B2(new_n898), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT120), .ZN(new_n933));
  INV_X1    g747(.A(new_n618), .ZN(new_n934));
  OR2_X1    g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n362), .B(KEYINPUT121), .Z(new_n936));
  NAND2_X1  g750(.A1(new_n933), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n935), .A2(new_n910), .A3(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT61), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n935), .A2(new_n937), .A3(KEYINPUT61), .A4(new_n910), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(G66));
  INV_X1    g756(.A(G224), .ZN(new_n943));
  OAI21_X1  g757(.A(G953), .B1(new_n520), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n944), .B1(new_n811), .B2(G953), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT122), .Z(new_n946));
  OAI21_X1  g760(.A(new_n884), .B1(G898), .B2(new_n434), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n946), .B(new_n947), .ZN(G69));
  NAND2_X1  g762(.A1(new_n279), .A2(new_n280), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n949), .B(KEYINPUT123), .Z(new_n950));
  NAND2_X1  g764(.A1(new_n397), .A2(new_n398), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n950), .B(new_n951), .Z(new_n952));
  NAND2_X1  g766(.A1(new_n761), .A2(new_n768), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n845), .A2(new_n807), .ZN(new_n954));
  NOR3_X1   g768(.A1(new_n954), .A2(new_n645), .A3(new_n733), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT62), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n826), .B(KEYINPUT124), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n956), .B1(new_n652), .B2(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(new_n650), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n960), .A2(new_n585), .A3(new_n619), .A4(new_n789), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n961), .A2(KEYINPUT62), .A3(new_n957), .ZN(new_n962));
  AOI211_X1 g776(.A(new_n953), .B(new_n955), .C1(new_n959), .C2(new_n962), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n952), .B1(new_n963), .B2(G953), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n434), .B1(G227), .B2(G900), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(KEYINPUT125), .ZN(new_n966));
  INV_X1    g780(.A(new_n952), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n768), .A2(new_n738), .A3(new_n741), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT126), .ZN(new_n969));
  INV_X1    g783(.A(new_n761), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n969), .B1(new_n970), .B2(new_n958), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n761), .A2(KEYINPUT126), .A3(new_n957), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n968), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n754), .A2(new_n735), .A3(new_n700), .ZN(new_n974));
  AOI21_X1  g788(.A(G953), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n434), .A2(G900), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n967), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  AND3_X1   g791(.A1(new_n964), .A2(new_n966), .A3(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n966), .B1(new_n964), .B2(new_n977), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n978), .A2(new_n979), .ZN(G72));
  XNOR2_X1  g794(.A(new_n282), .B(KEYINPUT127), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(new_n193), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n963), .A2(new_n811), .ZN(new_n983));
  NAND2_X1  g797(.A1(G472), .A2(G902), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n984), .B(KEYINPUT63), .Z(new_n985));
  AOI21_X1  g799(.A(new_n982), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n973), .A2(new_n811), .A3(new_n974), .ZN(new_n987));
  AOI211_X1 g801(.A(new_n193), .B(new_n981), .C1(new_n987), .C2(new_n985), .ZN(new_n988));
  INV_X1    g802(.A(new_n985), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n835), .A2(new_n852), .ZN(new_n990));
  INV_X1    g804(.A(new_n298), .ZN(new_n991));
  AOI211_X1 g805(.A(new_n989), .B(new_n990), .C1(new_n634), .C2(new_n991), .ZN(new_n992));
  NOR4_X1   g806(.A1(new_n986), .A2(new_n988), .A3(new_n887), .A4(new_n992), .ZN(G57));
endmodule


