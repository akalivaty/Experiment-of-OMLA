

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592;

  XNOR2_X1 U324 ( .A(n395), .B(KEYINPUT48), .ZN(n396) );
  XNOR2_X1 U325 ( .A(n483), .B(n482), .ZN(n500) );
  INV_X1 U326 ( .A(KEYINPUT100), .ZN(n482) );
  XOR2_X1 U327 ( .A(KEYINPUT28), .B(n477), .Z(n540) );
  XNOR2_X1 U328 ( .A(n453), .B(n452), .ZN(n455) );
  XNOR2_X1 U329 ( .A(n451), .B(n450), .ZN(n452) );
  XOR2_X1 U330 ( .A(n319), .B(n298), .Z(n292) );
  XOR2_X1 U331 ( .A(KEYINPUT22), .B(KEYINPUT92), .Z(n293) );
  AND2_X1 U332 ( .A1(G227GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U333 ( .A(KEYINPUT99), .B(KEYINPUT26), .ZN(n295) );
  XOR2_X1 U334 ( .A(n443), .B(n408), .Z(n296) );
  XNOR2_X1 U335 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U336 ( .A(n443), .B(n294), .ZN(n444) );
  XNOR2_X1 U337 ( .A(n382), .B(n341), .ZN(n342) );
  XNOR2_X1 U338 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U339 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U340 ( .A(n401), .B(n342), .ZN(n343) );
  NOR2_X1 U341 ( .A1(n590), .A2(n501), .ZN(n502) );
  XOR2_X1 U342 ( .A(n581), .B(KEYINPUT41), .Z(n559) );
  XNOR2_X1 U343 ( .A(n330), .B(n329), .ZN(n586) );
  XOR2_X1 U344 ( .A(n455), .B(n454), .Z(n542) );
  NOR2_X1 U345 ( .A1(n542), .A2(n512), .ZN(n509) );
  XNOR2_X1 U346 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U347 ( .A(n466), .B(n465), .ZN(G1351GAT) );
  XOR2_X1 U348 ( .A(G22GAT), .B(G155GAT), .Z(n319) );
  XNOR2_X1 U349 ( .A(KEYINPUT24), .B(G204GAT), .ZN(n297) );
  XNOR2_X1 U350 ( .A(n293), .B(n297), .ZN(n298) );
  NAND2_X1 U351 ( .A1(G228GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U352 ( .A(n292), .B(n299), .ZN(n300) );
  XOR2_X1 U353 ( .A(n300), .B(G211GAT), .Z(n303) );
  XNOR2_X1 U354 ( .A(G50GAT), .B(KEYINPUT80), .ZN(n301) );
  XNOR2_X1 U355 ( .A(n301), .B(G162GAT), .ZN(n384) );
  XNOR2_X1 U356 ( .A(n384), .B(KEYINPUT23), .ZN(n302) );
  XNOR2_X1 U357 ( .A(n303), .B(n302), .ZN(n305) );
  XNOR2_X1 U358 ( .A(G106GAT), .B(G78GAT), .ZN(n304) );
  XNOR2_X1 U359 ( .A(n304), .B(G148GAT), .ZN(n346) );
  XOR2_X1 U360 ( .A(n305), .B(n346), .Z(n312) );
  XOR2_X1 U361 ( .A(KEYINPUT3), .B(KEYINPUT95), .Z(n307) );
  XNOR2_X1 U362 ( .A(KEYINPUT2), .B(KEYINPUT94), .ZN(n306) );
  XNOR2_X1 U363 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U364 ( .A(G141GAT), .B(n308), .Z(n426) );
  XOR2_X1 U365 ( .A(KEYINPUT21), .B(KEYINPUT93), .Z(n310) );
  XNOR2_X1 U366 ( .A(G197GAT), .B(G218GAT), .ZN(n309) );
  XNOR2_X1 U367 ( .A(n310), .B(n309), .ZN(n400) );
  XNOR2_X1 U368 ( .A(n426), .B(n400), .ZN(n311) );
  XNOR2_X1 U369 ( .A(n312), .B(n311), .ZN(n476) );
  XOR2_X1 U370 ( .A(KEYINPUT87), .B(KEYINPUT83), .Z(n314) );
  XNOR2_X1 U371 ( .A(KEYINPUT85), .B(KEYINPUT86), .ZN(n313) );
  XOR2_X1 U372 ( .A(n314), .B(n313), .Z(n330) );
  XOR2_X1 U373 ( .A(G15GAT), .B(G127GAT), .Z(n443) );
  XNOR2_X1 U374 ( .A(G8GAT), .B(G183GAT), .ZN(n315) );
  XNOR2_X1 U375 ( .A(n315), .B(G211GAT), .ZN(n408) );
  NAND2_X1 U376 ( .A1(G231GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U377 ( .A(n296), .B(n316), .ZN(n323) );
  XOR2_X1 U378 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n318) );
  XNOR2_X1 U379 ( .A(G78GAT), .B(G64GAT), .ZN(n317) );
  XOR2_X1 U380 ( .A(n318), .B(n317), .Z(n321) );
  XOR2_X1 U381 ( .A(G1GAT), .B(KEYINPUT71), .Z(n354) );
  XNOR2_X1 U382 ( .A(n354), .B(n319), .ZN(n320) );
  XOR2_X1 U383 ( .A(n324), .B(KEYINPUT15), .Z(n328) );
  XOR2_X1 U384 ( .A(KEYINPUT13), .B(KEYINPUT72), .Z(n326) );
  XNOR2_X1 U385 ( .A(G71GAT), .B(G57GAT), .ZN(n325) );
  XNOR2_X1 U386 ( .A(n326), .B(n325), .ZN(n345) );
  XNOR2_X1 U387 ( .A(n345), .B(KEYINPUT84), .ZN(n327) );
  XNOR2_X1 U388 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U389 ( .A(n586), .B(KEYINPUT113), .ZN(n568) );
  NAND2_X1 U390 ( .A1(G230GAT), .A2(G233GAT), .ZN(n336) );
  XOR2_X1 U391 ( .A(KEYINPUT31), .B(KEYINPUT74), .Z(n332) );
  XNOR2_X1 U392 ( .A(KEYINPUT73), .B(KEYINPUT78), .ZN(n331) );
  XNOR2_X1 U393 ( .A(n332), .B(n331), .ZN(n334) );
  XOR2_X1 U394 ( .A(G120GAT), .B(KEYINPUT32), .Z(n333) );
  XNOR2_X1 U395 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U396 ( .A(n336), .B(n335), .ZN(n344) );
  XOR2_X1 U397 ( .A(G92GAT), .B(G64GAT), .Z(n338) );
  XNOR2_X1 U398 ( .A(G176GAT), .B(KEYINPUT77), .ZN(n337) );
  XNOR2_X1 U399 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U400 ( .A(G204GAT), .B(n339), .Z(n401) );
  XNOR2_X1 U401 ( .A(G99GAT), .B(G85GAT), .ZN(n340) );
  XNOR2_X1 U402 ( .A(n340), .B(KEYINPUT76), .ZN(n382) );
  XOR2_X1 U403 ( .A(KEYINPUT75), .B(KEYINPUT33), .Z(n341) );
  XNOR2_X1 U404 ( .A(n344), .B(n343), .ZN(n348) );
  XNOR2_X1 U405 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U406 ( .A(n348), .B(n347), .ZN(n581) );
  XOR2_X1 U407 ( .A(KEYINPUT68), .B(G8GAT), .Z(n350) );
  XNOR2_X1 U408 ( .A(G22GAT), .B(G141GAT), .ZN(n349) );
  XNOR2_X1 U409 ( .A(n350), .B(n349), .ZN(n367) );
  XOR2_X1 U410 ( .A(G15GAT), .B(G113GAT), .Z(n352) );
  XNOR2_X1 U411 ( .A(G50GAT), .B(G36GAT), .ZN(n351) );
  XNOR2_X1 U412 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U413 ( .A(n353), .B(G197GAT), .Z(n356) );
  XNOR2_X1 U414 ( .A(G169GAT), .B(n354), .ZN(n355) );
  XNOR2_X1 U415 ( .A(n356), .B(n355), .ZN(n360) );
  XOR2_X1 U416 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n358) );
  NAND2_X1 U417 ( .A1(G229GAT), .A2(G233GAT), .ZN(n357) );
  XNOR2_X1 U418 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U419 ( .A(n360), .B(n359), .Z(n365) );
  XOR2_X1 U420 ( .A(KEYINPUT8), .B(KEYINPUT70), .Z(n362) );
  XNOR2_X1 U421 ( .A(G43GAT), .B(G29GAT), .ZN(n361) );
  XNOR2_X1 U422 ( .A(n362), .B(n361), .ZN(n363) );
  XOR2_X1 U423 ( .A(KEYINPUT7), .B(n363), .Z(n385) );
  XNOR2_X1 U424 ( .A(n385), .B(KEYINPUT69), .ZN(n364) );
  XNOR2_X1 U425 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U426 ( .A(n367), .B(n366), .Z(n574) );
  INV_X1 U427 ( .A(n574), .ZN(n556) );
  NOR2_X1 U428 ( .A1(n559), .A2(n556), .ZN(n368) );
  XNOR2_X1 U429 ( .A(n368), .B(KEYINPUT46), .ZN(n369) );
  NOR2_X1 U430 ( .A1(n568), .A2(n369), .ZN(n388) );
  XOR2_X1 U431 ( .A(KEYINPUT65), .B(KEYINPUT81), .Z(n371) );
  XNOR2_X1 U432 ( .A(KEYINPUT11), .B(KEYINPUT9), .ZN(n370) );
  XNOR2_X1 U433 ( .A(n371), .B(n370), .ZN(n375) );
  XOR2_X1 U434 ( .A(KEYINPUT10), .B(G92GAT), .Z(n373) );
  XNOR2_X1 U435 ( .A(G134GAT), .B(G106GAT), .ZN(n372) );
  XNOR2_X1 U436 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U437 ( .A(n375), .B(n374), .Z(n381) );
  XNOR2_X1 U438 ( .A(G36GAT), .B(G190GAT), .ZN(n376) );
  XNOR2_X1 U439 ( .A(n376), .B(KEYINPUT82), .ZN(n402) );
  XOR2_X1 U440 ( .A(n402), .B(KEYINPUT66), .Z(n378) );
  NAND2_X1 U441 ( .A1(G232GAT), .A2(G233GAT), .ZN(n377) );
  XNOR2_X1 U442 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U443 ( .A(G218GAT), .B(n379), .ZN(n380) );
  XNOR2_X1 U444 ( .A(n381), .B(n380), .ZN(n383) );
  XNOR2_X1 U445 ( .A(n383), .B(n382), .ZN(n387) );
  XNOR2_X1 U446 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U447 ( .A(n387), .B(n386), .ZN(n468) );
  INV_X1 U448 ( .A(n468), .ZN(n565) );
  NAND2_X1 U449 ( .A1(n388), .A2(n565), .ZN(n389) );
  XNOR2_X1 U450 ( .A(n389), .B(KEYINPUT47), .ZN(n394) );
  XOR2_X1 U451 ( .A(KEYINPUT36), .B(n468), .Z(n590) );
  NOR2_X1 U452 ( .A1(n586), .A2(n590), .ZN(n390) );
  XNOR2_X1 U453 ( .A(KEYINPUT45), .B(n390), .ZN(n391) );
  NAND2_X1 U454 ( .A1(n391), .A2(n581), .ZN(n392) );
  NOR2_X1 U455 ( .A1(n392), .A2(n574), .ZN(n393) );
  NOR2_X1 U456 ( .A1(n394), .A2(n393), .ZN(n397) );
  INV_X1 U457 ( .A(KEYINPUT114), .ZN(n395) );
  XNOR2_X1 U458 ( .A(n397), .B(n396), .ZN(n537) );
  XOR2_X1 U459 ( .A(KEYINPUT18), .B(KEYINPUT19), .Z(n399) );
  XNOR2_X1 U460 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n398) );
  XNOR2_X1 U461 ( .A(n399), .B(n398), .ZN(n447) );
  XNOR2_X1 U462 ( .A(n447), .B(n400), .ZN(n406) );
  XOR2_X1 U463 ( .A(n402), .B(n401), .Z(n404) );
  NAND2_X1 U464 ( .A1(G226GAT), .A2(G233GAT), .ZN(n403) );
  XNOR2_X1 U465 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U466 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U467 ( .A(n408), .B(n407), .Z(n490) );
  NAND2_X1 U468 ( .A1(n537), .A2(n490), .ZN(n410) );
  INV_X1 U469 ( .A(KEYINPUT54), .ZN(n409) );
  XNOR2_X1 U470 ( .A(n410), .B(n409), .ZN(n432) );
  XOR2_X1 U471 ( .A(KEYINPUT0), .B(G134GAT), .Z(n412) );
  XNOR2_X1 U472 ( .A(KEYINPUT88), .B(G120GAT), .ZN(n411) );
  XNOR2_X1 U473 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U474 ( .A(G113GAT), .B(n413), .ZN(n454) );
  XOR2_X1 U475 ( .A(KEYINPUT6), .B(G155GAT), .Z(n415) );
  XNOR2_X1 U476 ( .A(G1GAT), .B(G148GAT), .ZN(n414) );
  XNOR2_X1 U477 ( .A(n415), .B(n414), .ZN(n419) );
  XOR2_X1 U478 ( .A(G85GAT), .B(G162GAT), .Z(n417) );
  XNOR2_X1 U479 ( .A(G29GAT), .B(G127GAT), .ZN(n416) );
  XNOR2_X1 U480 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U481 ( .A(n419), .B(n418), .ZN(n430) );
  XOR2_X1 U482 ( .A(KEYINPUT97), .B(KEYINPUT98), .Z(n421) );
  XNOR2_X1 U483 ( .A(KEYINPUT4), .B(G57GAT), .ZN(n420) );
  XNOR2_X1 U484 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U485 ( .A(KEYINPUT5), .B(n422), .Z(n424) );
  NAND2_X1 U486 ( .A1(G225GAT), .A2(G233GAT), .ZN(n423) );
  XNOR2_X1 U487 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U488 ( .A(n425), .B(KEYINPUT1), .Z(n428) );
  XNOR2_X1 U489 ( .A(n426), .B(KEYINPUT96), .ZN(n427) );
  XNOR2_X1 U490 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U491 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U492 ( .A(n454), .B(n431), .Z(n525) );
  NAND2_X1 U493 ( .A1(n432), .A2(n525), .ZN(n433) );
  XNOR2_X1 U494 ( .A(n433), .B(KEYINPUT64), .ZN(n573) );
  NOR2_X1 U495 ( .A1(n476), .A2(n573), .ZN(n436) );
  INV_X1 U496 ( .A(n436), .ZN(n435) );
  INV_X1 U497 ( .A(KEYINPUT118), .ZN(n434) );
  NAND2_X1 U498 ( .A1(n435), .A2(n434), .ZN(n438) );
  NAND2_X1 U499 ( .A1(KEYINPUT118), .A2(n436), .ZN(n437) );
  NAND2_X1 U500 ( .A1(n438), .A2(n437), .ZN(n440) );
  INV_X1 U501 ( .A(KEYINPUT55), .ZN(n439) );
  XNOR2_X1 U502 ( .A(n440), .B(n439), .ZN(n456) );
  XOR2_X1 U503 ( .A(KEYINPUT20), .B(G190GAT), .Z(n442) );
  XNOR2_X1 U504 ( .A(G43GAT), .B(G99GAT), .ZN(n441) );
  XNOR2_X1 U505 ( .A(n442), .B(n441), .ZN(n445) );
  XOR2_X1 U506 ( .A(n446), .B(KEYINPUT91), .Z(n453) );
  XNOR2_X1 U507 ( .A(n447), .B(KEYINPUT89), .ZN(n451) );
  XOR2_X1 U508 ( .A(KEYINPUT90), .B(G183GAT), .Z(n449) );
  XNOR2_X1 U509 ( .A(G176GAT), .B(G71GAT), .ZN(n448) );
  XNOR2_X1 U510 ( .A(n449), .B(n448), .ZN(n450) );
  INV_X1 U511 ( .A(n542), .ZN(n493) );
  NAND2_X1 U512 ( .A1(n456), .A2(n493), .ZN(n567) );
  NOR2_X1 U513 ( .A1(n567), .A2(n556), .ZN(n458) );
  XNOR2_X1 U514 ( .A(G169GAT), .B(KEYINPUT119), .ZN(n457) );
  XNOR2_X1 U515 ( .A(n458), .B(n457), .ZN(G1348GAT) );
  XNOR2_X1 U516 ( .A(n559), .B(KEYINPUT108), .ZN(n544) );
  NOR2_X1 U517 ( .A1(n567), .A2(n544), .ZN(n462) );
  XNOR2_X1 U518 ( .A(KEYINPUT57), .B(KEYINPUT120), .ZN(n460) );
  XNOR2_X1 U519 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n459) );
  XNOR2_X1 U520 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U521 ( .A(n462), .B(n461), .ZN(G1349GAT) );
  NOR2_X1 U522 ( .A1(n565), .A2(n567), .ZN(n466) );
  XNOR2_X1 U523 ( .A(KEYINPUT58), .B(KEYINPUT122), .ZN(n464) );
  INV_X1 U524 ( .A(G190GAT), .ZN(n463) );
  XOR2_X1 U525 ( .A(KEYINPUT34), .B(KEYINPUT102), .Z(n488) );
  NAND2_X1 U526 ( .A1(n581), .A2(n574), .ZN(n467) );
  XNOR2_X1 U527 ( .A(n467), .B(KEYINPUT79), .ZN(n503) );
  NOR2_X1 U528 ( .A1(n586), .A2(n468), .ZN(n469) );
  XNOR2_X1 U529 ( .A(KEYINPUT16), .B(n469), .ZN(n484) );
  INV_X1 U530 ( .A(n525), .ZN(n486) );
  INV_X1 U531 ( .A(n490), .ZN(n529) );
  NOR2_X1 U532 ( .A1(n542), .A2(n529), .ZN(n470) );
  NOR2_X1 U533 ( .A1(n476), .A2(n470), .ZN(n471) );
  XOR2_X1 U534 ( .A(KEYINPUT25), .B(n471), .Z(n474) );
  NAND2_X1 U535 ( .A1(n542), .A2(n476), .ZN(n472) );
  XNOR2_X1 U536 ( .A(n472), .B(n295), .ZN(n554) );
  INV_X1 U537 ( .A(n554), .ZN(n572) );
  XOR2_X1 U538 ( .A(KEYINPUT27), .B(n490), .Z(n478) );
  NOR2_X1 U539 ( .A1(n572), .A2(n478), .ZN(n473) );
  NOR2_X1 U540 ( .A1(n474), .A2(n473), .ZN(n475) );
  NOR2_X1 U541 ( .A1(n486), .A2(n475), .ZN(n481) );
  XOR2_X1 U542 ( .A(n476), .B(KEYINPUT67), .Z(n477) );
  INV_X1 U543 ( .A(n540), .ZN(n498) );
  NOR2_X1 U544 ( .A1(n478), .A2(n525), .ZN(n538) );
  NAND2_X1 U545 ( .A1(n538), .A2(n542), .ZN(n479) );
  NOR2_X1 U546 ( .A1(n498), .A2(n479), .ZN(n480) );
  NOR2_X1 U547 ( .A1(n481), .A2(n480), .ZN(n483) );
  AND2_X1 U548 ( .A1(n484), .A2(n500), .ZN(n515) );
  NAND2_X1 U549 ( .A1(n503), .A2(n515), .ZN(n485) );
  XNOR2_X1 U550 ( .A(KEYINPUT101), .B(n485), .ZN(n497) );
  NAND2_X1 U551 ( .A1(n497), .A2(n486), .ZN(n487) );
  XNOR2_X1 U552 ( .A(n488), .B(n487), .ZN(n489) );
  XOR2_X1 U553 ( .A(G1GAT), .B(n489), .Z(G1324GAT) );
  XOR2_X1 U554 ( .A(G8GAT), .B(KEYINPUT103), .Z(n492) );
  NAND2_X1 U555 ( .A1(n497), .A2(n490), .ZN(n491) );
  XNOR2_X1 U556 ( .A(n492), .B(n491), .ZN(G1325GAT) );
  XOR2_X1 U557 ( .A(KEYINPUT104), .B(KEYINPUT35), .Z(n495) );
  NAND2_X1 U558 ( .A1(n497), .A2(n493), .ZN(n494) );
  XNOR2_X1 U559 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U560 ( .A(G15GAT), .B(n496), .ZN(G1326GAT) );
  NAND2_X1 U561 ( .A1(n498), .A2(n497), .ZN(n499) );
  XNOR2_X1 U562 ( .A(n499), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U563 ( .A1(n586), .A2(n500), .ZN(n501) );
  XOR2_X1 U564 ( .A(KEYINPUT37), .B(n502), .Z(n524) );
  NAND2_X1 U565 ( .A1(n503), .A2(n524), .ZN(n504) );
  XNOR2_X2 U566 ( .A(n504), .B(KEYINPUT38), .ZN(n512) );
  NOR2_X1 U567 ( .A1(n512), .A2(n525), .ZN(n506) );
  XNOR2_X1 U568 ( .A(KEYINPUT39), .B(KEYINPUT105), .ZN(n505) );
  XNOR2_X1 U569 ( .A(n506), .B(n505), .ZN(n507) );
  XOR2_X1 U570 ( .A(G29GAT), .B(n507), .Z(G1328GAT) );
  NOR2_X1 U571 ( .A1(n512), .A2(n529), .ZN(n508) );
  XOR2_X1 U572 ( .A(G36GAT), .B(n508), .Z(G1329GAT) );
  XNOR2_X1 U573 ( .A(KEYINPUT40), .B(KEYINPUT106), .ZN(n510) );
  XNOR2_X1 U574 ( .A(n510), .B(n509), .ZN(n511) );
  XOR2_X1 U575 ( .A(n511), .B(G43GAT), .Z(G1330GAT) );
  XNOR2_X1 U576 ( .A(G50GAT), .B(KEYINPUT107), .ZN(n514) );
  NOR2_X1 U577 ( .A1(n540), .A2(n512), .ZN(n513) );
  XNOR2_X1 U578 ( .A(n514), .B(n513), .ZN(G1331GAT) );
  NOR2_X1 U579 ( .A1(n574), .A2(n544), .ZN(n523) );
  NAND2_X1 U580 ( .A1(n515), .A2(n523), .ZN(n520) );
  NOR2_X1 U581 ( .A1(n525), .A2(n520), .ZN(n516) );
  XOR2_X1 U582 ( .A(G57GAT), .B(n516), .Z(n517) );
  XNOR2_X1 U583 ( .A(KEYINPUT42), .B(n517), .ZN(G1332GAT) );
  NOR2_X1 U584 ( .A1(n529), .A2(n520), .ZN(n518) );
  XOR2_X1 U585 ( .A(G64GAT), .B(n518), .Z(G1333GAT) );
  NOR2_X1 U586 ( .A1(n542), .A2(n520), .ZN(n519) );
  XOR2_X1 U587 ( .A(G71GAT), .B(n519), .Z(G1334GAT) );
  NOR2_X1 U588 ( .A1(n540), .A2(n520), .ZN(n522) );
  XNOR2_X1 U589 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n521) );
  XNOR2_X1 U590 ( .A(n522), .B(n521), .ZN(G1335GAT) );
  NAND2_X1 U591 ( .A1(n524), .A2(n523), .ZN(n534) );
  NOR2_X1 U592 ( .A1(n525), .A2(n534), .ZN(n527) );
  XNOR2_X1 U593 ( .A(KEYINPUT109), .B(KEYINPUT110), .ZN(n526) );
  XNOR2_X1 U594 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U595 ( .A(G85GAT), .B(n528), .ZN(G1336GAT) );
  NOR2_X1 U596 ( .A1(n529), .A2(n534), .ZN(n531) );
  XNOR2_X1 U597 ( .A(G92GAT), .B(KEYINPUT111), .ZN(n530) );
  XNOR2_X1 U598 ( .A(n531), .B(n530), .ZN(G1337GAT) );
  NOR2_X1 U599 ( .A1(n542), .A2(n534), .ZN(n532) );
  XOR2_X1 U600 ( .A(KEYINPUT112), .B(n532), .Z(n533) );
  XNOR2_X1 U601 ( .A(G99GAT), .B(n533), .ZN(G1338GAT) );
  NOR2_X1 U602 ( .A1(n540), .A2(n534), .ZN(n535) );
  XOR2_X1 U603 ( .A(KEYINPUT44), .B(n535), .Z(n536) );
  XNOR2_X1 U604 ( .A(G106GAT), .B(n536), .ZN(G1339GAT) );
  NAND2_X1 U605 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U606 ( .A(KEYINPUT115), .B(n539), .ZN(n555) );
  NAND2_X1 U607 ( .A1(n540), .A2(n555), .ZN(n541) );
  NOR2_X1 U608 ( .A1(n542), .A2(n541), .ZN(n547) );
  NAND2_X1 U609 ( .A1(n574), .A2(n547), .ZN(n543) );
  XNOR2_X1 U610 ( .A(G113GAT), .B(n543), .ZN(G1340GAT) );
  INV_X1 U611 ( .A(n547), .ZN(n550) );
  NOR2_X1 U612 ( .A1(n544), .A2(n550), .ZN(n546) );
  XNOR2_X1 U613 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n545) );
  XNOR2_X1 U614 ( .A(n546), .B(n545), .ZN(G1341GAT) );
  NAND2_X1 U615 ( .A1(n568), .A2(n547), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n548), .B(KEYINPUT50), .ZN(n549) );
  XNOR2_X1 U617 ( .A(G127GAT), .B(n549), .ZN(G1342GAT) );
  NOR2_X1 U618 ( .A1(n565), .A2(n550), .ZN(n552) );
  XNOR2_X1 U619 ( .A(KEYINPUT116), .B(KEYINPUT51), .ZN(n551) );
  XNOR2_X1 U620 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U621 ( .A(G134GAT), .B(n553), .ZN(G1343GAT) );
  NAND2_X1 U622 ( .A1(n555), .A2(n554), .ZN(n564) );
  NOR2_X1 U623 ( .A1(n556), .A2(n564), .ZN(n558) );
  XNOR2_X1 U624 ( .A(G141GAT), .B(KEYINPUT117), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n558), .B(n557), .ZN(G1344GAT) );
  NOR2_X1 U626 ( .A1(n559), .A2(n564), .ZN(n561) );
  XNOR2_X1 U627 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n560) );
  XNOR2_X1 U628 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U629 ( .A(G148GAT), .B(n562), .ZN(G1345GAT) );
  NOR2_X1 U630 ( .A1(n586), .A2(n564), .ZN(n563) );
  XOR2_X1 U631 ( .A(G155GAT), .B(n563), .Z(G1346GAT) );
  NOR2_X1 U632 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U633 ( .A(G162GAT), .B(n566), .Z(G1347GAT) );
  XOR2_X1 U634 ( .A(G183GAT), .B(KEYINPUT121), .Z(n571) );
  INV_X1 U635 ( .A(n567), .ZN(n569) );
  NAND2_X1 U636 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(G1350GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT124), .B(KEYINPUT60), .Z(n576) );
  NOR2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n580) );
  NAND2_X1 U640 ( .A1(n580), .A2(n574), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(n577) );
  XOR2_X1 U642 ( .A(n577), .B(KEYINPUT123), .Z(n579) );
  XNOR2_X1 U643 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1352GAT) );
  INV_X1 U645 ( .A(n580), .ZN(n589) );
  NOR2_X1 U646 ( .A1(n589), .A2(n581), .ZN(n585) );
  XOR2_X1 U647 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n583) );
  XNOR2_X1 U648 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n582) );
  XNOR2_X1 U649 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n585), .B(n584), .ZN(G1353GAT) );
  NOR2_X1 U651 ( .A1(n586), .A2(n589), .ZN(n588) );
  XNOR2_X1 U652 ( .A(G211GAT), .B(KEYINPUT127), .ZN(n587) );
  XNOR2_X1 U653 ( .A(n588), .B(n587), .ZN(G1354GAT) );
  NOR2_X1 U654 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U655 ( .A(KEYINPUT62), .B(n591), .Z(n592) );
  XNOR2_X1 U656 ( .A(G218GAT), .B(n592), .ZN(G1355GAT) );
endmodule

