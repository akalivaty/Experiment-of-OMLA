

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752;

  XNOR2_X1 U377 ( .A(n510), .B(n435), .ZN(n434) );
  NAND2_X1 U378 ( .A1(n387), .A2(n385), .ZN(n376) );
  XNOR2_X1 U379 ( .A(n376), .B(n486), .ZN(n600) );
  INV_X1 U380 ( .A(G953), .ZN(n743) );
  XNOR2_X2 U381 ( .A(n394), .B(n497), .ZN(n529) );
  XNOR2_X2 U382 ( .A(KEYINPUT64), .B(G143), .ZN(n451) );
  OR2_X1 U383 ( .A1(n597), .A2(n690), .ZN(n379) );
  NAND2_X1 U384 ( .A1(n640), .A2(n639), .ZN(n393) );
  XNOR2_X1 U385 ( .A(n581), .B(KEYINPUT40), .ZN(n750) );
  AND2_X1 U386 ( .A1(n381), .A2(n382), .ZN(n369) );
  NAND2_X1 U387 ( .A1(n358), .A2(n527), .ZN(n380) );
  XNOR2_X1 U388 ( .A(n468), .B(KEYINPUT105), .ZN(n702) );
  OR2_X1 U389 ( .A1(n534), .A2(n533), .ZN(n686) );
  XNOR2_X1 U390 ( .A(n372), .B(n623), .ZN(n625) );
  XNOR2_X1 U391 ( .A(n467), .B(n466), .ZN(n554) );
  XNOR2_X1 U392 ( .A(n644), .B(n643), .ZN(n645) );
  XNOR2_X1 U393 ( .A(KEYINPUT3), .B(KEYINPUT90), .ZN(n409) );
  XNOR2_X1 U394 ( .A(G101), .B(G119), .ZN(n410) );
  INV_X1 U395 ( .A(KEYINPUT107), .ZN(n378) );
  BUF_X1 U396 ( .A(n684), .Z(n355) );
  XNOR2_X1 U397 ( .A(n433), .B(KEYINPUT72), .ZN(n684) );
  BUF_X1 U398 ( .A(n616), .Z(n731) );
  INV_X1 U399 ( .A(n383), .ZN(n527) );
  XNOR2_X1 U400 ( .A(n379), .B(n378), .ZN(n383) );
  XNOR2_X2 U401 ( .A(n546), .B(KEYINPUT1), .ZN(n530) );
  XNOR2_X2 U402 ( .A(n516), .B(G469), .ZN(n546) );
  NOR2_X1 U403 ( .A1(n576), .A2(n391), .ZN(n390) );
  OR2_X1 U404 ( .A1(G237), .A2(G902), .ZN(n485) );
  XNOR2_X1 U405 ( .A(n412), .B(n411), .ZN(n620) );
  INV_X1 U406 ( .A(KEYINPUT48), .ZN(n411) );
  NAND2_X1 U407 ( .A1(n416), .A2(n413), .ZN(n412) );
  XNOR2_X1 U408 ( .A(n417), .B(n364), .ZN(n416) );
  XNOR2_X1 U409 ( .A(G137), .B(G134), .ZN(n498) );
  XNOR2_X1 U410 ( .A(n736), .B(n484), .ZN(n624) );
  XNOR2_X1 U411 ( .A(n415), .B(n414), .ZN(n413) );
  INV_X1 U412 ( .A(KEYINPUT69), .ZN(n414) );
  NOR2_X1 U413 ( .A1(n607), .A2(n671), .ZN(n415) );
  AND2_X1 U414 ( .A1(G953), .A2(G902), .ZN(n490) );
  OR2_X1 U415 ( .A1(n651), .A2(G902), .ZN(n516) );
  XNOR2_X1 U416 ( .A(KEYINPUT65), .B(KEYINPUT22), .ZN(n497) );
  NAND2_X1 U417 ( .A1(n620), .A2(n614), .ZN(n742) );
  XNOR2_X1 U418 ( .A(n404), .B(n408), .ZN(n507) );
  XNOR2_X1 U419 ( .A(n476), .B(G113), .ZN(n408) );
  XNOR2_X1 U420 ( .A(n410), .B(n409), .ZN(n404) );
  INV_X1 U421 ( .A(G116), .ZN(n476) );
  XNOR2_X1 U422 ( .A(KEYINPUT67), .B(KEYINPUT8), .ZN(n446) );
  XNOR2_X1 U423 ( .A(G116), .B(G107), .ZN(n442) );
  INV_X1 U424 ( .A(G128), .ZN(n450) );
  INV_X1 U425 ( .A(KEYINPUT95), .ZN(n435) );
  XNOR2_X1 U426 ( .A(G104), .B(G107), .ZN(n475) );
  NAND2_X1 U427 ( .A1(n356), .A2(n590), .ZN(n609) );
  NOR2_X1 U428 ( .A1(n703), .A2(n702), .ZN(n582) );
  XNOR2_X1 U429 ( .A(n579), .B(n580), .ZN(n423) );
  XNOR2_X1 U430 ( .A(n530), .B(KEYINPUT87), .ZN(n597) );
  NAND2_X1 U431 ( .A1(n386), .A2(n576), .ZN(n385) );
  AND2_X1 U432 ( .A1(n388), .A2(n363), .ZN(n387) );
  XNOR2_X1 U433 ( .A(n609), .B(KEYINPUT114), .ZN(n594) );
  XNOR2_X1 U434 ( .A(n425), .B(n424), .ZN(n602) );
  INV_X1 U435 ( .A(KEYINPUT74), .ZN(n424) );
  NAND2_X1 U436 ( .A1(n428), .A2(n426), .ZN(n425) );
  XNOR2_X1 U437 ( .A(n567), .B(n429), .ZN(n428) );
  OR2_X1 U438 ( .A1(n631), .A2(G902), .ZN(n396) );
  XNOR2_X1 U439 ( .A(n453), .B(n452), .ZN(n553) );
  XNOR2_X1 U440 ( .A(n525), .B(KEYINPUT25), .ZN(n526) );
  BUF_X1 U441 ( .A(n529), .Z(n559) );
  BUF_X1 U442 ( .A(n530), .Z(n401) );
  XNOR2_X1 U443 ( .A(n422), .B(n421), .ZN(n420) );
  INV_X1 U444 ( .A(KEYINPUT81), .ZN(n421) );
  NAND2_X1 U445 ( .A1(n682), .A2(n683), .ZN(n422) );
  INV_X1 U446 ( .A(KEYINPUT34), .ZN(n538) );
  NOR2_X1 U447 ( .A1(G953), .A2(G237), .ZN(n503) );
  XOR2_X1 U448 ( .A(G146), .B(G125), .Z(n480) );
  NAND2_X1 U449 ( .A1(G234), .A2(G237), .ZN(n487) );
  AND2_X1 U450 ( .A1(n540), .A2(n554), .ZN(n468) );
  XNOR2_X1 U451 ( .A(n578), .B(KEYINPUT38), .ZN(n399) );
  INV_X1 U452 ( .A(KEYINPUT71), .ZN(n578) );
  NAND2_X1 U453 ( .A1(n576), .A2(n391), .ZN(n389) );
  XNOR2_X1 U454 ( .A(G902), .B(KEYINPUT89), .ZN(n470) );
  INV_X1 U455 ( .A(KEYINPUT110), .ZN(n429) );
  AND2_X1 U456 ( .A1(n571), .A2(n427), .ZN(n426) );
  INV_X1 U457 ( .A(n583), .ZN(n427) );
  INV_X1 U458 ( .A(G902), .ZN(n465) );
  XOR2_X1 U459 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n520) );
  XNOR2_X1 U460 ( .A(n480), .B(n455), .ZN(n523) );
  XNOR2_X1 U461 ( .A(n454), .B(KEYINPUT10), .ZN(n455) );
  INV_X1 U462 ( .A(G140), .ZN(n454) );
  XNOR2_X1 U463 ( .A(G143), .B(G122), .ZN(n458) );
  XOR2_X1 U464 ( .A(KEYINPUT12), .B(G104), .Z(n459) );
  INV_X1 U465 ( .A(G113), .ZN(n462) );
  XOR2_X1 U466 ( .A(KEYINPUT11), .B(KEYINPUT99), .Z(n457) );
  NOR2_X1 U467 ( .A1(n731), .A2(KEYINPUT2), .ZN(n677) );
  AND2_X1 U468 ( .A1(n681), .A2(n362), .ZN(n682) );
  INV_X1 U469 ( .A(KEYINPUT19), .ZN(n486) );
  XNOR2_X1 U470 ( .A(n631), .B(n630), .ZN(n632) );
  XNOR2_X1 U471 ( .A(n507), .B(G122), .ZN(n403) );
  XNOR2_X1 U472 ( .A(n449), .B(n398), .ZN(n722) );
  BUF_X1 U473 ( .A(n649), .Z(n726) );
  XNOR2_X1 U474 ( .A(n434), .B(n359), .ZN(n651) );
  XNOR2_X1 U475 ( .A(G146), .B(G140), .ZN(n512) );
  BUF_X1 U476 ( .A(n624), .Z(n372) );
  XNOR2_X1 U477 ( .A(n589), .B(n370), .ZN(n752) );
  XNOR2_X1 U478 ( .A(KEYINPUT42), .B(KEYINPUT113), .ZN(n370) );
  NAND2_X1 U479 ( .A1(n423), .A2(n590), .ZN(n581) );
  XNOR2_X1 U480 ( .A(KEYINPUT36), .B(KEYINPUT115), .ZN(n595) );
  XNOR2_X1 U481 ( .A(KEYINPUT112), .B(n605), .ZN(n751) );
  NOR2_X1 U482 ( .A1(n401), .A2(n557), .ZN(n558) );
  INV_X1 U483 ( .A(KEYINPUT53), .ZN(n418) );
  NAND2_X1 U484 ( .A1(n420), .A2(n721), .ZN(n419) );
  INV_X1 U485 ( .A(G122), .ZN(n438) );
  XOR2_X1 U486 ( .A(n593), .B(KEYINPUT109), .Z(n356) );
  NOR2_X1 U487 ( .A1(n540), .A2(n554), .ZN(n357) );
  AND2_X1 U488 ( .A1(n529), .A2(n436), .ZN(n358) );
  XOR2_X1 U489 ( .A(n515), .B(n514), .Z(n359) );
  AND2_X1 U490 ( .A1(G221), .A2(n517), .ZN(n360) );
  XOR2_X1 U491 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n361) );
  NAND2_X1 U492 ( .A1(n731), .A2(n621), .ZN(n362) );
  AND2_X1 U493 ( .A1(n389), .A2(n699), .ZN(n363) );
  XOR2_X1 U494 ( .A(KEYINPUT46), .B(KEYINPUT82), .Z(n364) );
  XNOR2_X1 U495 ( .A(n470), .B(n469), .ZN(n615) );
  INV_X1 U496 ( .A(n615), .ZN(n391) );
  INV_X1 U497 ( .A(n699), .ZN(n392) );
  XNOR2_X1 U498 ( .A(n403), .B(n477), .ZN(n736) );
  OR2_X1 U499 ( .A1(n615), .A2(n678), .ZN(n365) );
  NAND2_X1 U500 ( .A1(n543), .A2(KEYINPUT84), .ZN(n368) );
  XNOR2_X2 U501 ( .A(n542), .B(KEYINPUT35), .ZN(n543) );
  NAND2_X1 U502 ( .A1(n366), .A2(n544), .ZN(n432) );
  NAND2_X1 U503 ( .A1(n368), .A2(n367), .ZN(n366) );
  AND2_X2 U504 ( .A1(n402), .A2(KEYINPUT44), .ZN(n367) );
  XNOR2_X2 U505 ( .A(n393), .B(KEYINPUT85), .ZN(n402) );
  XNOR2_X1 U506 ( .A(n374), .B(n407), .ZN(n373) );
  XNOR2_X1 U507 ( .A(n371), .B(KEYINPUT45), .ZN(n616) );
  NAND2_X1 U508 ( .A1(n616), .A2(n391), .ZN(n374) );
  NAND2_X1 U509 ( .A1(n369), .A2(n380), .ZN(n640) );
  INV_X1 U510 ( .A(n742), .ZN(n406) );
  NAND2_X1 U511 ( .A1(n432), .A2(n566), .ZN(n371) );
  NAND2_X1 U512 ( .A1(n624), .A2(n390), .ZN(n388) );
  XNOR2_X1 U513 ( .A(n612), .B(n399), .ZN(n700) );
  NAND2_X1 U514 ( .A1(n372), .A2(n615), .ZN(n577) );
  AND2_X2 U515 ( .A1(n405), .A2(n362), .ZN(n649) );
  NAND2_X1 U516 ( .A1(n373), .A2(n406), .ZN(n375) );
  NAND2_X1 U517 ( .A1(n375), .A2(n365), .ZN(n405) );
  NOR2_X1 U518 ( .A1(n594), .A2(n376), .ZN(n596) );
  XNOR2_X2 U519 ( .A(n377), .B(n482), .ZN(n501) );
  XNOR2_X1 U520 ( .A(n377), .B(n448), .ZN(n398) );
  XNOR2_X2 U521 ( .A(n451), .B(n450), .ZN(n377) );
  NAND2_X1 U522 ( .A1(n384), .A2(n528), .ZN(n381) );
  NAND2_X1 U523 ( .A1(n383), .A2(n528), .ZN(n382) );
  NAND2_X1 U524 ( .A1(n529), .A2(n592), .ZN(n384) );
  INV_X1 U525 ( .A(n624), .ZN(n386) );
  NAND2_X1 U526 ( .A1(n549), .A2(n496), .ZN(n394) );
  XNOR2_X1 U527 ( .A(n395), .B(n461), .ZN(n464) );
  XNOR2_X1 U528 ( .A(n460), .B(n463), .ZN(n395) );
  XNOR2_X2 U529 ( .A(n396), .B(G472), .ZN(n568) );
  XNOR2_X1 U530 ( .A(n397), .B(n400), .ZN(n483) );
  XNOR2_X1 U531 ( .A(n479), .B(n481), .ZN(n397) );
  XNOR2_X1 U532 ( .A(n419), .B(n418), .ZN(G75) );
  INV_X1 U533 ( .A(n480), .ZN(n400) );
  NAND2_X1 U534 ( .A1(n649), .A2(G475), .ZN(n646) );
  NOR2_X2 U535 ( .A1(n634), .A2(n730), .ZN(n636) );
  NOR2_X2 U536 ( .A1(n628), .A2(n730), .ZN(n629) );
  NOR2_X2 U537 ( .A1(n647), .A2(n730), .ZN(n648) );
  NAND2_X1 U538 ( .A1(n402), .A2(n545), .ZN(n562) );
  INV_X1 U539 ( .A(KEYINPUT80), .ZN(n407) );
  NAND2_X1 U540 ( .A1(n750), .A2(n752), .ZN(n417) );
  NAND2_X1 U541 ( .A1(n423), .A2(n608), .ZN(n674) );
  XNOR2_X2 U542 ( .A(n526), .B(n430), .ZN(n690) );
  NOR2_X1 U543 ( .A1(n727), .A2(G902), .ZN(n430) );
  XNOR2_X1 U544 ( .A(n431), .B(n741), .ZN(n727) );
  XNOR2_X1 U545 ( .A(n522), .B(n360), .ZN(n431) );
  NOR2_X2 U546 ( .A1(n684), .A2(n592), .ZN(n537) );
  NAND2_X1 U547 ( .A1(n439), .A2(n530), .ZN(n433) );
  XNOR2_X1 U548 ( .A(n434), .B(n741), .ZN(n745) );
  AND2_X1 U549 ( .A1(n592), .A2(n437), .ZN(n436) );
  INV_X1 U550 ( .A(n528), .ZN(n437) );
  NAND2_X1 U551 ( .A1(n543), .A2(n563), .ZN(n564) );
  XNOR2_X1 U552 ( .A(n543), .B(n438), .ZN(G24) );
  INV_X1 U553 ( .A(n401), .ZN(n687) );
  INV_X1 U554 ( .A(n686), .ZN(n439) );
  XNOR2_X1 U555 ( .A(n501), .B(n483), .ZN(n484) );
  INV_X1 U556 ( .A(KEYINPUT4), .ZN(n482) );
  INV_X1 U557 ( .A(KEYINPUT79), .ZN(n679) );
  XNOR2_X1 U558 ( .A(n521), .B(n520), .ZN(n522) );
  BUF_X1 U559 ( .A(n546), .Z(n587) );
  XNOR2_X1 U560 ( .A(n596), .B(n595), .ZN(n598) );
  AND2_X1 U561 ( .A1(n720), .A2(n743), .ZN(n721) );
  INV_X1 U562 ( .A(KEYINPUT63), .ZN(n635) );
  XOR2_X1 U563 ( .A(KEYINPUT100), .B(KEYINPUT7), .Z(n441) );
  XNOR2_X1 U564 ( .A(G134), .B(G122), .ZN(n440) );
  XNOR2_X1 U565 ( .A(n441), .B(n440), .ZN(n445) );
  XOR2_X1 U566 ( .A(KEYINPUT9), .B(KEYINPUT101), .Z(n443) );
  XNOR2_X1 U567 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U568 ( .A(n445), .B(n444), .Z(n449) );
  NAND2_X1 U569 ( .A1(n743), .A2(G234), .ZN(n447) );
  XNOR2_X1 U570 ( .A(n447), .B(n446), .ZN(n517) );
  NAND2_X1 U571 ( .A1(G217), .A2(n517), .ZN(n448) );
  NAND2_X1 U572 ( .A1(n722), .A2(n465), .ZN(n453) );
  XNOR2_X1 U573 ( .A(KEYINPUT102), .B(G478), .ZN(n452) );
  INV_X1 U574 ( .A(n553), .ZN(n540) );
  NAND2_X1 U575 ( .A1(G214), .A2(n503), .ZN(n456) );
  XNOR2_X1 U576 ( .A(n457), .B(n456), .ZN(n461) );
  XNOR2_X1 U577 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X2 U578 ( .A(KEYINPUT68), .B(G131), .ZN(n499) );
  XNOR2_X1 U579 ( .A(n499), .B(n462), .ZN(n463) );
  XNOR2_X1 U580 ( .A(n523), .B(n464), .ZN(n644) );
  NAND2_X1 U581 ( .A1(n644), .A2(n465), .ZN(n467) );
  XNOR2_X1 U582 ( .A(KEYINPUT13), .B(G475), .ZN(n466) );
  XOR2_X1 U583 ( .A(KEYINPUT96), .B(KEYINPUT21), .Z(n473) );
  INV_X1 U584 ( .A(KEYINPUT15), .ZN(n469) );
  NAND2_X1 U585 ( .A1(n615), .A2(G234), .ZN(n471) );
  XNOR2_X1 U586 ( .A(n471), .B(KEYINPUT20), .ZN(n524) );
  NAND2_X1 U587 ( .A1(n524), .A2(G221), .ZN(n472) );
  XNOR2_X1 U588 ( .A(n473), .B(n472), .ZN(n689) );
  XNOR2_X1 U589 ( .A(n689), .B(KEYINPUT97), .ZN(n534) );
  NOR2_X1 U590 ( .A1(n702), .A2(n534), .ZN(n474) );
  XNOR2_X1 U591 ( .A(KEYINPUT106), .B(n474), .ZN(n496) );
  XNOR2_X1 U592 ( .A(n475), .B(G110), .ZN(n515) );
  XOR2_X1 U593 ( .A(n515), .B(KEYINPUT16), .Z(n477) );
  XNOR2_X1 U594 ( .A(KEYINPUT91), .B(KEYINPUT75), .ZN(n478) );
  XNOR2_X1 U595 ( .A(n361), .B(n478), .ZN(n479) );
  NAND2_X1 U596 ( .A1(G224), .A2(n743), .ZN(n481) );
  NAND2_X1 U597 ( .A1(G210), .A2(n485), .ZN(n576) );
  NAND2_X1 U598 ( .A1(G214), .A2(n485), .ZN(n699) );
  XNOR2_X1 U599 ( .A(n487), .B(KEYINPUT14), .ZN(n491) );
  NAND2_X1 U600 ( .A1(n491), .A2(G952), .ZN(n488) );
  XNOR2_X1 U601 ( .A(n488), .B(KEYINPUT92), .ZN(n715) );
  NOR2_X1 U602 ( .A1(G953), .A2(n715), .ZN(n489) );
  XOR2_X1 U603 ( .A(KEYINPUT93), .B(n489), .Z(n575) );
  NAND2_X1 U604 ( .A1(n491), .A2(n490), .ZN(n572) );
  NOR2_X1 U605 ( .A1(G898), .A2(n572), .ZN(n492) );
  NOR2_X1 U606 ( .A1(n575), .A2(n492), .ZN(n493) );
  XNOR2_X1 U607 ( .A(n493), .B(KEYINPUT94), .ZN(n494) );
  NOR2_X2 U608 ( .A1(n600), .A2(n494), .ZN(n495) );
  XNOR2_X2 U609 ( .A(n495), .B(KEYINPUT0), .ZN(n549) );
  XNOR2_X1 U610 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X2 U611 ( .A(n501), .B(n500), .ZN(n510) );
  XNOR2_X1 U612 ( .A(G146), .B(KEYINPUT5), .ZN(n502) );
  XNOR2_X1 U613 ( .A(n502), .B(KEYINPUT73), .ZN(n505) );
  NAND2_X1 U614 ( .A1(n503), .A2(G210), .ZN(n504) );
  XNOR2_X1 U615 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U616 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U617 ( .A(n510), .B(n508), .ZN(n631) );
  XNOR2_X1 U618 ( .A(KEYINPUT104), .B(KEYINPUT6), .ZN(n509) );
  XNOR2_X1 U619 ( .A(n568), .B(n509), .ZN(n592) );
  NAND2_X1 U620 ( .A1(n743), .A2(G227), .ZN(n511) );
  XNOR2_X1 U621 ( .A(n511), .B(G101), .ZN(n513) );
  XNOR2_X1 U622 ( .A(n513), .B(n512), .ZN(n514) );
  XOR2_X1 U623 ( .A(G110), .B(G128), .Z(n519) );
  XNOR2_X1 U624 ( .A(G119), .B(G137), .ZN(n518) );
  XNOR2_X1 U625 ( .A(n519), .B(n518), .ZN(n521) );
  INV_X1 U626 ( .A(n523), .ZN(n741) );
  NAND2_X1 U627 ( .A1(n524), .A2(G217), .ZN(n525) );
  XNOR2_X1 U628 ( .A(KEYINPUT76), .B(KEYINPUT32), .ZN(n528) );
  NOR2_X1 U629 ( .A1(n568), .A2(n690), .ZN(n531) );
  AND2_X1 U630 ( .A1(n531), .A2(n687), .ZN(n532) );
  NAND2_X1 U631 ( .A1(n559), .A2(n532), .ZN(n639) );
  INV_X1 U632 ( .A(n690), .ZN(n533) );
  INV_X1 U633 ( .A(KEYINPUT70), .ZN(n535) );
  XNOR2_X1 U634 ( .A(n535), .B(KEYINPUT33), .ZN(n536) );
  XNOR2_X1 U635 ( .A(n537), .B(n536), .ZN(n708) );
  NAND2_X1 U636 ( .A1(n708), .A2(n549), .ZN(n539) );
  XNOR2_X1 U637 ( .A(n539), .B(n538), .ZN(n541) );
  NAND2_X1 U638 ( .A1(n541), .A2(n357), .ZN(n542) );
  INV_X1 U639 ( .A(KEYINPUT44), .ZN(n545) );
  NAND2_X1 U640 ( .A1(n545), .A2(KEYINPUT84), .ZN(n544) );
  INV_X1 U641 ( .A(n549), .ZN(n547) );
  NAND2_X1 U642 ( .A1(n587), .A2(n439), .ZN(n567) );
  NOR2_X1 U643 ( .A1(n547), .A2(n567), .ZN(n548) );
  INV_X1 U644 ( .A(n568), .ZN(n585) );
  NAND2_X1 U645 ( .A1(n548), .A2(n585), .ZN(n656) );
  NAND2_X1 U646 ( .A1(n549), .A2(n568), .ZN(n550) );
  NOR2_X1 U647 ( .A1(n550), .A2(n355), .ZN(n552) );
  XNOR2_X1 U648 ( .A(KEYINPUT98), .B(KEYINPUT31), .ZN(n551) );
  XNOR2_X1 U649 ( .A(n552), .B(n551), .ZN(n669) );
  NAND2_X1 U650 ( .A1(n656), .A2(n669), .ZN(n556) );
  NOR2_X1 U651 ( .A1(n554), .A2(n553), .ZN(n590) );
  NAND2_X1 U652 ( .A1(n554), .A2(n553), .ZN(n668) );
  XNOR2_X1 U653 ( .A(KEYINPUT103), .B(n668), .ZN(n608) );
  NOR2_X1 U654 ( .A1(n590), .A2(n608), .ZN(n704) );
  INV_X1 U655 ( .A(n704), .ZN(n555) );
  NAND2_X1 U656 ( .A1(n556), .A2(n555), .ZN(n560) );
  NAND2_X1 U657 ( .A1(n592), .A2(n690), .ZN(n557) );
  NAND2_X1 U658 ( .A1(n559), .A2(n558), .ZN(n638) );
  AND2_X1 U659 ( .A1(n560), .A2(n638), .ZN(n563) );
  AND2_X1 U660 ( .A1(KEYINPUT84), .A2(n563), .ZN(n561) );
  NAND2_X1 U661 ( .A1(n562), .A2(n561), .ZN(n565) );
  NAND2_X1 U662 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U663 ( .A(KEYINPUT83), .B(KEYINPUT39), .Z(n580) );
  NAND2_X1 U664 ( .A1(n699), .A2(n568), .ZN(n569) );
  XNOR2_X1 U665 ( .A(n569), .B(KEYINPUT30), .ZN(n570) );
  XNOR2_X1 U666 ( .A(n570), .B(KEYINPUT111), .ZN(n571) );
  XNOR2_X1 U667 ( .A(KEYINPUT108), .B(n572), .ZN(n573) );
  NOR2_X1 U668 ( .A1(G900), .A2(n573), .ZN(n574) );
  NOR2_X1 U669 ( .A1(n575), .A2(n574), .ZN(n583) );
  XNOR2_X1 U670 ( .A(n577), .B(n576), .ZN(n612) );
  NAND2_X1 U671 ( .A1(n602), .A2(n700), .ZN(n579) );
  NAND2_X1 U672 ( .A1(n700), .A2(n699), .ZN(n703) );
  XNOR2_X1 U673 ( .A(n582), .B(KEYINPUT41), .ZN(n717) );
  NOR2_X1 U674 ( .A1(n583), .A2(n690), .ZN(n584) );
  NAND2_X1 U675 ( .A1(n689), .A2(n584), .ZN(n591) );
  NOR2_X1 U676 ( .A1(n591), .A2(n585), .ZN(n586) );
  XNOR2_X1 U677 ( .A(KEYINPUT28), .B(n586), .ZN(n588) );
  NAND2_X1 U678 ( .A1(n588), .A2(n587), .ZN(n599) );
  NOR2_X1 U679 ( .A1(n717), .A2(n599), .ZN(n589) );
  INV_X1 U680 ( .A(n590), .ZN(n666) );
  NOR2_X1 U681 ( .A1(n592), .A2(n591), .ZN(n593) );
  NOR2_X1 U682 ( .A1(n598), .A2(n597), .ZN(n671) );
  OR2_X1 U683 ( .A1(n600), .A2(n599), .ZN(n664) );
  NOR2_X1 U684 ( .A1(n704), .A2(n664), .ZN(n601) );
  XNOR2_X1 U685 ( .A(KEYINPUT47), .B(n601), .ZN(n606) );
  INV_X1 U686 ( .A(n612), .ZN(n603) );
  AND2_X1 U687 ( .A1(n603), .A2(n602), .ZN(n604) );
  NAND2_X1 U688 ( .A1(n357), .A2(n604), .ZN(n605) );
  NAND2_X1 U689 ( .A1(n606), .A2(n751), .ZN(n607) );
  NOR2_X1 U690 ( .A1(n609), .A2(n392), .ZN(n610) );
  NAND2_X1 U691 ( .A1(n610), .A2(n687), .ZN(n611) );
  XNOR2_X1 U692 ( .A(n611), .B(KEYINPUT43), .ZN(n613) );
  NAND2_X1 U693 ( .A1(n613), .A2(n612), .ZN(n676) );
  AND2_X1 U694 ( .A1(n674), .A2(n676), .ZN(n614) );
  INV_X1 U695 ( .A(KEYINPUT2), .ZN(n678) );
  NAND2_X1 U696 ( .A1(KEYINPUT2), .A2(n674), .ZN(n617) );
  XNOR2_X1 U697 ( .A(KEYINPUT77), .B(n617), .ZN(n618) );
  AND2_X1 U698 ( .A1(n618), .A2(n676), .ZN(n619) );
  AND2_X1 U699 ( .A1(n620), .A2(n619), .ZN(n621) );
  NAND2_X1 U700 ( .A1(n649), .A2(G210), .ZN(n626) );
  XNOR2_X1 U701 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n622) );
  XOR2_X1 U702 ( .A(n622), .B(KEYINPUT123), .Z(n623) );
  XNOR2_X1 U703 ( .A(n626), .B(n625), .ZN(n628) );
  INV_X1 U704 ( .A(G952), .ZN(n627) );
  AND2_X1 U705 ( .A1(n627), .A2(G953), .ZN(n730) );
  XNOR2_X1 U706 ( .A(n629), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U707 ( .A1(n649), .A2(G472), .ZN(n633) );
  XNOR2_X1 U708 ( .A(KEYINPUT86), .B(KEYINPUT62), .ZN(n630) );
  XNOR2_X1 U709 ( .A(n633), .B(n632), .ZN(n634) );
  XNOR2_X1 U710 ( .A(n636), .B(n635), .ZN(G57) );
  XNOR2_X1 U711 ( .A(G101), .B(KEYINPUT116), .ZN(n637) );
  XNOR2_X1 U712 ( .A(n638), .B(n637), .ZN(G3) );
  XNOR2_X1 U713 ( .A(n639), .B(G110), .ZN(G12) );
  XNOR2_X1 U714 ( .A(n640), .B(G119), .ZN(G21) );
  XNOR2_X1 U715 ( .A(KEYINPUT88), .B(KEYINPUT124), .ZN(n642) );
  XNOR2_X1 U716 ( .A(KEYINPUT59), .B(KEYINPUT66), .ZN(n641) );
  XNOR2_X1 U717 ( .A(n642), .B(n641), .ZN(n643) );
  XNOR2_X1 U718 ( .A(n646), .B(n645), .ZN(n647) );
  XNOR2_X1 U719 ( .A(n648), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U720 ( .A1(n726), .A2(G469), .ZN(n653) );
  XOR2_X1 U721 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n650) );
  XNOR2_X1 U722 ( .A(n651), .B(n650), .ZN(n652) );
  XNOR2_X1 U723 ( .A(n653), .B(n652), .ZN(n654) );
  NOR2_X1 U724 ( .A1(n654), .A2(n730), .ZN(G54) );
  NOR2_X1 U725 ( .A1(n666), .A2(n656), .ZN(n655) );
  XOR2_X1 U726 ( .A(G104), .B(n655), .Z(G6) );
  NOR2_X1 U727 ( .A1(n668), .A2(n656), .ZN(n661) );
  XOR2_X1 U728 ( .A(KEYINPUT27), .B(KEYINPUT118), .Z(n658) );
  XNOR2_X1 U729 ( .A(G107), .B(KEYINPUT117), .ZN(n657) );
  XNOR2_X1 U730 ( .A(n658), .B(n657), .ZN(n659) );
  XNOR2_X1 U731 ( .A(KEYINPUT26), .B(n659), .ZN(n660) );
  XNOR2_X1 U732 ( .A(n661), .B(n660), .ZN(G9) );
  NOR2_X1 U733 ( .A1(n668), .A2(n664), .ZN(n663) );
  XNOR2_X1 U734 ( .A(G128), .B(KEYINPUT29), .ZN(n662) );
  XNOR2_X1 U735 ( .A(n663), .B(n662), .ZN(G30) );
  NOR2_X1 U736 ( .A1(n666), .A2(n664), .ZN(n665) );
  XOR2_X1 U737 ( .A(G146), .B(n665), .Z(G48) );
  NOR2_X1 U738 ( .A1(n669), .A2(n666), .ZN(n667) );
  XOR2_X1 U739 ( .A(G113), .B(n667), .Z(G15) );
  NOR2_X1 U740 ( .A1(n669), .A2(n668), .ZN(n670) );
  XOR2_X1 U741 ( .A(G116), .B(n670), .Z(G18) );
  XOR2_X1 U742 ( .A(KEYINPUT37), .B(KEYINPUT119), .Z(n673) );
  XNOR2_X1 U743 ( .A(n671), .B(G125), .ZN(n672) );
  XNOR2_X1 U744 ( .A(n673), .B(n672), .ZN(G27) );
  XNOR2_X1 U745 ( .A(G134), .B(KEYINPUT120), .ZN(n675) );
  XNOR2_X1 U746 ( .A(n675), .B(n674), .ZN(G36) );
  XNOR2_X1 U747 ( .A(G140), .B(n676), .ZN(G42) );
  XOR2_X1 U748 ( .A(KEYINPUT78), .B(n677), .Z(n683) );
  NAND2_X1 U749 ( .A1(n678), .A2(n742), .ZN(n680) );
  XNOR2_X1 U750 ( .A(n680), .B(n679), .ZN(n681) );
  INV_X1 U751 ( .A(n355), .ZN(n685) );
  NAND2_X1 U752 ( .A1(n685), .A2(n568), .ZN(n696) );
  NAND2_X1 U753 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U754 ( .A(n688), .B(KEYINPUT50), .ZN(n694) );
  NOR2_X1 U755 ( .A1(n690), .A2(n689), .ZN(n691) );
  XOR2_X1 U756 ( .A(KEYINPUT49), .B(n691), .Z(n692) );
  NOR2_X1 U757 ( .A1(n568), .A2(n692), .ZN(n693) );
  NAND2_X1 U758 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U759 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U760 ( .A(KEYINPUT51), .B(n697), .ZN(n698) );
  NOR2_X1 U761 ( .A1(n698), .A2(n717), .ZN(n711) );
  NOR2_X1 U762 ( .A1(n700), .A2(n699), .ZN(n701) );
  NOR2_X1 U763 ( .A1(n702), .A2(n701), .ZN(n707) );
  NOR2_X1 U764 ( .A1(n704), .A2(n703), .ZN(n705) );
  XOR2_X1 U765 ( .A(KEYINPUT121), .B(n705), .Z(n706) );
  NOR2_X1 U766 ( .A1(n707), .A2(n706), .ZN(n709) );
  INV_X1 U767 ( .A(n708), .ZN(n716) );
  NOR2_X1 U768 ( .A1(n709), .A2(n716), .ZN(n710) );
  NOR2_X1 U769 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U770 ( .A(n712), .B(KEYINPUT122), .ZN(n713) );
  XNOR2_X1 U771 ( .A(KEYINPUT52), .B(n713), .ZN(n714) );
  NOR2_X1 U772 ( .A1(n715), .A2(n714), .ZN(n719) );
  NOR2_X1 U773 ( .A1(n717), .A2(n716), .ZN(n718) );
  NOR2_X1 U774 ( .A1(n719), .A2(n718), .ZN(n720) );
  NAND2_X1 U775 ( .A1(n726), .A2(G478), .ZN(n724) );
  XNOR2_X1 U776 ( .A(n722), .B(KEYINPUT125), .ZN(n723) );
  XNOR2_X1 U777 ( .A(n724), .B(n723), .ZN(n725) );
  NOR2_X1 U778 ( .A1(n730), .A2(n725), .ZN(G63) );
  NAND2_X1 U779 ( .A1(n726), .A2(G217), .ZN(n728) );
  XNOR2_X1 U780 ( .A(n728), .B(n727), .ZN(n729) );
  NOR2_X1 U781 ( .A1(n730), .A2(n729), .ZN(G66) );
  NAND2_X1 U782 ( .A1(n731), .A2(n743), .ZN(n735) );
  NAND2_X1 U783 ( .A1(G953), .A2(G224), .ZN(n732) );
  XNOR2_X1 U784 ( .A(KEYINPUT61), .B(n732), .ZN(n733) );
  NAND2_X1 U785 ( .A1(n733), .A2(G898), .ZN(n734) );
  NAND2_X1 U786 ( .A1(n735), .A2(n734), .ZN(n739) );
  NOR2_X1 U787 ( .A1(G898), .A2(n743), .ZN(n737) );
  NOR2_X1 U788 ( .A1(n736), .A2(n737), .ZN(n738) );
  XNOR2_X1 U789 ( .A(n739), .B(n738), .ZN(n740) );
  XNOR2_X1 U790 ( .A(KEYINPUT126), .B(n740), .ZN(G69) );
  XNOR2_X1 U791 ( .A(n742), .B(n745), .ZN(n744) );
  NAND2_X1 U792 ( .A1(n744), .A2(n743), .ZN(n749) );
  XNOR2_X1 U793 ( .A(n745), .B(G227), .ZN(n746) );
  NAND2_X1 U794 ( .A1(n746), .A2(G900), .ZN(n747) );
  NAND2_X1 U795 ( .A1(n747), .A2(G953), .ZN(n748) );
  NAND2_X1 U796 ( .A1(n749), .A2(n748), .ZN(G72) );
  XNOR2_X1 U797 ( .A(G131), .B(n750), .ZN(G33) );
  XNOR2_X1 U798 ( .A(G143), .B(n751), .ZN(G45) );
  XNOR2_X1 U799 ( .A(n752), .B(G137), .ZN(G39) );
endmodule

