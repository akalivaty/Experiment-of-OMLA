

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744;

  XNOR2_X1 U371 ( .A(n390), .B(n389), .ZN(n602) );
  XNOR2_X1 U372 ( .A(n484), .B(n485), .ZN(n713) );
  XNOR2_X2 U373 ( .A(n392), .B(KEYINPUT19), .ZN(n576) );
  NAND2_X2 U374 ( .A1(n550), .A2(n658), .ZN(n392) );
  NOR2_X2 U375 ( .A1(n562), .A2(n561), .ZN(n563) );
  INV_X2 U376 ( .A(G143), .ZN(n370) );
  NOR2_X2 U377 ( .A1(n552), .A2(n582), .ZN(n632) );
  XNOR2_X2 U378 ( .A(n502), .B(n513), .ZN(n725) );
  INV_X2 U379 ( .A(G953), .ZN(n729) );
  AND2_X1 U380 ( .A1(n611), .A2(n743), .ZN(n612) );
  XNOR2_X1 U381 ( .A(n483), .B(KEYINPUT77), .ZN(n551) );
  XNOR2_X2 U382 ( .A(n510), .B(n441), .ZN(n723) );
  INV_X1 U383 ( .A(KEYINPUT91), .ZN(n389) );
  INV_X1 U384 ( .A(KEYINPUT66), .ZN(n391) );
  NOR2_X1 U385 ( .A1(n615), .A2(n614), .ZN(n616) );
  NOR2_X1 U386 ( .A1(n564), .A2(n542), .ZN(n519) );
  XNOR2_X1 U387 ( .A(n495), .B(n494), .ZN(n564) );
  AND2_X1 U388 ( .A1(n551), .A2(n525), .ZN(n495) );
  OR2_X1 U389 ( .A1(n668), .A2(n667), .ZN(n399) );
  XNOR2_X1 U390 ( .A(n384), .B(G472), .ZN(n671) );
  NOR2_X1 U391 ( .A1(G902), .A2(n697), .ZN(n437) );
  XOR2_X1 U392 ( .A(G119), .B(KEYINPUT71), .Z(n467) );
  XNOR2_X1 U393 ( .A(n649), .B(n650), .ZN(n347) );
  BUF_X1 U394 ( .A(n691), .Z(n348) );
  XNOR2_X1 U395 ( .A(n649), .B(n650), .ZN(n620) );
  NAND2_X1 U396 ( .A1(n409), .A2(n408), .ZN(n486) );
  XNOR2_X1 U397 ( .A(KEYINPUT4), .B(G101), .ZN(n468) );
  XNOR2_X1 U398 ( .A(n538), .B(KEYINPUT1), .ZN(n668) );
  XNOR2_X1 U399 ( .A(n479), .B(n480), .ZN(n356) );
  XNOR2_X1 U400 ( .A(n671), .B(n383), .ZN(n609) );
  INV_X1 U401 ( .A(KEYINPUT6), .ZN(n383) );
  XNOR2_X1 U402 ( .A(n725), .B(G146), .ZN(n469) );
  XNOR2_X1 U403 ( .A(G137), .B(G140), .ZN(n441) );
  BUF_X1 U404 ( .A(n619), .Z(n373) );
  XOR2_X1 U405 ( .A(KEYINPUT20), .B(KEYINPUT89), .Z(n451) );
  NAND2_X1 U406 ( .A1(n388), .A2(n387), .ZN(n510) );
  NAND2_X1 U407 ( .A1(n486), .A2(n440), .ZN(n387) );
  XNOR2_X1 U408 ( .A(G902), .B(KEYINPUT15), .ZN(n619) );
  INV_X1 U409 ( .A(KEYINPUT74), .ZN(n580) );
  XNOR2_X1 U410 ( .A(n517), .B(n425), .ZN(n548) );
  XNOR2_X1 U411 ( .A(n516), .B(n426), .ZN(n425) );
  OR2_X1 U412 ( .A1(n621), .A2(G902), .ZN(n384) );
  XNOR2_X1 U413 ( .A(n563), .B(KEYINPUT48), .ZN(n386) );
  XNOR2_X1 U414 ( .A(G113), .B(KEYINPUT3), .ZN(n466) );
  XNOR2_X1 U415 ( .A(G119), .B(G128), .ZN(n442) );
  XNOR2_X1 U416 ( .A(n512), .B(n511), .ZN(n423) );
  XNOR2_X1 U417 ( .A(G113), .B(KEYINPUT12), .ZN(n507) );
  INV_X1 U418 ( .A(n510), .ZN(n421) );
  XNOR2_X1 U419 ( .A(n487), .B(n357), .ZN(n427) );
  XNOR2_X1 U420 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n357) );
  BUF_X1 U421 ( .A(n668), .Z(n371) );
  NOR2_X1 U422 ( .A1(n532), .A2(n531), .ZN(n533) );
  INV_X1 U423 ( .A(KEYINPUT22), .ZN(n411) );
  AND2_X1 U424 ( .A1(n585), .A2(n664), .ZN(n410) );
  NOR2_X1 U425 ( .A1(n371), .A2(n609), .ZN(n585) );
  NAND2_X1 U426 ( .A1(n415), .A2(n413), .ZN(n412) );
  NOR2_X1 U427 ( .A1(n414), .A2(n710), .ZN(n413) );
  NAND2_X1 U428 ( .A1(n419), .A2(n354), .ZN(n415) );
  XOR2_X1 U429 ( .A(G110), .B(KEYINPUT16), .Z(n485) );
  NOR2_X1 U430 ( .A1(n373), .A2(n379), .ZN(n378) );
  INV_X1 U431 ( .A(G469), .ZN(n379) );
  XNOR2_X1 U432 ( .A(n469), .B(n406), .ZN(n697) );
  XNOR2_X1 U433 ( .A(n407), .B(n431), .ZN(n406) );
  XNOR2_X1 U434 ( .A(n434), .B(n435), .ZN(n407) );
  XNOR2_X1 U435 ( .A(n453), .B(n452), .ZN(n455) );
  XOR2_X1 U436 ( .A(G116), .B(KEYINPUT93), .Z(n471) );
  XNOR2_X1 U437 ( .A(KEYINPUT94), .B(KEYINPUT76), .ZN(n472) );
  XOR2_X1 U438 ( .A(KEYINPUT92), .B(KEYINPUT5), .Z(n473) );
  XNOR2_X1 U439 ( .A(n424), .B(KEYINPUT103), .ZN(n657) );
  OR2_X1 U440 ( .A1(n548), .A2(n549), .ZN(n424) );
  NOR2_X1 U441 ( .A1(G902), .A2(G237), .ZN(n478) );
  NOR2_X1 U442 ( .A1(n373), .A2(n418), .ZN(n417) );
  INV_X1 U443 ( .A(G472), .ZN(n418) );
  INV_X1 U444 ( .A(G134), .ZN(n429) );
  XNOR2_X1 U445 ( .A(n498), .B(n363), .ZN(n362) );
  INV_X1 U446 ( .A(KEYINPUT7), .ZN(n363) );
  XNOR2_X1 U447 ( .A(G122), .B(KEYINPUT9), .ZN(n498) );
  XNOR2_X1 U448 ( .A(n433), .B(n432), .ZN(n434) );
  INV_X1 U449 ( .A(G110), .ZN(n432) );
  XOR2_X1 U450 ( .A(G107), .B(G104), .Z(n435) );
  INV_X1 U451 ( .A(KEYINPUT33), .ZN(n368) );
  NOR2_X1 U452 ( .A1(n356), .A2(n520), .ZN(n481) );
  INV_X1 U453 ( .A(KEYINPUT0), .ZN(n578) );
  BUF_X1 U454 ( .A(n671), .Z(n375) );
  XOR2_X1 U455 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n447) );
  XNOR2_X1 U456 ( .A(n422), .B(n420), .ZN(n700) );
  XNOR2_X1 U457 ( .A(n515), .B(n421), .ZN(n420) );
  XNOR2_X1 U458 ( .A(n514), .B(n423), .ZN(n422) );
  XNOR2_X1 U459 ( .A(n489), .B(n488), .ZN(n490) );
  INV_X1 U460 ( .A(G210), .ZN(n381) );
  NOR2_X1 U461 ( .A1(n539), .A2(n371), .ZN(n643) );
  INV_X1 U462 ( .A(KEYINPUT36), .ZN(n536) );
  INV_X1 U463 ( .A(KEYINPUT35), .ZN(n400) );
  INV_X1 U464 ( .A(n582), .ZN(n402) );
  XNOR2_X1 U465 ( .A(n586), .B(n364), .ZN(n740) );
  XNOR2_X1 U466 ( .A(n365), .B(KEYINPUT32), .ZN(n364) );
  INV_X1 U467 ( .A(KEYINPUT64), .ZN(n365) );
  XNOR2_X1 U468 ( .A(KEYINPUT102), .B(n541), .ZN(n641) );
  INV_X1 U469 ( .A(KEYINPUT105), .ZN(n393) );
  INV_X1 U470 ( .A(n664), .ZN(n610) );
  INV_X1 U471 ( .A(KEYINPUT63), .ZN(n366) );
  NOR2_X1 U472 ( .A1(n416), .A2(n412), .ZN(n622) );
  XNOR2_X1 U473 ( .A(n695), .B(n372), .ZN(n698) );
  XNOR2_X1 U474 ( .A(n697), .B(n696), .ZN(n372) );
  XNOR2_X1 U475 ( .A(n404), .B(n403), .ZN(G75) );
  XNOR2_X1 U476 ( .A(KEYINPUT53), .B(KEYINPUT123), .ZN(n403) );
  OR2_X1 U477 ( .A1(n653), .A2(n405), .ZN(n404) );
  NAND2_X1 U478 ( .A1(n690), .A2(n729), .ZN(n405) );
  XOR2_X1 U479 ( .A(n492), .B(KEYINPUT86), .Z(n349) );
  XOR2_X1 U480 ( .A(n476), .B(n475), .Z(n350) );
  AND2_X1 U481 ( .A1(n409), .A2(KEYINPUT10), .ZN(n351) );
  XOR2_X1 U482 ( .A(n455), .B(n454), .Z(n352) );
  XOR2_X1 U483 ( .A(n621), .B(KEYINPUT62), .Z(n353) );
  AND2_X1 U484 ( .A1(n353), .A2(n417), .ZN(n354) );
  NOR2_X1 U485 ( .A1(n373), .A2(n381), .ZN(n355) );
  NOR2_X1 U486 ( .A1(G952), .A2(n729), .ZN(n710) );
  INV_X1 U487 ( .A(G475), .ZN(n426) );
  NOR2_X2 U488 ( .A1(n587), .A2(n665), .ZN(n458) );
  XNOR2_X2 U489 ( .A(n370), .B(G128), .ZN(n487) );
  INV_X1 U490 ( .A(n620), .ZN(n377) );
  BUF_X1 U491 ( .A(n587), .Z(n358) );
  XNOR2_X1 U492 ( .A(n359), .B(KEYINPUT34), .ZN(n581) );
  NOR2_X2 U493 ( .A1(n687), .A2(n599), .ZN(n359) );
  XNOR2_X2 U494 ( .A(n360), .B(n411), .ZN(n588) );
  NAND2_X1 U495 ( .A1(n601), .A2(n584), .ZN(n360) );
  XOR2_X2 U496 ( .A(G116), .B(G107), .Z(n497) );
  XNOR2_X2 U497 ( .A(n497), .B(n505), .ZN(n484) );
  XNOR2_X2 U498 ( .A(n361), .B(n352), .ZN(n587) );
  OR2_X2 U499 ( .A1(n708), .A2(G902), .ZN(n361) );
  NOR2_X1 U500 ( .A1(n590), .A2(n591), .ZN(n628) );
  XNOR2_X1 U501 ( .A(n497), .B(n362), .ZN(n499) );
  NAND2_X1 U502 ( .A1(n576), .A2(n577), .ZN(n579) );
  XOR2_X2 U503 ( .A(G122), .B(G104), .Z(n505) );
  XNOR2_X1 U504 ( .A(n622), .B(n366), .ZN(G57) );
  XNOR2_X1 U505 ( .A(n367), .B(KEYINPUT60), .ZN(G60) );
  NOR2_X2 U506 ( .A1(n703), .A2(n710), .ZN(n367) );
  XNOR2_X1 U507 ( .A(n632), .B(KEYINPUT82), .ZN(n553) );
  XNOR2_X2 U508 ( .A(n369), .B(n368), .ZN(n687) );
  NAND2_X1 U509 ( .A1(n597), .A2(n609), .ZN(n369) );
  XNOR2_X2 U510 ( .A(n487), .B(n429), .ZN(n502) );
  NAND2_X2 U511 ( .A1(n386), .A2(n385), .ZN(n649) );
  XNOR2_X1 U512 ( .A(n477), .B(n350), .ZN(n621) );
  XNOR2_X1 U513 ( .A(n374), .B(KEYINPUT56), .ZN(G51) );
  NOR2_X2 U514 ( .A1(n694), .A2(n710), .ZN(n374) );
  NAND2_X1 U515 ( .A1(n588), .A2(n410), .ZN(n586) );
  XNOR2_X2 U516 ( .A(n467), .B(n466), .ZN(n711) );
  XNOR2_X2 U517 ( .A(n711), .B(n468), .ZN(n489) );
  NOR2_X2 U518 ( .A1(n608), .A2(n375), .ZN(n589) );
  XNOR2_X1 U519 ( .A(n602), .B(n459), .ZN(n482) );
  NOR2_X2 U520 ( .A1(n667), .A2(n538), .ZN(n390) );
  NAND2_X1 U521 ( .A1(n617), .A2(n616), .ZN(n618) );
  AND2_X2 U522 ( .A1(n376), .A2(n571), .ZN(n385) );
  NAND2_X1 U523 ( .A1(n376), .A2(n729), .ZN(n716) );
  XNOR2_X2 U524 ( .A(n618), .B(KEYINPUT45), .ZN(n376) );
  NAND2_X1 U525 ( .A1(n419), .A2(n378), .ZN(n695) );
  NAND2_X1 U526 ( .A1(n377), .A2(n355), .ZN(n693) );
  NAND2_X1 U527 ( .A1(n377), .A2(n380), .ZN(n702) );
  NOR2_X1 U528 ( .A1(n347), .A2(n373), .ZN(n382) );
  NOR2_X1 U529 ( .A1(n373), .A2(n426), .ZN(n380) );
  NAND2_X1 U530 ( .A1(n382), .A2(G478), .ZN(n704) );
  NAND2_X1 U531 ( .A1(n382), .A2(G217), .ZN(n707) );
  AND2_X1 U532 ( .A1(n386), .A2(n571), .ZN(n727) );
  NAND2_X1 U533 ( .A1(n351), .A2(n408), .ZN(n388) );
  XNOR2_X2 U534 ( .A(n458), .B(n391), .ZN(n667) );
  INV_X1 U535 ( .A(n550), .ZN(n544) );
  XNOR2_X2 U536 ( .A(n493), .B(n349), .ZN(n550) );
  XNOR2_X2 U537 ( .A(n394), .B(n393), .ZN(n743) );
  NAND2_X1 U538 ( .A1(n395), .A2(n610), .ZN(n394) );
  XNOR2_X1 U539 ( .A(n396), .B(KEYINPUT84), .ZN(n395) );
  NOR2_X1 U540 ( .A1(n608), .A2(n609), .ZN(n396) );
  XNOR2_X1 U541 ( .A(n397), .B(n490), .ZN(n691) );
  XNOR2_X1 U542 ( .A(n398), .B(n713), .ZN(n397) );
  XNOR2_X1 U543 ( .A(n427), .B(n486), .ZN(n398) );
  XNOR2_X2 U544 ( .A(n399), .B(n580), .ZN(n597) );
  XNOR2_X2 U545 ( .A(n437), .B(n436), .ZN(n538) );
  NAND2_X1 U546 ( .A1(n595), .A2(n742), .ZN(n592) );
  XNOR2_X2 U547 ( .A(n401), .B(n400), .ZN(n742) );
  NAND2_X1 U548 ( .A1(n581), .A2(n402), .ZN(n401) );
  NAND2_X1 U549 ( .A1(n438), .A2(G146), .ZN(n408) );
  NAND2_X1 U550 ( .A1(n439), .A2(G125), .ZN(n409) );
  NOR2_X1 U551 ( .A1(n353), .A2(n417), .ZN(n414) );
  NOR2_X1 U552 ( .A1(n419), .A2(n353), .ZN(n416) );
  INV_X1 U553 ( .A(n347), .ZN(n419) );
  XNOR2_X1 U554 ( .A(n693), .B(n692), .ZN(n694) );
  XNOR2_X1 U555 ( .A(n702), .B(n701), .ZN(n703) );
  XNOR2_X1 U556 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n428) );
  INV_X1 U557 ( .A(n665), .ZN(n583) );
  AND2_X1 U558 ( .A1(n657), .A2(n583), .ZN(n584) );
  INV_X1 U559 ( .A(KEYINPUT109), .ZN(n459) );
  INV_X1 U560 ( .A(KEYINPUT25), .ZN(n452) );
  INV_X1 U561 ( .A(n646), .ZN(n570) );
  XNOR2_X1 U562 ( .A(n430), .B(n441), .ZN(n431) );
  NOR2_X1 U563 ( .A1(n739), .A2(n570), .ZN(n571) );
  INV_X1 U564 ( .A(KEYINPUT59), .ZN(n699) );
  XNOR2_X1 U565 ( .A(n700), .B(n699), .ZN(n701) );
  XOR2_X1 U566 ( .A(KEYINPUT68), .B(G131), .Z(n513) );
  INV_X1 U567 ( .A(n468), .ZN(n430) );
  AND2_X1 U568 ( .A1(G227), .A2(n729), .ZN(n433) );
  XNOR2_X1 U569 ( .A(KEYINPUT70), .B(G469), .ZN(n436) );
  INV_X1 U570 ( .A(G125), .ZN(n438) );
  INV_X1 U571 ( .A(G146), .ZN(n439) );
  INV_X1 U572 ( .A(KEYINPUT10), .ZN(n440) );
  XOR2_X1 U573 ( .A(KEYINPUT72), .B(G110), .Z(n443) );
  XNOR2_X1 U574 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U575 ( .A(n723), .B(n444), .ZN(n449) );
  NAND2_X1 U576 ( .A1(G234), .A2(n729), .ZN(n445) );
  XOR2_X1 U577 ( .A(KEYINPUT8), .B(n445), .Z(n496) );
  NAND2_X1 U578 ( .A1(G221), .A2(n496), .ZN(n446) );
  XNOR2_X1 U579 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U580 ( .A(n449), .B(n448), .ZN(n708) );
  NAND2_X1 U581 ( .A1(G234), .A2(n619), .ZN(n450) );
  XNOR2_X1 U582 ( .A(n451), .B(n450), .ZN(n456) );
  NAND2_X1 U583 ( .A1(n456), .A2(G217), .ZN(n453) );
  XNOR2_X1 U584 ( .A(KEYINPUT88), .B(KEYINPUT90), .ZN(n454) );
  NAND2_X1 U585 ( .A1(n456), .A2(G221), .ZN(n457) );
  XNOR2_X1 U586 ( .A(n457), .B(KEYINPUT21), .ZN(n665) );
  NAND2_X1 U587 ( .A1(G234), .A2(G237), .ZN(n460) );
  XNOR2_X1 U588 ( .A(n460), .B(KEYINPUT14), .ZN(n461) );
  NAND2_X1 U589 ( .A1(G952), .A2(n461), .ZN(n684) );
  NOR2_X1 U590 ( .A1(G953), .A2(n684), .ZN(n573) );
  NAND2_X1 U591 ( .A1(n461), .A2(G902), .ZN(n462) );
  XNOR2_X1 U592 ( .A(n462), .B(KEYINPUT87), .ZN(n572) );
  NAND2_X1 U593 ( .A1(n572), .A2(G953), .ZN(n463) );
  NOR2_X1 U594 ( .A1(G900), .A2(n463), .ZN(n464) );
  NOR2_X1 U595 ( .A1(n573), .A2(n464), .ZN(n520) );
  XOR2_X1 U596 ( .A(KEYINPUT111), .B(KEYINPUT30), .Z(n465) );
  XNOR2_X1 U597 ( .A(KEYINPUT110), .B(n465), .ZN(n480) );
  XNOR2_X1 U598 ( .A(n469), .B(n489), .ZN(n477) );
  NOR2_X1 U599 ( .A1(G953), .A2(G237), .ZN(n509) );
  NAND2_X1 U600 ( .A1(n509), .A2(G210), .ZN(n470) );
  XNOR2_X1 U601 ( .A(n471), .B(n470), .ZN(n476) );
  XNOR2_X1 U602 ( .A(n473), .B(n472), .ZN(n474) );
  XOR2_X1 U603 ( .A(n474), .B(G137), .Z(n475) );
  XNOR2_X1 U604 ( .A(n478), .B(KEYINPUT75), .ZN(n491) );
  NAND2_X1 U605 ( .A1(G214), .A2(n491), .ZN(n658) );
  NAND2_X1 U606 ( .A1(n671), .A2(n658), .ZN(n479) );
  NAND2_X1 U607 ( .A1(n482), .A2(n481), .ZN(n483) );
  NAND2_X1 U608 ( .A1(G224), .A2(n729), .ZN(n488) );
  NAND2_X1 U609 ( .A1(n691), .A2(n373), .ZN(n493) );
  NAND2_X1 U610 ( .A1(n491), .A2(G210), .ZN(n492) );
  XOR2_X1 U611 ( .A(KEYINPUT38), .B(n544), .Z(n655) );
  INV_X1 U612 ( .A(n655), .ZN(n525) );
  XOR2_X1 U613 ( .A(KEYINPUT73), .B(KEYINPUT39), .Z(n494) );
  NAND2_X1 U614 ( .A1(n496), .A2(G217), .ZN(n500) );
  XNOR2_X1 U615 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U616 ( .A(n502), .B(n501), .ZN(n705) );
  NOR2_X1 U617 ( .A1(G902), .A2(n705), .ZN(n504) );
  XNOR2_X1 U618 ( .A(KEYINPUT101), .B(G478), .ZN(n503) );
  XNOR2_X1 U619 ( .A(n504), .B(n503), .ZN(n549) );
  XNOR2_X1 U620 ( .A(G143), .B(G140), .ZN(n506) );
  XNOR2_X1 U621 ( .A(n506), .B(n505), .ZN(n515) );
  XOR2_X1 U622 ( .A(KEYINPUT11), .B(KEYINPUT97), .Z(n508) );
  XNOR2_X1 U623 ( .A(n508), .B(n507), .ZN(n512) );
  NAND2_X1 U624 ( .A1(G214), .A2(n509), .ZN(n511) );
  XNOR2_X1 U625 ( .A(n513), .B(KEYINPUT98), .ZN(n514) );
  NOR2_X1 U626 ( .A1(G902), .A2(n700), .ZN(n517) );
  XNOR2_X1 U627 ( .A(KEYINPUT13), .B(KEYINPUT99), .ZN(n516) );
  XOR2_X1 U628 ( .A(KEYINPUT100), .B(n548), .Z(n540) );
  OR2_X1 U629 ( .A1(n549), .A2(n540), .ZN(n542) );
  XNOR2_X1 U630 ( .A(KEYINPUT112), .B(KEYINPUT40), .ZN(n518) );
  XNOR2_X1 U631 ( .A(n519), .B(n518), .ZN(n737) );
  INV_X1 U632 ( .A(n375), .ZN(n522) );
  NOR2_X1 U633 ( .A1(n520), .A2(n665), .ZN(n521) );
  NAND2_X1 U634 ( .A1(n358), .A2(n521), .ZN(n532) );
  NOR2_X1 U635 ( .A1(n522), .A2(n532), .ZN(n523) );
  XOR2_X1 U636 ( .A(KEYINPUT28), .B(n523), .Z(n524) );
  NOR2_X1 U637 ( .A1(n538), .A2(n524), .ZN(n545) );
  AND2_X1 U638 ( .A1(n525), .A2(n657), .ZN(n662) );
  NAND2_X1 U639 ( .A1(n662), .A2(n658), .ZN(n526) );
  XNOR2_X1 U640 ( .A(KEYINPUT41), .B(n526), .ZN(n685) );
  NAND2_X1 U641 ( .A1(n545), .A2(n685), .ZN(n527) );
  XNOR2_X1 U642 ( .A(n527), .B(KEYINPUT42), .ZN(n528) );
  XNOR2_X1 U643 ( .A(KEYINPUT113), .B(n528), .ZN(n744) );
  NOR2_X1 U644 ( .A1(n737), .A2(n744), .ZN(n530) );
  XNOR2_X1 U645 ( .A(KEYINPUT46), .B(KEYINPUT83), .ZN(n529) );
  XNOR2_X1 U646 ( .A(n530), .B(n529), .ZN(n562) );
  XNOR2_X1 U647 ( .A(n542), .B(KEYINPUT106), .ZN(n637) );
  INV_X1 U648 ( .A(n609), .ZN(n531) );
  XNOR2_X1 U649 ( .A(n533), .B(KEYINPUT107), .ZN(n534) );
  NOR2_X1 U650 ( .A1(n637), .A2(n534), .ZN(n535) );
  NAND2_X1 U651 ( .A1(n535), .A2(n658), .ZN(n566) );
  NOR2_X1 U652 ( .A1(n566), .A2(n544), .ZN(n537) );
  XNOR2_X1 U653 ( .A(n537), .B(n536), .ZN(n539) );
  NAND2_X1 U654 ( .A1(n540), .A2(n549), .ZN(n541) );
  AND2_X1 U655 ( .A1(n542), .A2(n641), .ZN(n654) );
  NAND2_X1 U656 ( .A1(n654), .A2(KEYINPUT47), .ZN(n543) );
  XNOR2_X1 U657 ( .A(n543), .B(KEYINPUT80), .ZN(n547) );
  NAND2_X1 U658 ( .A1(n545), .A2(n576), .ZN(n634) );
  NAND2_X1 U659 ( .A1(n634), .A2(KEYINPUT47), .ZN(n546) );
  NAND2_X1 U660 ( .A1(n547), .A2(n546), .ZN(n554) );
  NAND2_X1 U661 ( .A1(n549), .A2(n548), .ZN(n582) );
  NAND2_X1 U662 ( .A1(n551), .A2(n550), .ZN(n552) );
  NOR2_X1 U663 ( .A1(n554), .A2(n553), .ZN(n558) );
  XNOR2_X1 U664 ( .A(KEYINPUT47), .B(KEYINPUT67), .ZN(n556) );
  XOR2_X1 U665 ( .A(n654), .B(KEYINPUT81), .Z(n605) );
  NOR2_X1 U666 ( .A1(n634), .A2(n605), .ZN(n555) );
  NAND2_X1 U667 ( .A1(n556), .A2(n555), .ZN(n557) );
  NAND2_X1 U668 ( .A1(n558), .A2(n557), .ZN(n559) );
  NOR2_X1 U669 ( .A1(n643), .A2(n559), .ZN(n560) );
  XNOR2_X1 U670 ( .A(n560), .B(KEYINPUT69), .ZN(n561) );
  OR2_X1 U671 ( .A1(n564), .A2(n641), .ZN(n565) );
  XOR2_X1 U672 ( .A(KEYINPUT114), .B(n565), .Z(n739) );
  XOR2_X1 U673 ( .A(KEYINPUT108), .B(n566), .Z(n567) );
  NAND2_X1 U674 ( .A1(n567), .A2(n371), .ZN(n568) );
  XNOR2_X1 U675 ( .A(KEYINPUT43), .B(n568), .ZN(n569) );
  NAND2_X1 U676 ( .A1(n569), .A2(n544), .ZN(n646) );
  NOR2_X1 U677 ( .A1(G898), .A2(n729), .ZN(n715) );
  NAND2_X1 U678 ( .A1(n715), .A2(n572), .ZN(n575) );
  INV_X1 U679 ( .A(n573), .ZN(n574) );
  NAND2_X1 U680 ( .A1(n575), .A2(n574), .ZN(n577) );
  XNOR2_X2 U681 ( .A(n579), .B(n578), .ZN(n601) );
  INV_X1 U682 ( .A(n601), .ZN(n599) );
  XNOR2_X1 U683 ( .A(n358), .B(KEYINPUT104), .ZN(n664) );
  INV_X1 U684 ( .A(n358), .ZN(n591) );
  NAND2_X1 U685 ( .A1(n588), .A2(n371), .ZN(n608) );
  XNOR2_X1 U686 ( .A(n589), .B(KEYINPUT65), .ZN(n590) );
  NOR2_X1 U687 ( .A1(n740), .A2(n628), .ZN(n595) );
  XNOR2_X1 U688 ( .A(n592), .B(KEYINPUT44), .ZN(n594) );
  INV_X1 U689 ( .A(KEYINPUT85), .ZN(n593) );
  NAND2_X1 U690 ( .A1(n594), .A2(n593), .ZN(n617) );
  NAND2_X1 U691 ( .A1(KEYINPUT44), .A2(n595), .ZN(n596) );
  NAND2_X1 U692 ( .A1(n596), .A2(KEYINPUT85), .ZN(n613) );
  NAND2_X1 U693 ( .A1(n597), .A2(n375), .ZN(n598) );
  XNOR2_X1 U694 ( .A(n598), .B(KEYINPUT96), .ZN(n676) );
  NOR2_X1 U695 ( .A1(n676), .A2(n599), .ZN(n600) );
  XNOR2_X1 U696 ( .A(n600), .B(KEYINPUT31), .ZN(n640) );
  NAND2_X1 U697 ( .A1(n602), .A2(n601), .ZN(n603) );
  NOR2_X1 U698 ( .A1(n375), .A2(n603), .ZN(n604) );
  XNOR2_X1 U699 ( .A(n604), .B(KEYINPUT95), .ZN(n624) );
  NAND2_X1 U700 ( .A1(n640), .A2(n624), .ZN(n607) );
  INV_X1 U701 ( .A(n605), .ZN(n606) );
  NAND2_X1 U702 ( .A1(n607), .A2(n606), .ZN(n611) );
  NAND2_X1 U703 ( .A1(n613), .A2(n612), .ZN(n615) );
  AND2_X1 U704 ( .A1(n742), .A2(KEYINPUT85), .ZN(n614) );
  INV_X1 U705 ( .A(KEYINPUT2), .ZN(n650) );
  NOR2_X1 U706 ( .A1(n637), .A2(n624), .ZN(n623) );
  XOR2_X1 U707 ( .A(G104), .B(n623), .Z(G6) );
  NOR2_X1 U708 ( .A1(n641), .A2(n624), .ZN(n626) );
  XNOR2_X1 U709 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n625) );
  XNOR2_X1 U710 ( .A(n626), .B(n625), .ZN(n627) );
  XNOR2_X1 U711 ( .A(G107), .B(n627), .ZN(G9) );
  XOR2_X1 U712 ( .A(n628), .B(G110), .Z(G12) );
  NOR2_X1 U713 ( .A1(n641), .A2(n634), .ZN(n630) );
  XNOR2_X1 U714 ( .A(KEYINPUT115), .B(KEYINPUT29), .ZN(n629) );
  XNOR2_X1 U715 ( .A(n630), .B(n629), .ZN(n631) );
  XOR2_X1 U716 ( .A(G128), .B(n631), .Z(G30) );
  XOR2_X1 U717 ( .A(G143), .B(n632), .Z(n633) );
  XNOR2_X1 U718 ( .A(KEYINPUT116), .B(n633), .ZN(G45) );
  NOR2_X1 U719 ( .A1(n637), .A2(n634), .ZN(n636) );
  XNOR2_X1 U720 ( .A(G146), .B(KEYINPUT117), .ZN(n635) );
  XNOR2_X1 U721 ( .A(n636), .B(n635), .ZN(G48) );
  NOR2_X1 U722 ( .A1(n637), .A2(n640), .ZN(n638) );
  XOR2_X1 U723 ( .A(KEYINPUT118), .B(n638), .Z(n639) );
  XNOR2_X1 U724 ( .A(G113), .B(n639), .ZN(G15) );
  NOR2_X1 U725 ( .A1(n641), .A2(n640), .ZN(n642) );
  XOR2_X1 U726 ( .A(G116), .B(n642), .Z(G18) );
  XOR2_X1 U727 ( .A(KEYINPUT37), .B(KEYINPUT119), .Z(n645) );
  XNOR2_X1 U728 ( .A(G125), .B(n643), .ZN(n644) );
  XNOR2_X1 U729 ( .A(n645), .B(n644), .ZN(G27) );
  XNOR2_X1 U730 ( .A(G140), .B(n646), .ZN(G42) );
  XNOR2_X1 U731 ( .A(KEYINPUT79), .B(KEYINPUT2), .ZN(n647) );
  NAND2_X1 U732 ( .A1(n647), .A2(n649), .ZN(n648) );
  XOR2_X1 U733 ( .A(KEYINPUT78), .B(n648), .Z(n652) );
  NOR2_X1 U734 ( .A1(n650), .A2(n649), .ZN(n651) );
  NOR2_X1 U735 ( .A1(n652), .A2(n651), .ZN(n653) );
  NOR2_X1 U736 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U737 ( .A1(n657), .A2(n656), .ZN(n660) );
  INV_X1 U738 ( .A(n658), .ZN(n659) );
  NOR2_X1 U739 ( .A1(n660), .A2(n659), .ZN(n661) );
  NOR2_X1 U740 ( .A1(n662), .A2(n661), .ZN(n663) );
  NOR2_X1 U741 ( .A1(n687), .A2(n663), .ZN(n681) );
  NAND2_X1 U742 ( .A1(n665), .A2(n664), .ZN(n666) );
  XOR2_X1 U743 ( .A(KEYINPUT49), .B(n666), .Z(n674) );
  NAND2_X1 U744 ( .A1(n371), .A2(n667), .ZN(n669) );
  XNOR2_X1 U745 ( .A(n669), .B(KEYINPUT50), .ZN(n670) );
  XNOR2_X1 U746 ( .A(KEYINPUT121), .B(n670), .ZN(n672) );
  NOR2_X1 U747 ( .A1(n672), .A2(n375), .ZN(n673) );
  NAND2_X1 U748 ( .A1(n674), .A2(n673), .ZN(n675) );
  NAND2_X1 U749 ( .A1(n676), .A2(n675), .ZN(n677) );
  XOR2_X1 U750 ( .A(KEYINPUT51), .B(n677), .Z(n678) );
  NAND2_X1 U751 ( .A1(n685), .A2(n678), .ZN(n679) );
  XOR2_X1 U752 ( .A(KEYINPUT122), .B(n679), .Z(n680) );
  NOR2_X1 U753 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U754 ( .A(n682), .B(KEYINPUT52), .ZN(n683) );
  NOR2_X1 U755 ( .A1(n684), .A2(n683), .ZN(n689) );
  INV_X1 U756 ( .A(n685), .ZN(n686) );
  NOR2_X1 U757 ( .A1(n687), .A2(n686), .ZN(n688) );
  NOR2_X1 U758 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U759 ( .A(n348), .B(n428), .ZN(n692) );
  XOR2_X1 U760 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n696) );
  NOR2_X1 U761 ( .A1(n710), .A2(n698), .ZN(G54) );
  XNOR2_X1 U762 ( .A(n705), .B(n704), .ZN(n706) );
  NOR2_X1 U763 ( .A1(n710), .A2(n706), .ZN(G63) );
  XNOR2_X1 U764 ( .A(n708), .B(n707), .ZN(n709) );
  NOR2_X1 U765 ( .A1(n710), .A2(n709), .ZN(G66) );
  XOR2_X1 U766 ( .A(G101), .B(n711), .Z(n712) );
  XNOR2_X1 U767 ( .A(n713), .B(n712), .ZN(n714) );
  NOR2_X1 U768 ( .A1(n715), .A2(n714), .ZN(n722) );
  XNOR2_X1 U769 ( .A(KEYINPUT124), .B(n716), .ZN(n720) );
  NAND2_X1 U770 ( .A1(G953), .A2(G224), .ZN(n717) );
  XNOR2_X1 U771 ( .A(KEYINPUT61), .B(n717), .ZN(n718) );
  NAND2_X1 U772 ( .A1(n718), .A2(G898), .ZN(n719) );
  NAND2_X1 U773 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U774 ( .A(n722), .B(n721), .ZN(G69) );
  XOR2_X1 U775 ( .A(n723), .B(KEYINPUT125), .Z(n724) );
  XNOR2_X1 U776 ( .A(n725), .B(n724), .ZN(n726) );
  XNOR2_X1 U777 ( .A(KEYINPUT4), .B(n726), .ZN(n731) );
  INV_X1 U778 ( .A(n731), .ZN(n728) );
  XNOR2_X1 U779 ( .A(n728), .B(n727), .ZN(n730) );
  NAND2_X1 U780 ( .A1(n730), .A2(n729), .ZN(n736) );
  XNOR2_X1 U781 ( .A(G227), .B(KEYINPUT126), .ZN(n732) );
  XNOR2_X1 U782 ( .A(n732), .B(n731), .ZN(n733) );
  NAND2_X1 U783 ( .A1(G900), .A2(n733), .ZN(n734) );
  NAND2_X1 U784 ( .A1(n734), .A2(G953), .ZN(n735) );
  NAND2_X1 U785 ( .A1(n736), .A2(n735), .ZN(G72) );
  XOR2_X1 U786 ( .A(n737), .B(G131), .Z(G33) );
  XOR2_X1 U787 ( .A(G134), .B(KEYINPUT120), .Z(n738) );
  XNOR2_X1 U788 ( .A(n739), .B(n738), .ZN(G36) );
  XOR2_X1 U789 ( .A(n740), .B(G119), .Z(G21) );
  XOR2_X1 U790 ( .A(G122), .B(KEYINPUT127), .Z(n741) );
  XNOR2_X1 U791 ( .A(n742), .B(n741), .ZN(G24) );
  XNOR2_X1 U792 ( .A(n743), .B(G101), .ZN(G3) );
  XOR2_X1 U793 ( .A(G137), .B(n744), .Z(G39) );
endmodule

