//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 1 0 0 1 1 0 1 1 0 1 0 0 0 0 1 1 0 0 0 1 0 0 1 1 0 0 1 0 0 1 0 0 1 0 1 1 1 1 1 1 0 0 1 1 1 0 1 1 1 1 0 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:59 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n681, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n909, new_n910, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n929,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  INV_X1    g001(.A(G119), .ZN(new_n188));
  OAI21_X1  g002(.A(KEYINPUT67), .B1(new_n188), .B2(G116), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT67), .ZN(new_n190));
  INV_X1    g004(.A(G116), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n190), .A2(new_n191), .A3(G119), .ZN(new_n192));
  AND2_X1   g006(.A1(new_n189), .A2(new_n192), .ZN(new_n193));
  XOR2_X1   g007(.A(KEYINPUT2), .B(G113), .Z(new_n194));
  OAI21_X1  g008(.A(KEYINPUT66), .B1(new_n191), .B2(G119), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT66), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n196), .A2(new_n188), .A3(G116), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n193), .A2(new_n194), .A3(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n194), .B1(new_n193), .B2(new_n198), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  NOR2_X1   g017(.A1(KEYINPUT0), .A2(G128), .ZN(new_n204));
  XNOR2_X1  g018(.A(G143), .B(G146), .ZN(new_n205));
  NAND2_X1  g019(.A1(KEYINPUT0), .A2(G128), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G143), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n208), .A2(G146), .ZN(new_n209));
  INV_X1    g023(.A(G146), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n210), .A2(G143), .ZN(new_n211));
  OAI211_X1 g025(.A(KEYINPUT0), .B(G128), .C1(new_n209), .C2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n207), .A2(new_n212), .ZN(new_n213));
  XOR2_X1   g027(.A(KEYINPUT65), .B(G131), .Z(new_n214));
  INV_X1    g028(.A(G134), .ZN(new_n215));
  OAI21_X1  g029(.A(KEYINPUT64), .B1(new_n215), .B2(G137), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(KEYINPUT11), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT11), .ZN(new_n218));
  OAI211_X1 g032(.A(KEYINPUT64), .B(new_n218), .C1(new_n215), .C2(G137), .ZN(new_n219));
  INV_X1    g033(.A(G137), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n220), .A2(G134), .ZN(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  AND4_X1   g036(.A1(new_n214), .A2(new_n217), .A3(new_n219), .A4(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G131), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n221), .B1(new_n216), .B2(KEYINPUT11), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n224), .B1(new_n225), .B2(new_n219), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n213), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT30), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT1), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n229), .B1(G143), .B2(new_n210), .ZN(new_n230));
  INV_X1    g044(.A(G128), .ZN(new_n231));
  OAI22_X1  g045(.A1(new_n230), .A2(new_n231), .B1(new_n209), .B2(new_n211), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n210), .A2(G143), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n208), .A2(G146), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n233), .A2(new_n234), .A3(new_n229), .A4(G128), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n232), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n225), .A2(new_n214), .A3(new_n219), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n215), .A2(G137), .ZN(new_n238));
  OAI21_X1  g052(.A(G131), .B1(new_n238), .B2(new_n221), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n236), .A2(new_n237), .A3(new_n239), .ZN(new_n240));
  AND3_X1   g054(.A1(new_n227), .A2(new_n228), .A3(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT68), .ZN(new_n242));
  INV_X1    g056(.A(new_n235), .ZN(new_n243));
  OAI21_X1  g057(.A(KEYINPUT1), .B1(new_n208), .B2(G146), .ZN(new_n244));
  AOI22_X1  g058(.A1(new_n244), .A2(G128), .B1(new_n233), .B2(new_n234), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n242), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n232), .A2(KEYINPUT68), .A3(new_n235), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n246), .A2(new_n237), .A3(new_n247), .A4(new_n239), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n228), .B1(new_n248), .B2(new_n227), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n203), .B1(new_n241), .B2(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n248), .A2(new_n202), .A3(new_n227), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NOR2_X1   g066(.A1(G237), .A2(G953), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G210), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n254), .B(KEYINPUT27), .ZN(new_n255));
  XNOR2_X1  g069(.A(KEYINPUT26), .B(G101), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n255), .B(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n252), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT29), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n251), .A2(KEYINPUT28), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT28), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n248), .A2(new_n202), .A3(new_n227), .A4(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n227), .A2(new_n240), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(new_n203), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n264), .A2(new_n266), .A3(new_n257), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n259), .A2(new_n260), .A3(new_n267), .ZN(new_n268));
  XNOR2_X1  g082(.A(KEYINPUT71), .B(G902), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n248), .A2(new_n227), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(new_n203), .ZN(new_n272));
  AND2_X1   g086(.A1(new_n264), .A2(new_n272), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n258), .A2(new_n260), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n270), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n187), .B1(new_n268), .B2(new_n275), .ZN(new_n276));
  XNOR2_X1  g090(.A(new_n276), .B(KEYINPUT72), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT32), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT31), .ZN(new_n279));
  AND2_X1   g093(.A1(new_n251), .A2(new_n257), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n250), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(KEYINPUT69), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT69), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n250), .A2(new_n283), .A3(new_n280), .A4(new_n279), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n257), .B1(new_n264), .B2(new_n266), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n279), .B1(new_n250), .B2(new_n280), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(KEYINPUT70), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT70), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n285), .A2(new_n291), .A3(new_n288), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  NOR2_X1   g107(.A1(G472), .A2(G902), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n278), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  AND3_X1   g109(.A1(new_n285), .A2(new_n291), .A3(new_n288), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n291), .B1(new_n285), .B2(new_n288), .ZN(new_n297));
  OAI211_X1 g111(.A(new_n278), .B(new_n294), .C1(new_n296), .C2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n277), .B1(new_n295), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT96), .ZN(new_n301));
  INV_X1    g115(.A(G475), .ZN(new_n302));
  INV_X1    g116(.A(G902), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G237), .ZN(new_n305));
  INV_X1    g119(.A(G953), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n305), .A2(new_n306), .A3(G214), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(new_n208), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n253), .A2(G143), .A3(G214), .ZN(new_n309));
  NAND3_X1  g123(.A1(KEYINPUT92), .A2(KEYINPUT18), .A3(G131), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n310), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n307), .A2(new_n208), .ZN(new_n313));
  AOI21_X1  g127(.A(G143), .B1(new_n253), .B2(G214), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n312), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G140), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G125), .ZN(new_n317));
  INV_X1    g131(.A(G125), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G140), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  OAI21_X1  g134(.A(KEYINPUT76), .B1(new_n320), .B2(G146), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT76), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n317), .A2(new_n319), .A3(new_n322), .A4(new_n210), .ZN(new_n323));
  AND2_X1   g137(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n210), .B1(new_n317), .B2(new_n319), .ZN(new_n325));
  OAI211_X1 g139(.A(new_n311), .B(new_n315), .C1(new_n324), .C2(new_n325), .ZN(new_n326));
  XOR2_X1   g140(.A(G113), .B(G122), .Z(new_n327));
  XOR2_X1   g141(.A(KEYINPUT93), .B(G104), .Z(new_n328));
  XOR2_X1   g142(.A(new_n327), .B(new_n328), .Z(new_n329));
  INV_X1    g143(.A(KEYINPUT94), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n317), .A2(new_n319), .A3(KEYINPUT16), .ZN(new_n331));
  OR3_X1    g145(.A1(new_n318), .A2(KEYINPUT16), .A3(G140), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n331), .A2(new_n332), .A3(G146), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(G146), .B1(new_n331), .B2(new_n332), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n330), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n331), .A2(new_n332), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(new_n210), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n338), .A2(KEYINPUT94), .A3(new_n333), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  XNOR2_X1  g154(.A(KEYINPUT65), .B(G131), .ZN(new_n341));
  OAI211_X1 g155(.A(KEYINPUT17), .B(new_n341), .C1(new_n313), .C2(new_n314), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n341), .B1(new_n313), .B2(new_n314), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n214), .A2(new_n308), .A3(new_n309), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n342), .B1(new_n345), .B2(KEYINPUT17), .ZN(new_n346));
  OAI211_X1 g160(.A(new_n326), .B(new_n329), .C1(new_n340), .C2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n329), .ZN(new_n348));
  AND3_X1   g162(.A1(new_n317), .A2(new_n319), .A3(KEYINPUT19), .ZN(new_n349));
  AOI21_X1  g163(.A(KEYINPUT19), .B1(new_n317), .B2(new_n319), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n210), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  AND3_X1   g165(.A1(new_n345), .A2(new_n333), .A3(new_n351), .ZN(new_n352));
  AOI22_X1  g166(.A1(new_n321), .A2(new_n323), .B1(G146), .B2(new_n320), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n315), .A2(new_n311), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n348), .B1(new_n352), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n347), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT95), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n347), .A2(new_n356), .A3(KEYINPUT95), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n304), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT20), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n301), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  AND3_X1   g177(.A1(new_n347), .A2(KEYINPUT95), .A3(new_n356), .ZN(new_n364));
  AOI21_X1  g178(.A(KEYINPUT95), .B1(new_n347), .B2(new_n356), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n302), .B(new_n303), .C1(new_n364), .C2(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n366), .A2(KEYINPUT96), .A3(KEYINPUT20), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n304), .A2(KEYINPUT20), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n357), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n363), .A2(new_n367), .A3(new_n369), .ZN(new_n370));
  OR2_X1    g184(.A1(new_n340), .A2(new_n346), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n329), .B1(new_n371), .B2(new_n326), .ZN(new_n372));
  INV_X1    g186(.A(new_n347), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n303), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(G475), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n208), .A2(G128), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n231), .A2(G143), .ZN(new_n377));
  AND2_X1   g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n378), .B(new_n215), .ZN(new_n379));
  INV_X1    g193(.A(G122), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(G116), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n191), .A2(G122), .ZN(new_n382));
  AND2_X1   g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(G107), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OR2_X1    g199(.A1(new_n382), .A2(KEYINPUT14), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n382), .A2(KEYINPUT14), .ZN(new_n387));
  AND3_X1   g201(.A1(new_n386), .A2(new_n381), .A3(new_n387), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n379), .B(new_n385), .C1(new_n384), .C2(new_n388), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n383), .B(new_n384), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT13), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n376), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(new_n377), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n376), .A2(new_n391), .ZN(new_n394));
  OAI21_X1  g208(.A(G134), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n378), .A2(new_n215), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n390), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  XNOR2_X1  g211(.A(KEYINPUT9), .B(G234), .ZN(new_n398));
  INV_X1    g212(.A(G217), .ZN(new_n399));
  NOR3_X1   g213(.A1(new_n398), .A2(new_n399), .A3(G953), .ZN(new_n400));
  AND3_X1   g214(.A1(new_n389), .A2(new_n397), .A3(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n400), .B1(new_n389), .B2(new_n397), .ZN(new_n402));
  OR2_X1    g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(G478), .ZN(new_n404));
  OAI211_X1 g218(.A(new_n403), .B(new_n269), .C1(KEYINPUT15), .C2(new_n404), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n404), .A2(KEYINPUT15), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n401), .A2(new_n402), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n406), .B1(new_n407), .B2(new_n270), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n405), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(G952), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n411), .A2(G953), .ZN(new_n412));
  INV_X1    g226(.A(G234), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n412), .B1(new_n413), .B2(new_n305), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  AOI211_X1 g229(.A(new_n306), .B(new_n269), .C1(G234), .C2(G237), .ZN(new_n416));
  XNOR2_X1  g230(.A(KEYINPUT21), .B(G898), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n370), .A2(new_n375), .A3(new_n410), .A4(new_n419), .ZN(new_n420));
  OAI21_X1  g234(.A(G210), .B1(G237), .B2(G902), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n198), .A2(KEYINPUT5), .A3(new_n189), .A4(new_n192), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(KEYINPUT88), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT5), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n425), .A2(new_n188), .A3(G116), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(G113), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT89), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n427), .B(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT88), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n193), .A2(new_n430), .A3(KEYINPUT5), .A4(new_n198), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n424), .A2(new_n429), .A3(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(G104), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n433), .A2(G107), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n384), .A2(G104), .ZN(new_n435));
  OAI21_X1  g249(.A(G101), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g250(.A(KEYINPUT3), .B1(new_n433), .B2(G107), .ZN(new_n437));
  AOI21_X1  g251(.A(G101), .B1(new_n433), .B2(G107), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT3), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n439), .A2(new_n384), .A3(G104), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n437), .A2(new_n438), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n436), .A2(new_n441), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n200), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n432), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n423), .A2(G113), .A3(new_n426), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n199), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(new_n442), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  XNOR2_X1  g262(.A(G110), .B(G122), .ZN(new_n449));
  XOR2_X1   g263(.A(new_n449), .B(KEYINPUT8), .Z(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n448), .A2(new_n451), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n243), .A2(new_n245), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT90), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n453), .A2(new_n454), .A3(new_n318), .ZN(new_n455));
  OAI21_X1  g269(.A(KEYINPUT90), .B1(new_n236), .B2(G125), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n207), .A2(new_n212), .A3(G125), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(G224), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n459), .A2(G953), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(KEYINPUT7), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n458), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n457), .A2(KEYINPUT87), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n453), .A2(new_n318), .ZN(new_n465));
  INV_X1    g279(.A(new_n462), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT87), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n207), .A2(new_n212), .A3(new_n467), .A4(G125), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n464), .A2(new_n465), .A3(new_n466), .A4(new_n468), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n452), .A2(KEYINPUT91), .A3(new_n463), .A4(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT91), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n463), .A2(new_n469), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n450), .B1(new_n444), .B2(new_n447), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n433), .A2(G107), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n437), .A2(new_n440), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(G101), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n477), .A2(KEYINPUT4), .A3(new_n441), .ZN(new_n478));
  XNOR2_X1  g292(.A(KEYINPUT81), .B(KEYINPUT4), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n476), .A2(G101), .A3(new_n479), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n478), .B(new_n480), .C1(new_n200), .C2(new_n201), .ZN(new_n481));
  AND2_X1   g295(.A1(new_n436), .A2(new_n441), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n445), .A2(new_n199), .A3(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n481), .A2(new_n483), .A3(new_n449), .ZN(new_n484));
  AND3_X1   g298(.A1(new_n470), .A2(new_n474), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n481), .A2(new_n483), .ZN(new_n486));
  INV_X1    g300(.A(new_n449), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT6), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n489), .A2(KEYINPUT86), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n488), .A2(new_n484), .A3(new_n490), .ZN(new_n491));
  OAI211_X1 g305(.A(new_n486), .B(new_n487), .C1(KEYINPUT86), .C2(new_n489), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n464), .A2(new_n465), .A3(new_n468), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n493), .B(new_n460), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n491), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n303), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n422), .B1(new_n485), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n470), .A2(new_n474), .A3(new_n484), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n498), .A2(new_n303), .A3(new_n495), .A4(new_n421), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(G214), .B1(G237), .B2(G902), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(G469), .ZN(new_n503));
  OR2_X1    g317(.A1(new_n223), .A2(new_n226), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT83), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n442), .A2(new_n505), .A3(new_n235), .A4(new_n232), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n441), .B(new_n436), .C1(new_n243), .C2(new_n245), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n505), .B1(new_n453), .B2(new_n442), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n504), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  XNOR2_X1  g324(.A(KEYINPUT84), .B(KEYINPUT12), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  XNOR2_X1  g326(.A(G110), .B(G140), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n306), .A2(G227), .ZN(new_n514));
  XOR2_X1   g328(.A(new_n513), .B(new_n514), .Z(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n246), .A2(KEYINPUT10), .A3(new_n247), .A4(new_n482), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n478), .A2(new_n213), .A3(new_n480), .ZN(new_n518));
  XNOR2_X1  g332(.A(KEYINPUT82), .B(KEYINPUT10), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n507), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n223), .A2(new_n226), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n517), .A2(new_n518), .A3(new_n520), .A4(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT84), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n523), .A2(KEYINPUT12), .ZN(new_n524));
  OAI211_X1 g338(.A(new_n504), .B(new_n524), .C1(new_n508), .C2(new_n509), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n512), .A2(new_n516), .A3(new_n522), .A4(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n517), .A2(new_n518), .A3(new_n520), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(new_n504), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n516), .B1(new_n528), .B2(new_n522), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n526), .B1(new_n529), .B2(KEYINPUT85), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT85), .ZN(new_n531));
  AOI211_X1 g345(.A(new_n531), .B(new_n516), .C1(new_n528), .C2(new_n522), .ZN(new_n532));
  OAI211_X1 g346(.A(new_n503), .B(new_n269), .C1(new_n530), .C2(new_n532), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n503), .A2(new_n303), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n512), .A2(new_n522), .A3(new_n525), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(new_n515), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n528), .A2(new_n516), .A3(new_n522), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n537), .A2(G469), .A3(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n533), .A2(new_n535), .A3(new_n539), .ZN(new_n540));
  OAI21_X1  g354(.A(G221), .B1(new_n398), .B2(G902), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NOR3_X1   g356(.A1(new_n420), .A2(new_n502), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n399), .B1(new_n269), .B2(G234), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT79), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n545), .A2(KEYINPUT25), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n306), .A2(G221), .A3(G234), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n548), .B(KEYINPUT77), .ZN(new_n549));
  XNOR2_X1  g363(.A(KEYINPUT22), .B(G137), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n549), .B(new_n550), .ZN(new_n551));
  OAI21_X1  g365(.A(KEYINPUT74), .B1(new_n188), .B2(G128), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(KEYINPUT23), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT23), .ZN(new_n554));
  OAI211_X1 g368(.A(KEYINPUT74), .B(new_n554), .C1(new_n188), .C2(G128), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n188), .A2(G128), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n553), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(KEYINPUT75), .B1(new_n557), .B2(G110), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n557), .A2(KEYINPUT75), .A3(G110), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  OR3_X1    g375(.A1(new_n231), .A2(KEYINPUT73), .A3(G119), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n556), .A2(KEYINPUT73), .ZN(new_n563));
  AOI22_X1  g377(.A1(new_n562), .A2(new_n563), .B1(G119), .B2(new_n231), .ZN(new_n564));
  XOR2_X1   g378(.A(KEYINPUT24), .B(G110), .Z(new_n565));
  AOI22_X1  g379(.A1(new_n338), .A2(new_n333), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  OAI22_X1  g380(.A1(new_n564), .A2(new_n565), .B1(new_n557), .B2(G110), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n334), .B1(new_n323), .B2(new_n321), .ZN(new_n568));
  AOI22_X1  g382(.A1(new_n561), .A2(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT78), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n551), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  AND3_X1   g385(.A1(new_n557), .A2(KEYINPUT75), .A3(G110), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n566), .B1(new_n558), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n568), .A2(new_n567), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(KEYINPUT78), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n573), .A2(new_n574), .A3(new_n570), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n571), .B1(new_n578), .B2(new_n551), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n547), .B1(new_n579), .B2(new_n269), .ZN(new_n580));
  AND3_X1   g394(.A1(new_n573), .A2(new_n574), .A3(new_n570), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n570), .B1(new_n573), .B2(new_n574), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n551), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n551), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n577), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n583), .A2(new_n269), .A3(new_n585), .A4(new_n547), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n544), .B1(new_n580), .B2(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n544), .A2(G902), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n589), .B(KEYINPUT80), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n579), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n588), .A2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n300), .A2(new_n543), .A3(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n595), .B(G101), .ZN(G3));
  OAI21_X1  g410(.A(new_n269), .B1(new_n296), .B2(new_n297), .ZN(new_n597));
  AOI22_X1  g411(.A1(new_n597), .A2(G472), .B1(new_n293), .B2(new_n294), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n593), .A2(new_n542), .ZN(new_n599));
  AND2_X1   g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n370), .A2(new_n375), .ZN(new_n601));
  XNOR2_X1  g415(.A(KEYINPUT97), .B(KEYINPUT33), .ZN(new_n602));
  OR3_X1    g416(.A1(new_n401), .A2(new_n402), .A3(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT33), .ZN(new_n604));
  OAI22_X1  g418(.A1(new_n401), .A2(new_n402), .B1(KEYINPUT97), .B2(new_n604), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n603), .A2(G478), .A3(new_n269), .A4(new_n605), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n404), .B1(new_n407), .B2(new_n270), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n601), .A2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n501), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n610), .B1(new_n497), .B2(new_n499), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(new_n419), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n600), .A2(new_n613), .ZN(new_n614));
  XOR2_X1   g428(.A(KEYINPUT34), .B(G104), .Z(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(G6));
  NAND2_X1  g430(.A1(new_n359), .A2(new_n360), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(new_n368), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n363), .A2(new_n367), .A3(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n619), .A2(new_n375), .A3(new_n409), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n612), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n600), .A2(new_n621), .ZN(new_n622));
  XOR2_X1   g436(.A(KEYINPUT35), .B(G107), .Z(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(G9));
  NOR2_X1   g438(.A1(new_n420), .A2(new_n542), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n584), .A2(KEYINPUT36), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(new_n575), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(new_n591), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n588), .A2(KEYINPUT98), .A3(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT98), .ZN(new_n630));
  INV_X1    g444(.A(new_n544), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n583), .A2(new_n269), .A3(new_n585), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(new_n546), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n631), .B1(new_n633), .B2(new_n586), .ZN(new_n634));
  INV_X1    g448(.A(new_n628), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n630), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n629), .A2(new_n636), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n598), .A2(new_n611), .A3(new_n625), .A4(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT37), .B(G110), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G12));
  INV_X1    g454(.A(new_n542), .ZN(new_n641));
  AND3_X1   g455(.A1(new_n637), .A2(new_n611), .A3(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(G900), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n415), .B1(new_n416), .B2(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n620), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n300), .A2(new_n642), .A3(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(G128), .ZN(G30));
  OAI21_X1  g461(.A(new_n294), .B1(new_n296), .B2(new_n297), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(KEYINPUT32), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n298), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n250), .A2(new_n280), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n257), .B1(new_n272), .B2(new_n251), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n303), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(G472), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n650), .A2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n637), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n658), .A2(new_n501), .A3(new_n601), .A4(new_n409), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n657), .B1(KEYINPUT99), .B2(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(KEYINPUT100), .B(KEYINPUT39), .ZN(new_n661));
  XOR2_X1   g475(.A(new_n644), .B(new_n661), .Z(new_n662));
  NOR2_X1   g476(.A1(new_n542), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(KEYINPUT40), .ZN(new_n664));
  OR2_X1    g478(.A1(new_n659), .A2(KEYINPUT99), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n500), .B(KEYINPUT38), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n660), .A2(new_n664), .A3(new_n665), .A4(new_n666), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT101), .B(G143), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G45));
  INV_X1    g483(.A(new_n608), .ZN(new_n670));
  AOI211_X1 g484(.A(new_n644), .B(new_n670), .C1(new_n370), .C2(new_n375), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n300), .A2(new_n642), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G146), .ZN(G48));
  OAI21_X1  g487(.A(new_n269), .B1(new_n530), .B2(new_n532), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(G469), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n675), .A2(new_n541), .A3(new_n533), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n300), .A2(new_n594), .A3(new_n613), .A4(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(KEYINPUT41), .B(G113), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G15));
  NAND4_X1  g494(.A1(new_n300), .A2(new_n594), .A3(new_n621), .A4(new_n677), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G116), .ZN(G18));
  INV_X1    g496(.A(KEYINPUT102), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n683), .B1(new_n502), .B2(new_n676), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n677), .A2(KEYINPUT102), .A3(new_n611), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n420), .B1(new_n636), .B2(new_n629), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n300), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G119), .ZN(G21));
  NAND4_X1  g503(.A1(new_n601), .A2(new_n501), .A3(new_n500), .A4(new_n409), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n294), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n273), .A2(new_n257), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n693), .A2(new_n287), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n692), .B1(new_n694), .B2(new_n285), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n695), .B1(new_n597), .B2(G472), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n676), .A2(new_n418), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n691), .A2(new_n696), .A3(new_n594), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G122), .ZN(G24));
  AND3_X1   g513(.A1(new_n696), .A2(new_n637), .A3(new_n671), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(new_n686), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G125), .ZN(G27));
  AND3_X1   g516(.A1(new_n497), .A2(new_n499), .A3(new_n501), .ZN(new_n703));
  OR2_X1    g517(.A1(new_n538), .A2(KEYINPUT103), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n538), .A2(KEYINPUT103), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n704), .A2(new_n537), .A3(G469), .A4(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n533), .A2(new_n535), .A3(new_n706), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n703), .A2(KEYINPUT104), .A3(new_n541), .A4(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT104), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n707), .A2(new_n541), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n497), .A2(new_n499), .A3(new_n501), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n709), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n708), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n300), .A2(new_n594), .A3(new_n671), .A4(new_n713), .ZN(new_n714));
  XOR2_X1   g528(.A(KEYINPUT105), .B(KEYINPUT42), .Z(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(new_n644), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n601), .A2(new_n608), .A3(KEYINPUT42), .A4(new_n717), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n718), .B1(new_n708), .B2(new_n712), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n649), .A2(KEYINPUT106), .A3(new_n298), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(new_n277), .ZN(new_n721));
  AOI21_X1  g535(.A(KEYINPUT106), .B1(new_n649), .B2(new_n298), .ZN(new_n722));
  OAI211_X1 g536(.A(new_n594), .B(new_n719), .C1(new_n721), .C2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n716), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G131), .ZN(G33));
  NAND4_X1  g539(.A1(new_n300), .A2(new_n594), .A3(new_n645), .A4(new_n713), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G134), .ZN(G36));
  INV_X1    g541(.A(new_n541), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n704), .A2(KEYINPUT45), .A3(new_n537), .A4(new_n705), .ZN(new_n729));
  AND2_X1   g543(.A1(new_n537), .A2(new_n538), .ZN(new_n730));
  OAI211_X1 g544(.A(new_n729), .B(G469), .C1(KEYINPUT45), .C2(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n731), .A2(KEYINPUT46), .A3(new_n535), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n533), .ZN(new_n733));
  OR2_X1    g547(.A1(new_n733), .A2(KEYINPUT107), .ZN(new_n734));
  AOI21_X1  g548(.A(KEYINPUT46), .B1(new_n731), .B2(new_n535), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n735), .B1(new_n733), .B2(KEYINPUT107), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n728), .B1(new_n734), .B2(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(new_n662), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  OR2_X1    g553(.A1(new_n598), .A2(new_n658), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n370), .A2(new_n375), .A3(new_n608), .ZN(new_n741));
  OR2_X1    g555(.A1(new_n741), .A2(KEYINPUT43), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(KEYINPUT43), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n740), .A2(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT108), .ZN(new_n746));
  OR3_X1    g560(.A1(new_n745), .A2(new_n746), .A3(KEYINPUT44), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n746), .B1(new_n745), .B2(KEYINPUT44), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n711), .B1(new_n745), .B2(KEYINPUT44), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n747), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n739), .B1(new_n750), .B2(KEYINPUT109), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n751), .B1(KEYINPUT109), .B2(new_n750), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G137), .ZN(G39));
  OR2_X1    g567(.A1(new_n737), .A2(KEYINPUT47), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n737), .A2(KEYINPUT47), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT72), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n276), .B(new_n757), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n758), .B1(new_n649), .B2(new_n298), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n594), .A2(new_n711), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n756), .A2(new_n759), .A3(new_n671), .A4(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G140), .ZN(G42));
  OR4_X1    g576(.A1(new_n593), .A2(new_n666), .A3(new_n610), .A4(new_n728), .ZN(new_n763));
  AND2_X1   g577(.A1(new_n675), .A2(new_n533), .ZN(new_n764));
  XOR2_X1   g578(.A(new_n764), .B(KEYINPUT49), .Z(new_n765));
  OR4_X1    g579(.A1(new_n656), .A2(new_n763), .A3(new_n741), .A4(new_n765), .ZN(new_n766));
  OAI211_X1 g580(.A(new_n300), .B(new_n642), .C1(new_n645), .C2(new_n671), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n588), .A2(new_n628), .A3(new_n717), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n690), .A2(new_n710), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n656), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n767), .A2(new_n701), .A3(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(KEYINPUT52), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n678), .A2(new_n681), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n595), .A2(new_n688), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n609), .B1(new_n601), .B2(new_n410), .ZN(new_n775));
  INV_X1    g589(.A(new_n612), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n775), .A2(new_n598), .A3(new_n776), .A4(new_n599), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n777), .A2(new_n698), .A3(new_n638), .ZN(new_n778));
  NOR3_X1   g592(.A1(new_n773), .A2(new_n774), .A3(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT111), .ZN(new_n780));
  INV_X1    g594(.A(new_n726), .ZN(new_n781));
  INV_X1    g595(.A(new_n713), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n696), .A2(new_n637), .A3(new_n671), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n542), .A2(new_n711), .ZN(new_n784));
  AND4_X1   g598(.A1(new_n375), .A2(new_n408), .A3(new_n405), .A4(new_n717), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n619), .A2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT110), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n619), .A2(new_n785), .A3(KEYINPUT110), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n637), .A2(new_n784), .A3(new_n788), .A4(new_n789), .ZN(new_n790));
  OAI22_X1  g604(.A1(new_n782), .A2(new_n783), .B1(new_n759), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n780), .B1(new_n781), .B2(new_n791), .ZN(new_n792));
  AND4_X1   g606(.A1(new_n637), .A2(new_n784), .A3(new_n789), .A4(new_n788), .ZN(new_n793));
  AOI22_X1  g607(.A1(new_n700), .A2(new_n713), .B1(new_n793), .B2(new_n300), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n794), .A2(KEYINPUT111), .A3(new_n726), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n779), .A2(new_n724), .A3(new_n792), .A4(new_n795), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n772), .B1(new_n796), .B2(KEYINPUT112), .ZN(new_n797));
  AOI21_X1  g611(.A(KEYINPUT111), .B1(new_n794), .B2(new_n726), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n713), .A2(new_n637), .A3(new_n671), .A4(new_n696), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n793), .A2(new_n300), .ZN(new_n800));
  AND4_X1   g614(.A1(KEYINPUT111), .A2(new_n726), .A3(new_n799), .A4(new_n800), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT112), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n802), .A2(new_n803), .A3(new_n724), .A4(new_n779), .ZN(new_n804));
  AOI21_X1  g618(.A(KEYINPUT53), .B1(new_n797), .B2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT53), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n796), .A2(new_n772), .A3(new_n806), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n805), .A2(KEYINPUT54), .A3(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT54), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n774), .A2(new_n778), .ZN(new_n810));
  INV_X1    g624(.A(new_n773), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n810), .A2(new_n724), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n792), .A2(new_n795), .ZN(new_n813));
  OAI21_X1  g627(.A(KEYINPUT112), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(new_n772), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n804), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(new_n806), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n797), .A2(KEYINPUT53), .A3(new_n804), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n809), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n808), .A2(new_n819), .A3(KEYINPUT113), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT113), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n816), .A2(new_n806), .ZN(new_n822));
  OAI21_X1  g636(.A(KEYINPUT54), .B1(new_n822), .B2(new_n805), .ZN(new_n823));
  INV_X1    g637(.A(new_n807), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n817), .A2(new_n809), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n821), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n820), .A2(new_n826), .ZN(new_n827));
  OR2_X1    g641(.A1(new_n721), .A2(new_n722), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n742), .A2(new_n415), .A3(new_n743), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n829), .A2(new_n676), .A3(new_n711), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n828), .A2(new_n594), .A3(new_n830), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(KEYINPUT48), .ZN(new_n832));
  NOR4_X1   g646(.A1(new_n593), .A2(new_n676), .A3(new_n711), .A4(new_n414), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n657), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n412), .B1(new_n834), .B2(new_n609), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n696), .A2(new_n594), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n829), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n835), .B1(new_n686), .B2(new_n837), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n764), .A2(new_n728), .ZN(new_n839));
  OAI211_X1 g653(.A(new_n703), .B(new_n837), .C1(new_n756), .C2(new_n839), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n834), .A2(new_n601), .A3(new_n608), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n696), .A2(new_n637), .ZN(new_n842));
  INV_X1    g656(.A(new_n842), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n841), .B1(new_n843), .B2(new_n830), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n840), .A2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT50), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n666), .B1(KEYINPUT115), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n677), .A2(new_n610), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(KEYINPUT114), .ZN(new_n849));
  OR2_X1    g663(.A1(new_n848), .A2(KEYINPUT114), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n847), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(new_n837), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n846), .A2(KEYINPUT115), .ZN(new_n853));
  OR2_X1    g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n852), .A2(new_n853), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n854), .A2(KEYINPUT51), .A3(new_n855), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n832), .B(new_n838), .C1(new_n845), .C2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(new_n855), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n852), .A2(new_n853), .ZN(new_n859));
  OAI21_X1  g673(.A(KEYINPUT116), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT116), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n854), .A2(new_n861), .A3(new_n855), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n860), .A2(new_n862), .A3(new_n840), .A4(new_n844), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT51), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(KEYINPUT117), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT117), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n863), .A2(new_n867), .A3(new_n864), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n857), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(KEYINPUT118), .B1(new_n827), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g684(.A(KEYINPUT113), .B1(new_n808), .B2(new_n819), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n823), .A2(new_n821), .A3(new_n825), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n871), .A2(new_n872), .A3(new_n869), .A4(KEYINPUT118), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n411), .A2(new_n306), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n766), .B1(new_n870), .B2(new_n875), .ZN(G75));
  NOR2_X1   g690(.A1(new_n306), .A2(G952), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT56), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n491), .A2(new_n492), .ZN(new_n880));
  XOR2_X1   g694(.A(new_n880), .B(new_n494), .Z(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(KEYINPUT55), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n817), .A2(new_n824), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n883), .A2(new_n270), .A3(new_n422), .ZN(new_n884));
  OAI211_X1 g698(.A(new_n879), .B(new_n882), .C1(new_n884), .C2(KEYINPUT120), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n884), .A2(KEYINPUT120), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n878), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT119), .ZN(new_n888));
  OR2_X1    g702(.A1(new_n884), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(KEYINPUT56), .B1(new_n884), .B2(new_n888), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n882), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n887), .A2(new_n891), .ZN(G51));
  OAI21_X1  g706(.A(KEYINPUT54), .B1(new_n805), .B2(new_n807), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n893), .A2(KEYINPUT121), .A3(new_n825), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT121), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n883), .A2(new_n895), .A3(KEYINPUT54), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n534), .B(KEYINPUT57), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n894), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT122), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  OR2_X1    g714(.A1(new_n530), .A2(new_n532), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n894), .A2(KEYINPUT122), .A3(new_n896), .A4(new_n897), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(new_n883), .ZN(new_n904));
  OR3_X1    g718(.A1(new_n904), .A2(new_n269), .A3(new_n731), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n877), .B1(new_n903), .B2(new_n905), .ZN(G54));
  NAND4_X1  g720(.A1(new_n883), .A2(KEYINPUT58), .A3(G475), .A4(new_n270), .ZN(new_n907));
  INV_X1    g721(.A(new_n617), .ZN(new_n908));
  AND2_X1   g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n907), .A2(new_n908), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n909), .A2(new_n910), .A3(new_n877), .ZN(G60));
  NAND2_X1  g725(.A1(new_n603), .A2(new_n605), .ZN(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(G478), .A2(G902), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(KEYINPUT59), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n894), .A2(new_n913), .A3(new_n896), .A4(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(new_n878), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n915), .B1(new_n820), .B2(new_n826), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n917), .B1(new_n912), .B2(new_n918), .ZN(G63));
  NAND2_X1  g733(.A1(G217), .A2(G902), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(KEYINPUT60), .ZN(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n883), .A2(new_n627), .A3(new_n922), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n904), .A2(new_n921), .ZN(new_n924));
  OAI211_X1 g738(.A(new_n878), .B(new_n923), .C1(new_n924), .C2(new_n579), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n923), .A2(KEYINPUT123), .A3(new_n878), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(KEYINPUT61), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n925), .B(new_n927), .ZN(G66));
  NOR3_X1   g742(.A1(new_n417), .A2(new_n459), .A3(new_n306), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n929), .B1(new_n779), .B2(new_n306), .ZN(new_n930));
  INV_X1    g744(.A(G898), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n880), .B1(new_n931), .B2(G953), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n930), .B(new_n932), .Z(G69));
  NOR2_X1   g747(.A1(new_n241), .A2(new_n249), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n349), .A2(new_n350), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n934), .B(new_n935), .Z(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(G227), .Z(new_n937));
  NOR3_X1   g751(.A1(new_n937), .A2(new_n643), .A3(new_n306), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n759), .A2(new_n593), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n939), .A2(new_n738), .A3(new_n775), .A4(new_n784), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n752), .A2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT125), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n752), .A2(KEYINPUT125), .A3(new_n940), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  AND2_X1   g759(.A1(new_n767), .A2(new_n701), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n667), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n947), .B1(KEYINPUT124), .B2(KEYINPUT62), .ZN(new_n948));
  XNOR2_X1  g762(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n948), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n945), .A2(new_n761), .A3(new_n936), .A4(new_n950), .ZN(new_n951));
  AND2_X1   g765(.A1(new_n946), .A2(new_n726), .ZN(new_n952));
  INV_X1    g766(.A(new_n739), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n953), .A2(new_n594), .A3(new_n691), .A4(new_n828), .ZN(new_n954));
  AND4_X1   g768(.A1(new_n724), .A2(new_n761), .A3(new_n952), .A4(new_n954), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n752), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n951), .B1(new_n956), .B2(new_n936), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n938), .B1(new_n957), .B2(new_n306), .ZN(G72));
  XOR2_X1   g772(.A(new_n252), .B(KEYINPUT126), .Z(new_n959));
  NOR2_X1   g773(.A1(new_n959), .A2(new_n258), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n950), .A2(new_n761), .A3(new_n779), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n961), .B1(new_n943), .B2(new_n944), .ZN(new_n962));
  NAND2_X1  g776(.A1(G472), .A2(G902), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT63), .Z(new_n964));
  INV_X1    g778(.A(new_n964), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n960), .B1(new_n962), .B2(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n965), .B1(new_n259), .B2(new_n651), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n967), .B1(new_n822), .B2(new_n805), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n959), .A2(new_n258), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n956), .A2(new_n779), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n970), .B1(new_n971), .B2(new_n964), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT127), .ZN(new_n973));
  OR3_X1    g787(.A1(new_n972), .A2(new_n973), .A3(new_n877), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n973), .B1(new_n972), .B2(new_n877), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n969), .B1(new_n974), .B2(new_n975), .ZN(G57));
endmodule


