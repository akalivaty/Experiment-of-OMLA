//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 1 0 0 1 1 0 1 1 1 0 0 0 1 0 0 0 1 0 1 0 0 1 1 1 1 1 1 1 1 0 0 1 0 1 0 0 0 0 0 1 0 0 1 0 1 0 0 1 1 0 0 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:24 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n448, new_n450, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n549,
    new_n551, new_n552, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n611, new_n612, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1118,
    new_n1119;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT64), .B(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT65), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  NAND2_X1  g022(.A1(G94), .A2(G452), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT66), .ZN(G173));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g026(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n454));
  XNOR2_X1  g029(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n454), .B(new_n455), .ZN(new_n456));
  OR4_X1    g031(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n456), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n456), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  AOI22_X1  g036(.A1(new_n461), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n462));
  XOR2_X1   g037(.A(KEYINPUT68), .B(G2105), .Z(new_n463));
  NOR2_X1   g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n465), .A2(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G101), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT68), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n471));
  AND2_X1   g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  NOR2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  OAI211_X1 g048(.A(new_n470), .B(new_n471), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G137), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n467), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n464), .A2(new_n476), .ZN(new_n477));
  XNOR2_X1  g052(.A(new_n477), .B(KEYINPUT69), .ZN(G160));
  NAND2_X1  g053(.A1(new_n470), .A2(new_n471), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(new_n461), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n461), .A2(new_n469), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  AOI22_X1  g058(.A1(G124), .A2(new_n481), .B1(new_n483), .B2(G136), .ZN(new_n484));
  OAI221_X1 g059(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n463), .C2(G112), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  XOR2_X1   g061(.A(new_n486), .B(KEYINPUT70), .Z(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  NAND2_X1  g063(.A1(G114), .A2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(G102), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n489), .B1(new_n490), .B2(G2105), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G2104), .ZN(new_n492));
  AND2_X1   g067(.A1(G126), .A2(G2105), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n493), .B1(new_n472), .B2(new_n473), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT71), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT71), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n492), .A2(new_n497), .A3(new_n494), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(G138), .ZN(new_n500));
  OAI21_X1  g075(.A(KEYINPUT4), .B1(new_n474), .B2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n463), .A2(new_n461), .A3(new_n502), .A4(G138), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n499), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(G164));
  AND2_X1   g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  OR2_X1    g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(KEYINPUT72), .A2(KEYINPUT5), .ZN(new_n510));
  INV_X1    g085(.A(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g087(.A1(KEYINPUT72), .A2(KEYINPUT5), .A3(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n509), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G88), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n509), .A2(G543), .ZN(new_n517));
  INV_X1    g092(.A(G50), .ZN(new_n518));
  OAI22_X1  g093(.A1(new_n515), .A2(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n514), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n520));
  INV_X1    g095(.A(G651), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n519), .A2(new_n522), .ZN(G166));
  INV_X1    g098(.A(new_n515), .ZN(new_n524));
  AND2_X1   g099(.A1(new_n524), .A2(G89), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n526), .B(KEYINPUT7), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n514), .A2(G63), .A3(G651), .ZN(new_n528));
  INV_X1    g103(.A(G51), .ZN(new_n529));
  OAI211_X1 g104(.A(new_n527), .B(new_n528), .C1(new_n517), .C2(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n525), .A2(new_n530), .ZN(G168));
  INV_X1    g106(.A(G90), .ZN(new_n532));
  INV_X1    g107(.A(G52), .ZN(new_n533));
  OAI22_X1  g108(.A1(new_n515), .A2(new_n532), .B1(new_n517), .B2(new_n533), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n514), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n535), .A2(new_n521), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n534), .A2(new_n536), .ZN(G171));
  NAND2_X1  g112(.A1(new_n514), .A2(G56), .ZN(new_n538));
  INV_X1    g113(.A(G68), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n539), .B2(new_n511), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT73), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n521), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n542), .B1(new_n541), .B2(new_n540), .ZN(new_n543));
  INV_X1    g118(.A(new_n517), .ZN(new_n544));
  AOI22_X1  g119(.A1(G81), .A2(new_n524), .B1(new_n544), .B2(G43), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  AND3_X1   g123(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G36), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n549), .A2(new_n552), .ZN(G188));
  INV_X1    g128(.A(KEYINPUT9), .ZN(new_n554));
  OAI211_X1 g129(.A(G53), .B(G543), .C1(new_n507), .C2(new_n508), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(KEYINPUT74), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT74), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g134(.A(new_n554), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(KEYINPUT75), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT75), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n562), .B1(new_n556), .B2(new_n554), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n561), .B1(new_n560), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(G78), .A2(G543), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT76), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n514), .B(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(G65), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n565), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n569), .A2(G651), .B1(G91), .B2(new_n524), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n564), .A2(new_n570), .ZN(G299));
  INV_X1    g146(.A(G171), .ZN(G301));
  INV_X1    g147(.A(G168), .ZN(G286));
  INV_X1    g148(.A(G166), .ZN(G303));
  NAND2_X1  g149(.A1(new_n524), .A2(G87), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n544), .A2(G49), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(G288));
  INV_X1    g153(.A(G86), .ZN(new_n579));
  INV_X1    g154(.A(G48), .ZN(new_n580));
  OAI22_X1  g155(.A1(new_n515), .A2(new_n579), .B1(new_n517), .B2(new_n580), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n514), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n582), .A2(new_n521), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(G305));
  INV_X1    g160(.A(G85), .ZN(new_n586));
  INV_X1    g161(.A(G47), .ZN(new_n587));
  OAI22_X1  g162(.A1(new_n515), .A2(new_n586), .B1(new_n517), .B2(new_n587), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n589), .A2(new_n521), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(G290));
  INV_X1    g167(.A(G66), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n567), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(G79), .A2(G543), .ZN(new_n595));
  XOR2_X1   g170(.A(new_n595), .B(KEYINPUT77), .Z(new_n596));
  OAI21_X1  g171(.A(G651), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n524), .A2(KEYINPUT10), .A3(G92), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT10), .ZN(new_n599));
  INV_X1    g174(.A(G92), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n515), .B2(new_n600), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n598), .A2(new_n601), .B1(G54), .B2(new_n544), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n597), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(G868), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(G171), .A2(G868), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(G284));
  XNOR2_X1  g184(.A(new_n608), .B(KEYINPUT78), .ZN(G321));
  NOR2_X1   g185(.A1(G286), .A2(new_n605), .ZN(new_n611));
  INV_X1    g186(.A(G299), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n611), .B1(new_n612), .B2(new_n605), .ZN(G297));
  AOI21_X1  g188(.A(new_n611), .B1(new_n612), .B2(new_n605), .ZN(G280));
  XNOR2_X1  g189(.A(KEYINPUT79), .B(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n604), .B1(G860), .B2(new_n615), .ZN(G148));
  NAND2_X1  g191(.A1(new_n547), .A2(new_n605), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n604), .A2(new_n615), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(new_n605), .ZN(new_n619));
  XNOR2_X1  g194(.A(KEYINPUT80), .B(KEYINPUT11), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n619), .B(new_n620), .ZN(G282));
  INV_X1    g196(.A(new_n619), .ZN(G323));
  AOI22_X1  g197(.A1(G123), .A2(new_n481), .B1(new_n483), .B2(G135), .ZN(new_n623));
  OAI221_X1 g198(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n463), .C2(G111), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT82), .ZN(new_n626));
  INV_X1    g201(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(G2096), .ZN(new_n628));
  INV_X1    g203(.A(G2096), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n482), .A2(new_n465), .ZN(new_n631));
  XOR2_X1   g206(.A(KEYINPUT81), .B(KEYINPUT12), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT13), .B(G2100), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n628), .A2(new_n630), .A3(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(KEYINPUT83), .Z(G156));
  XOR2_X1   g212(.A(G2451), .B(G2454), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT16), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT84), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2443), .B(G2446), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G1341), .B(G1348), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(KEYINPUT15), .B(G2435), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2438), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(G2427), .Z(new_n647));
  OAI21_X1  g222(.A(KEYINPUT14), .B1(new_n647), .B2(G2430), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n648), .B1(G2430), .B2(new_n647), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n644), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n644), .A2(new_n649), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n650), .A2(G14), .A3(new_n651), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(G401));
  XNOR2_X1  g228(.A(G2067), .B(G2678), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(KEYINPUT85), .Z(new_n655));
  NOR2_X1   g230(.A1(G2072), .A2(G2078), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n444), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2084), .B(G2090), .Z(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n657), .B(KEYINPUT17), .ZN(new_n661));
  OAI211_X1 g236(.A(new_n658), .B(new_n660), .C1(new_n655), .C2(new_n661), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n661), .A2(new_n655), .A3(new_n659), .ZN(new_n663));
  OAI211_X1 g238(.A(new_n659), .B(new_n654), .C1(new_n444), .C2(new_n656), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(KEYINPUT18), .Z(new_n665));
  NAND3_X1  g240(.A1(new_n662), .A2(new_n663), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(new_n629), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n667), .B(G2100), .Z(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(G227));
  XOR2_X1   g244(.A(G1971), .B(G1976), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT19), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1956), .B(G2474), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1961), .B(G1966), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  AND2_X1   g249(.A1(new_n672), .A2(new_n673), .ZN(new_n675));
  NOR3_X1   g250(.A1(new_n671), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n671), .A2(new_n674), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(KEYINPUT20), .Z(new_n678));
  AOI211_X1 g253(.A(new_n676), .B(new_n678), .C1(new_n671), .C2(new_n675), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1981), .B(G1986), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n679), .B(new_n680), .Z(new_n681));
  XNOR2_X1  g256(.A(G1991), .B(G1996), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT87), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT86), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n683), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n681), .B(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(G229));
  NOR2_X1   g263(.A1(G16), .A2(G24), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n689), .B1(new_n591), .B2(G16), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n690), .B(G1986), .Z(new_n691));
  AOI22_X1  g266(.A1(G119), .A2(new_n481), .B1(new_n483), .B2(G131), .ZN(new_n692));
  OAI221_X1 g267(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n463), .C2(G107), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  MUX2_X1   g269(.A(G25), .B(new_n694), .S(G29), .Z(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT89), .Z(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT35), .B(G1991), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(KEYINPUT88), .Z(new_n698));
  OAI21_X1  g273(.A(new_n691), .B1(new_n696), .B2(new_n698), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n699), .B1(new_n698), .B2(new_n696), .ZN(new_n700));
  NOR2_X1   g275(.A1(G6), .A2(G16), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n701), .B1(new_n584), .B2(G16), .ZN(new_n702));
  XOR2_X1   g277(.A(KEYINPUT32), .B(G1981), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  NOR2_X1   g279(.A1(G16), .A2(G23), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(KEYINPUT90), .Z(new_n706));
  INV_X1    g281(.A(G16), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n706), .B1(G288), .B2(new_n707), .ZN(new_n708));
  XOR2_X1   g283(.A(KEYINPUT33), .B(G1976), .Z(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  NOR2_X1   g285(.A1(G16), .A2(G22), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(G166), .B2(G16), .ZN(new_n712));
  INV_X1    g287(.A(G1971), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n704), .A2(new_n710), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(KEYINPUT34), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n715), .A2(KEYINPUT34), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n700), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(KEYINPUT36), .Z(new_n719));
  INV_X1    g294(.A(G29), .ZN(new_n720));
  AND2_X1   g295(.A1(new_n720), .A2(G33), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT25), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  AND2_X1   g299(.A1(new_n461), .A2(G127), .ZN(new_n725));
  AND2_X1   g300(.A1(G115), .A2(G2104), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n479), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n483), .A2(G139), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n724), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT93), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n721), .B1(new_n730), .B2(G29), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n731), .A2(new_n442), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT94), .Z(new_n733));
  NAND2_X1  g308(.A1(new_n707), .A2(G5), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G171), .B2(new_n707), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(G1961), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n707), .A2(G21), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G168), .B2(new_n707), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(G1966), .ZN(new_n739));
  AOI211_X1 g314(.A(new_n736), .B(new_n739), .C1(new_n731), .C2(new_n442), .ZN(new_n740));
  NAND2_X1  g315(.A1(G160), .A2(G29), .ZN(new_n741));
  AND2_X1   g316(.A1(KEYINPUT24), .A2(G34), .ZN(new_n742));
  NOR2_X1   g317(.A1(KEYINPUT24), .A2(G34), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n720), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n741), .A2(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(G2084), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT96), .ZN(new_n748));
  AOI22_X1  g323(.A1(G129), .A2(new_n481), .B1(new_n483), .B2(G141), .ZN(new_n749));
  NAND3_X1  g324(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT26), .ZN(new_n751));
  OR2_X1    g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n750), .A2(new_n751), .ZN(new_n753));
  AOI22_X1  g328(.A1(new_n752), .A2(new_n753), .B1(G105), .B2(new_n466), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n749), .A2(new_n754), .ZN(new_n755));
  MUX2_X1   g330(.A(G32), .B(new_n755), .S(G29), .Z(new_n756));
  XNOR2_X1  g331(.A(KEYINPUT27), .B(G1996), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(KEYINPUT95), .Z(new_n758));
  XNOR2_X1  g333(.A(new_n756), .B(new_n758), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n745), .A2(new_n746), .ZN(new_n760));
  XOR2_X1   g335(.A(KEYINPUT31), .B(G11), .Z(new_n761));
  XNOR2_X1  g336(.A(KEYINPUT30), .B(G28), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n761), .B1(new_n720), .B2(new_n762), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(new_n627), .B2(new_n720), .ZN(new_n764));
  NOR2_X1   g339(.A1(G27), .A2(G29), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(G164), .B2(G29), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(G2078), .ZN(new_n767));
  NOR4_X1   g342(.A1(new_n759), .A2(new_n760), .A3(new_n764), .A4(new_n767), .ZN(new_n768));
  NAND4_X1  g343(.A1(new_n733), .A2(new_n740), .A3(new_n748), .A4(new_n768), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n769), .A2(KEYINPUT97), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n720), .A2(G35), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G162), .B2(new_n720), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT29), .Z(new_n773));
  INV_X1    g348(.A(G2090), .ZN(new_n774));
  AND2_X1   g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n773), .A2(new_n774), .ZN(new_n776));
  NOR2_X1   g351(.A1(G4), .A2(G16), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT91), .Z(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(new_n603), .B2(new_n707), .ZN(new_n779));
  INV_X1    g354(.A(G1348), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(G16), .A2(G19), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(new_n547), .B2(G16), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(G1341), .Z(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT98), .B(KEYINPUT23), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n707), .A2(G20), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(G299), .B2(G16), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(G1956), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n720), .A2(G26), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(KEYINPUT92), .Z(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT28), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n481), .A2(G128), .ZN(new_n793));
  OAI221_X1 g368(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n463), .C2(G116), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n483), .A2(G140), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n793), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n792), .B1(new_n796), .B2(G29), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(G2067), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n784), .A2(new_n789), .A3(new_n798), .ZN(new_n799));
  NOR4_X1   g374(.A1(new_n775), .A2(new_n776), .A3(new_n781), .A4(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n769), .A2(KEYINPUT97), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n770), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  OR2_X1    g377(.A1(new_n802), .A2(KEYINPUT99), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n802), .A2(KEYINPUT99), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n719), .B1(new_n803), .B2(new_n804), .ZN(G311));
  INV_X1    g380(.A(G311), .ZN(G150));
  AOI22_X1  g381(.A1(G93), .A2(new_n524), .B1(new_n544), .B2(G55), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n807), .A2(KEYINPUT100), .ZN(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n807), .A2(KEYINPUT100), .ZN(new_n810));
  AOI22_X1  g385(.A1(new_n514), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n811));
  OAI22_X1  g386(.A1(new_n809), .A2(new_n810), .B1(new_n521), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n812), .A2(G860), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(KEYINPUT37), .Z(new_n814));
  XNOR2_X1  g389(.A(new_n812), .B(new_n546), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT38), .ZN(new_n816));
  AND2_X1   g391(.A1(new_n604), .A2(G559), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n818), .A2(KEYINPUT39), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT101), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT102), .ZN(new_n821));
  AOI21_X1  g396(.A(G860), .B1(new_n818), .B2(KEYINPUT39), .ZN(new_n822));
  AND3_X1   g397(.A1(new_n820), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n821), .B1(new_n820), .B2(new_n822), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n814), .B1(new_n823), .B2(new_n824), .ZN(G145));
  XOR2_X1   g400(.A(new_n730), .B(new_n755), .Z(new_n826));
  INV_X1    g401(.A(KEYINPUT103), .ZN(new_n827));
  INV_X1    g402(.A(new_n495), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n827), .B1(new_n504), .B2(new_n828), .ZN(new_n829));
  AOI211_X1 g404(.A(KEYINPUT103), .B(new_n495), .C1(new_n501), .C2(new_n503), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  XOR2_X1   g406(.A(new_n831), .B(new_n796), .Z(new_n832));
  OR2_X1    g407(.A1(new_n826), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n826), .A2(new_n832), .ZN(new_n834));
  AOI22_X1  g409(.A1(G130), .A2(new_n481), .B1(new_n483), .B2(G142), .ZN(new_n835));
  OAI221_X1 g410(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n463), .C2(G118), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n694), .B(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(new_n633), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n839), .A2(KEYINPUT104), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n833), .A2(new_n834), .A3(new_n840), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n839), .A2(KEYINPUT104), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n841), .B(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n487), .B(G160), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(new_n627), .ZN(new_n845));
  OR2_X1    g420(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g421(.A(G37), .B1(new_n843), .B2(new_n845), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g424(.A1(new_n812), .A2(new_n605), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT111), .ZN(new_n851));
  XOR2_X1   g426(.A(G166), .B(new_n584), .Z(new_n852));
  XNOR2_X1  g427(.A(G288), .B(new_n591), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n854), .B(KEYINPUT109), .Z(new_n855));
  OR2_X1    g430(.A1(new_n852), .A2(new_n853), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT42), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n857), .A2(KEYINPUT110), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT110), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n861), .B1(new_n855), .B2(new_n856), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n859), .B1(new_n863), .B2(new_n858), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n604), .A2(G299), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT106), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n604), .A2(G299), .A3(KEYINPUT106), .ZN(new_n869));
  AOI22_X1  g444(.A1(new_n868), .A2(new_n869), .B1(new_n612), .B2(new_n603), .ZN(new_n870));
  OR3_X1    g445(.A1(new_n870), .A2(KEYINPUT107), .A3(KEYINPUT41), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(KEYINPUT41), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT108), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n870), .A2(KEYINPUT108), .A3(KEYINPUT41), .ZN(new_n875));
  OAI21_X1  g450(.A(KEYINPUT107), .B1(new_n870), .B2(KEYINPUT41), .ZN(new_n876));
  NAND4_X1  g451(.A1(new_n871), .A2(new_n874), .A3(new_n875), .A4(new_n876), .ZN(new_n877));
  XOR2_X1   g452(.A(new_n618), .B(KEYINPUT105), .Z(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(new_n815), .ZN(new_n879));
  OR2_X1    g454(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n870), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n851), .B1(new_n865), .B2(new_n882), .ZN(new_n883));
  NAND4_X1  g458(.A1(new_n864), .A2(new_n880), .A3(KEYINPUT111), .A4(new_n881), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n865), .A2(new_n882), .ZN(new_n885));
  AND3_X1   g460(.A1(new_n883), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n850), .B1(new_n886), .B2(new_n605), .ZN(G295));
  OAI21_X1  g462(.A(new_n850), .B1(new_n886), .B2(new_n605), .ZN(G331));
  INV_X1    g463(.A(KEYINPUT44), .ZN(new_n889));
  XNOR2_X1  g464(.A(G168), .B(G171), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n815), .B(new_n890), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n891), .A2(new_n870), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n892), .B1(new_n877), .B2(new_n891), .ZN(new_n893));
  AOI21_X1  g468(.A(G37), .B1(new_n893), .B2(new_n863), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n870), .B(KEYINPUT41), .ZN(new_n895));
  AND2_X1   g470(.A1(new_n895), .A2(new_n891), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n896), .A2(new_n892), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n894), .B1(new_n863), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(KEYINPUT43), .ZN(new_n899));
  OR2_X1    g474(.A1(new_n893), .A2(new_n863), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT43), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n900), .A2(new_n901), .A3(new_n894), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n889), .B1(new_n899), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n898), .A2(new_n901), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n900), .A2(new_n894), .A3(KEYINPUT43), .ZN(new_n905));
  AOI21_X1  g480(.A(KEYINPUT44), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n903), .A2(new_n906), .ZN(G397));
  INV_X1    g482(.A(G1384), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n831), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT45), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(G40), .ZN(new_n912));
  NOR3_X1   g487(.A1(new_n464), .A2(new_n912), .A3(new_n476), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  XOR2_X1   g490(.A(new_n915), .B(KEYINPUT112), .Z(new_n916));
  INV_X1    g491(.A(G1996), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n755), .B(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(G2067), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n796), .B(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n698), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n922), .A2(new_n692), .A3(new_n693), .ZN(new_n923));
  OAI22_X1  g498(.A1(new_n921), .A2(new_n923), .B1(G2067), .B2(new_n796), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n916), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g500(.A1(G290), .A2(G1986), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n916), .A2(new_n926), .ZN(new_n927));
  XNOR2_X1  g502(.A(KEYINPUT127), .B(KEYINPUT48), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n921), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n694), .B(new_n922), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n916), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n929), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n927), .A2(new_n928), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n925), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n916), .A2(new_n917), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n937), .B(KEYINPUT46), .ZN(new_n938));
  INV_X1    g513(.A(new_n920), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n916), .B1(new_n755), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  XOR2_X1   g516(.A(KEYINPUT126), .B(KEYINPUT47), .Z(new_n942));
  OR2_X1    g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n941), .A2(new_n942), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n936), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT125), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT54), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n504), .A2(new_n828), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(new_n908), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT50), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(G1384), .B1(new_n499), .B2(new_n504), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(KEYINPUT50), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(G1961), .B1(new_n954), .B2(new_n913), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n913), .B1(new_n952), .B2(KEYINPUT45), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT113), .ZN(new_n958));
  NOR3_X1   g533(.A1(new_n829), .A2(new_n830), .A3(G1384), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n958), .B1(new_n959), .B2(KEYINPUT45), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n948), .A2(KEYINPUT103), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n495), .B1(new_n501), .B2(new_n503), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(new_n827), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n961), .A2(KEYINPUT45), .A3(new_n908), .A4(new_n963), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n964), .A2(KEYINPUT113), .ZN(new_n965));
  OAI211_X1 g540(.A(new_n443), .B(new_n957), .C1(new_n960), .C2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT53), .ZN(new_n967));
  AOI211_X1 g542(.A(G171), .B(new_n955), .C1(new_n966), .C2(new_n967), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n962), .A2(G1384), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n913), .B1(new_n969), .B2(KEYINPUT45), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(KEYINPUT116), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT117), .ZN(new_n972));
  INV_X1    g547(.A(new_n952), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n972), .B1(new_n973), .B2(new_n910), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT116), .ZN(new_n975));
  OAI211_X1 g550(.A(new_n975), .B(new_n913), .C1(new_n969), .C2(KEYINPUT45), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n952), .A2(KEYINPUT117), .A3(KEYINPUT45), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n971), .A2(new_n974), .A3(new_n976), .A4(new_n977), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n967), .A2(G2078), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  OR2_X1    g555(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n947), .B1(new_n968), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n966), .A2(new_n967), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT122), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n959), .A2(KEYINPUT45), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n984), .B1(new_n985), .B2(new_n914), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n911), .A2(KEYINPUT122), .A3(new_n913), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n964), .A2(KEYINPUT113), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n831), .A2(new_n958), .A3(KEYINPUT45), .A4(new_n908), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n980), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n986), .A2(new_n987), .A3(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT123), .ZN(new_n992));
  INV_X1    g567(.A(new_n955), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n983), .A2(new_n991), .A3(new_n992), .A4(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(G171), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n955), .B1(new_n966), .B2(new_n967), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n992), .B1(new_n996), .B2(new_n991), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n982), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n954), .A2(new_n774), .A3(new_n913), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n956), .B1(new_n988), .B2(new_n989), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n999), .B1(new_n1000), .B2(G1971), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(KEYINPUT114), .ZN(new_n1002));
  NAND2_X1  g577(.A1(G303), .A2(G8), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT115), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT55), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1003), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1006), .B1(new_n1005), .B2(new_n1003), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1004), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT114), .ZN(new_n1011));
  OAI211_X1 g586(.A(new_n1011), .B(new_n999), .C1(new_n1000), .C2(G1971), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1002), .A2(G8), .A3(new_n1010), .A4(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n957), .B1(new_n960), .B2(new_n965), .ZN(new_n1014));
  OR2_X1    g589(.A1(new_n952), .A2(KEYINPUT50), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n969), .A2(KEYINPUT50), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n914), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  AOI22_X1  g592(.A1(new_n1014), .A2(new_n713), .B1(new_n774), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(G8), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1009), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(G305), .A2(G1981), .ZN(new_n1021));
  OR3_X1    g596(.A1(new_n581), .A2(new_n583), .A3(G1981), .ZN(new_n1022));
  AND2_X1   g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  OR2_X1    g598(.A1(new_n1023), .A2(KEYINPUT49), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n914), .A2(new_n949), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1025), .A2(new_n1019), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1023), .A2(KEYINPUT49), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1024), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(G1976), .ZN(new_n1029));
  AOI21_X1  g604(.A(KEYINPUT52), .B1(G288), .B2(new_n1029), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n1026), .B(new_n1030), .C1(new_n1029), .C2(G288), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1026), .ZN(new_n1032));
  NOR2_X1   g607(.A1(G288), .A2(new_n1029), .ZN(new_n1033));
  OAI21_X1  g608(.A(KEYINPUT52), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  AND3_X1   g609(.A1(new_n1028), .A2(new_n1031), .A3(new_n1034), .ZN(new_n1035));
  AND3_X1   g610(.A1(new_n1013), .A2(new_n1020), .A3(new_n1035), .ZN(new_n1036));
  AND3_X1   g611(.A1(new_n996), .A2(G301), .A3(new_n991), .ZN(new_n1037));
  AOI21_X1  g612(.A(G301), .B1(new_n996), .B2(new_n981), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n947), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  AOI211_X1 g614(.A(G2084), .B(new_n914), .C1(new_n951), .C2(new_n953), .ZN(new_n1040));
  INV_X1    g615(.A(G1966), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1040), .B1(new_n978), .B2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(KEYINPUT51), .B1(new_n1042), .B2(G168), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1019), .B1(new_n1042), .B2(G168), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  AOI211_X1 g620(.A(G286), .B(new_n1040), .C1(new_n978), .C2(new_n1041), .ZN(new_n1046));
  OAI21_X1  g621(.A(KEYINPUT51), .B1(new_n1046), .B2(new_n1019), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n998), .A2(new_n1036), .A3(new_n1039), .A4(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(KEYINPUT124), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n983), .A2(new_n981), .A3(new_n993), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(G171), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n996), .A2(G301), .A3(new_n991), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  AOI22_X1  g629(.A1(new_n1054), .A2(new_n947), .B1(new_n1047), .B2(new_n1045), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT124), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1055), .A2(new_n1056), .A3(new_n1036), .A4(new_n998), .ZN(new_n1057));
  XNOR2_X1  g632(.A(KEYINPUT56), .B(G2072), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1000), .A2(new_n1058), .ZN(new_n1059));
  OR2_X1    g634(.A1(new_n1017), .A2(G1956), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT119), .ZN(new_n1062));
  XNOR2_X1  g637(.A(new_n1061), .B(new_n1062), .ZN(new_n1063));
  XOR2_X1   g638(.A(G299), .B(KEYINPUT57), .Z(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1064), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n954), .A2(new_n913), .ZN(new_n1067));
  AOI22_X1  g642(.A1(new_n1067), .A2(new_n780), .B1(new_n919), .B2(new_n1025), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1068), .A2(new_n603), .ZN(new_n1069));
  AOI22_X1  g644(.A1(new_n1063), .A2(new_n1065), .B1(new_n1066), .B2(new_n1069), .ZN(new_n1070));
  XNOR2_X1  g645(.A(KEYINPUT58), .B(G1341), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1025), .A2(new_n1071), .ZN(new_n1072));
  XNOR2_X1  g647(.A(KEYINPUT120), .B(G1996), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1072), .B1(new_n1000), .B2(new_n1073), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1074), .A2(new_n546), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT59), .ZN(new_n1076));
  XNOR2_X1  g651(.A(new_n1075), .B(new_n1076), .ZN(new_n1077));
  XOR2_X1   g652(.A(KEYINPUT121), .B(KEYINPUT61), .Z(new_n1078));
  INV_X1    g653(.A(new_n1066), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1064), .B1(new_n1060), .B2(new_n1059), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1078), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  XNOR2_X1  g656(.A(new_n1068), .B(new_n603), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n603), .A2(KEYINPUT60), .ZN(new_n1083));
  AOI22_X1  g658(.A1(new_n1082), .A2(KEYINPUT60), .B1(new_n1068), .B2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1077), .A2(new_n1081), .A3(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1066), .A2(KEYINPUT61), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1086), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1070), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1050), .A2(new_n1057), .A3(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1048), .A2(KEYINPUT62), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT62), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1045), .A2(new_n1047), .A3(new_n1091), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1090), .A2(new_n1036), .A3(new_n1038), .A4(new_n1092), .ZN(new_n1093));
  NOR3_X1   g668(.A1(new_n1042), .A2(new_n1019), .A3(G286), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1013), .A2(new_n1020), .A3(new_n1035), .A4(new_n1094), .ZN(new_n1095));
  XNOR2_X1  g670(.A(KEYINPUT118), .B(KEYINPUT63), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1002), .A2(G8), .A3(new_n1012), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(new_n1009), .ZN(new_n1099));
  AND2_X1   g674(.A1(new_n1094), .A2(KEYINPUT63), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1099), .A2(new_n1100), .A3(new_n1013), .A4(new_n1035), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1097), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(G288), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1028), .A2(new_n1029), .A3(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1032), .B1(new_n1104), .B2(new_n1022), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1013), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1105), .B1(new_n1106), .B2(new_n1035), .ZN(new_n1107));
  AND3_X1   g682(.A1(new_n1093), .A2(new_n1102), .A3(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1089), .A2(new_n1108), .ZN(new_n1109));
  AND2_X1   g684(.A1(G290), .A2(G1986), .ZN(new_n1110));
  OR3_X1    g685(.A1(new_n932), .A2(new_n926), .A3(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n916), .A2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n946), .B1(new_n1109), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1112), .ZN(new_n1114));
  AOI211_X1 g689(.A(KEYINPUT125), .B(new_n1114), .C1(new_n1089), .C2(new_n1108), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n945), .B1(new_n1113), .B2(new_n1115), .ZN(G329));
  assign    G231 = 1'b0;
  NAND4_X1  g691(.A1(new_n687), .A2(G319), .A3(new_n652), .A4(new_n668), .ZN(new_n1118));
  AOI21_X1  g692(.A(new_n1118), .B1(new_n846), .B2(new_n847), .ZN(new_n1119));
  NAND3_X1  g693(.A1(new_n1119), .A2(new_n904), .A3(new_n905), .ZN(G225));
  INV_X1    g694(.A(G225), .ZN(G308));
endmodule


