//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 1 0 0 1 0 0 0 0 1 1 1 1 1 0 1 0 0 1 0 1 1 0 1 1 1 0 0 1 1 1 1 0 0 1 1 1 1 1 0 1 1 0 1 1 0 1 0 1 1 1 0 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n630, new_n631,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n807,
    new_n808, new_n809, new_n810, new_n812, new_n813, new_n814, new_n815,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n860,
    new_n861, new_n863, new_n864, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n874, new_n875, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n913, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925;
  XNOR2_X1  g000(.A(G197gat), .B(G204gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT70), .ZN(new_n203));
  XNOR2_X1  g002(.A(G211gat), .B(G218gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT22), .ZN(new_n205));
  AOI22_X1  g004(.A1(new_n205), .A2(KEYINPUT71), .B1(G211gat), .B2(G218gat), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n206), .B1(KEYINPUT71), .B2(new_n205), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n203), .A2(new_n204), .A3(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  AOI21_X1  g008(.A(new_n204), .B1(new_n203), .B2(new_n207), .ZN(new_n210));
  OR2_X1    g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT29), .ZN(new_n212));
  XNOR2_X1  g011(.A(G155gat), .B(G162gat), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G141gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(G148gat), .ZN(new_n216));
  INV_X1    g015(.A(G148gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(G141gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(KEYINPUT75), .ZN(new_n220));
  INV_X1    g019(.A(G155gat), .ZN(new_n221));
  INV_X1    g020(.A(G162gat), .ZN(new_n222));
  OAI21_X1  g021(.A(KEYINPUT2), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n220), .A2(new_n223), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n219), .A2(KEYINPUT75), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n214), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  OR2_X1    g025(.A1(new_n213), .A2(KEYINPUT77), .ZN(new_n227));
  OR3_X1    g026(.A1(new_n215), .A2(KEYINPUT76), .A3(G148gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n218), .A2(KEYINPUT76), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n228), .A2(new_n229), .A3(new_n216), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n213), .A2(KEYINPUT77), .ZN(new_n231));
  NAND4_X1  g030(.A1(new_n227), .A2(new_n230), .A3(new_n223), .A4(new_n231), .ZN(new_n232));
  AND2_X1   g031(.A1(new_n226), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT3), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n211), .B1(new_n212), .B2(new_n235), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n212), .B1(new_n209), .B2(new_n210), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n233), .B1(new_n237), .B2(new_n234), .ZN(new_n238));
  OAI21_X1  g037(.A(KEYINPUT81), .B1(new_n236), .B2(new_n238), .ZN(new_n239));
  XOR2_X1   g038(.A(KEYINPUT79), .B(KEYINPUT31), .Z(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n240), .ZN(new_n242));
  OAI211_X1 g041(.A(KEYINPUT81), .B(new_n242), .C1(new_n236), .C2(new_n238), .ZN(new_n243));
  XOR2_X1   g042(.A(G78gat), .B(G106gat), .Z(new_n244));
  XNOR2_X1  g043(.A(new_n244), .B(KEYINPUT80), .ZN(new_n245));
  INV_X1    g044(.A(G50gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n245), .B(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(G228gat), .A2(G233gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n248), .B(G22gat), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n247), .B(new_n249), .ZN(new_n250));
  AND3_X1   g049(.A1(new_n241), .A2(new_n243), .A3(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n250), .B1(new_n241), .B2(new_n243), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NOR2_X1   g052(.A1(G169gat), .A2(G176gat), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(KEYINPUT23), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT23), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n256), .B1(G169gat), .B2(G176gat), .ZN(new_n257));
  INV_X1    g056(.A(G169gat), .ZN(new_n258));
  INV_X1    g057(.A(G176gat), .ZN(new_n259));
  OAI211_X1 g058(.A(new_n255), .B(new_n257), .C1(new_n258), .C2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT25), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(G183gat), .A2(G190gat), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n264), .B1(KEYINPUT64), .B2(KEYINPUT24), .ZN(new_n265));
  AND2_X1   g064(.A1(KEYINPUT64), .A2(KEYINPUT24), .ZN(new_n266));
  OAI221_X1 g065(.A(new_n263), .B1(G183gat), .B2(G190gat), .C1(new_n265), .C2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n262), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT65), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n262), .A2(KEYINPUT65), .A3(new_n267), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n263), .B1(G183gat), .B2(G190gat), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT24), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n272), .B1(new_n273), .B2(new_n264), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n261), .B1(new_n274), .B2(new_n260), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n270), .A2(new_n271), .A3(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(KEYINPUT27), .B(G183gat), .ZN(new_n277));
  INV_X1    g076(.A(G190gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT28), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(KEYINPUT66), .ZN(new_n281));
  OR2_X1    g080(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  OR2_X1    g081(.A1(new_n280), .A2(KEYINPUT66), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n279), .A2(new_n281), .A3(new_n283), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n254), .A2(KEYINPUT26), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n285), .B1(new_n258), .B2(new_n259), .ZN(new_n286));
  AOI22_X1  g085(.A1(new_n254), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n282), .A2(new_n284), .A3(new_n286), .A4(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n276), .A2(new_n288), .ZN(new_n289));
  XOR2_X1   g088(.A(G113gat), .B(G120gat), .Z(new_n290));
  INV_X1    g089(.A(KEYINPUT1), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(G127gat), .B(G134gat), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n292), .B(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n294), .B(KEYINPUT67), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n289), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(G227gat), .ZN(new_n297));
  INV_X1    g096(.A(G233gat), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  OR2_X1    g098(.A1(new_n294), .A2(KEYINPUT67), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n294), .A2(KEYINPUT67), .ZN(new_n301));
  NAND4_X1  g100(.A1(new_n300), .A2(new_n276), .A3(new_n301), .A4(new_n288), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n296), .A2(new_n299), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT32), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT33), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  XOR2_X1   g105(.A(G15gat), .B(G43gat), .Z(new_n307));
  XNOR2_X1  g106(.A(G71gat), .B(G99gat), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n307), .B(new_n308), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n304), .A2(new_n306), .A3(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n309), .ZN(new_n311));
  OAI211_X1 g110(.A(new_n303), .B(KEYINPUT32), .C1(new_n305), .C2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n296), .A2(new_n302), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  OAI21_X1  g114(.A(KEYINPUT34), .B1(new_n315), .B2(new_n299), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT34), .ZN(new_n317));
  OAI211_X1 g116(.A(new_n314), .B(new_n317), .C1(new_n297), .C2(new_n298), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  AND2_X1   g118(.A1(new_n313), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT69), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n321), .B1(new_n313), .B2(new_n319), .ZN(new_n322));
  INV_X1    g121(.A(new_n319), .ZN(new_n323));
  NAND4_X1  g122(.A1(new_n323), .A2(KEYINPUT69), .A3(new_n310), .A4(new_n312), .ZN(new_n324));
  AOI211_X1 g123(.A(new_n253), .B(new_n320), .C1(new_n322), .C2(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n295), .A2(KEYINPUT4), .A3(new_n233), .ZN(new_n326));
  NAND2_X1  g125(.A1(G225gat), .A2(G233gat), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n226), .A2(new_n232), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n294), .B1(new_n329), .B2(KEYINPUT3), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n328), .B1(new_n235), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n233), .A2(new_n294), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT4), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n326), .A2(new_n331), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(KEYINPUT78), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT78), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n326), .A2(new_n331), .A3(new_n337), .A4(new_n334), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n329), .B(new_n294), .ZN(new_n340));
  OAI21_X1  g139(.A(KEYINPUT5), .B1(new_n340), .B2(new_n327), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  XNOR2_X1  g142(.A(G1gat), .B(G29gat), .ZN(new_n344));
  XNOR2_X1  g143(.A(new_n344), .B(KEYINPUT0), .ZN(new_n345));
  XNOR2_X1  g144(.A(G57gat), .B(G85gat), .ZN(new_n346));
  XOR2_X1   g145(.A(new_n345), .B(new_n346), .Z(new_n347));
  NOR2_X1   g146(.A1(new_n332), .A2(new_n333), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n295), .A2(new_n233), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n348), .B1(new_n349), .B2(new_n333), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT5), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n350), .A2(new_n351), .A3(new_n331), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n343), .A2(new_n347), .A3(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n347), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n341), .B1(new_n336), .B2(new_n338), .ZN(new_n355));
  INV_X1    g154(.A(new_n352), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n354), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT6), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n353), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT82), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n357), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(KEYINPUT6), .ZN(new_n363));
  NAND4_X1  g162(.A1(new_n353), .A2(new_n357), .A3(KEYINPUT82), .A4(new_n358), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n361), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT35), .ZN(new_n366));
  INV_X1    g165(.A(G226gat), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n367), .A2(new_n298), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(new_n212), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n289), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n276), .A2(new_n288), .A3(new_n369), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n211), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n371), .A2(new_n211), .A3(new_n372), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT72), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n375), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  OR2_X1    g177(.A1(new_n376), .A2(new_n377), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  XOR2_X1   g179(.A(G8gat), .B(G36gat), .Z(new_n381));
  XNOR2_X1  g180(.A(new_n381), .B(KEYINPUT73), .ZN(new_n382));
  XNOR2_X1  g181(.A(G64gat), .B(G92gat), .ZN(new_n383));
  XOR2_X1   g182(.A(new_n382), .B(new_n383), .Z(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(KEYINPUT30), .B1(new_n380), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n380), .A2(new_n385), .ZN(new_n387));
  XOR2_X1   g186(.A(new_n384), .B(KEYINPUT74), .Z(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n387), .B1(new_n380), .B2(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n386), .B1(new_n390), .B2(KEYINPUT30), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n325), .A2(new_n365), .A3(new_n366), .A4(new_n391), .ZN(new_n392));
  AND3_X1   g191(.A1(new_n316), .A2(KEYINPUT68), .A3(new_n318), .ZN(new_n393));
  AOI21_X1  g192(.A(KEYINPUT68), .B1(new_n316), .B2(new_n318), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AOI22_X1  g194(.A1(new_n322), .A2(new_n324), .B1(new_n395), .B2(new_n313), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n363), .A2(new_n359), .ZN(new_n397));
  INV_X1    g196(.A(new_n253), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n396), .A2(new_n397), .A3(new_n391), .A4(new_n398), .ZN(new_n399));
  AOI22_X1  g198(.A1(new_n392), .A2(KEYINPUT83), .B1(KEYINPUT35), .B2(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n320), .B1(new_n324), .B2(new_n322), .ZN(new_n401));
  AND3_X1   g200(.A1(new_n391), .A2(new_n401), .A3(new_n398), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT83), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n402), .A2(new_n403), .A3(new_n366), .A4(new_n365), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT38), .ZN(new_n405));
  AND2_X1   g204(.A1(new_n375), .A2(new_n376), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT37), .ZN(new_n407));
  OAI211_X1 g206(.A(new_n405), .B(new_n388), .C1(new_n406), .C2(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(KEYINPUT37), .B1(new_n378), .B2(new_n379), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n387), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n384), .B1(new_n380), .B2(new_n407), .ZN(new_n411));
  OR2_X1    g210(.A1(new_n411), .A2(new_n409), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n410), .B1(new_n412), .B2(KEYINPUT38), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n413), .A2(new_n363), .A3(new_n361), .A4(new_n364), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n235), .A2(new_n330), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n350), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(new_n328), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT39), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n418), .B1(new_n340), .B2(new_n327), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n420), .B(new_n347), .C1(KEYINPUT39), .C2(new_n417), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT40), .ZN(new_n422));
  AND2_X1   g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n421), .A2(new_n422), .ZN(new_n424));
  NOR3_X1   g223(.A1(new_n423), .A2(new_n424), .A3(new_n362), .ZN(new_n425));
  INV_X1    g224(.A(new_n391), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n414), .A2(new_n427), .A3(new_n398), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n398), .B1(new_n397), .B2(new_n391), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT36), .ZN(new_n430));
  AND2_X1   g229(.A1(new_n401), .A2(new_n430), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n396), .A2(new_n430), .ZN(new_n432));
  NOR3_X1   g231(.A1(new_n429), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  AOI22_X1  g232(.A1(new_n400), .A2(new_n404), .B1(new_n428), .B2(new_n433), .ZN(new_n434));
  OR3_X1    g233(.A1(KEYINPUT84), .A2(G29gat), .A3(G36gat), .ZN(new_n435));
  OAI21_X1  g234(.A(KEYINPUT84), .B1(G29gat), .B2(G36gat), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n435), .A2(KEYINPUT14), .A3(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(G29gat), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(KEYINPUT85), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT85), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(G29gat), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(G36gat), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n246), .A2(G43gat), .ZN(new_n444));
  INV_X1    g243(.A(G43gat), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(G50gat), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT15), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  OR2_X1    g248(.A1(new_n436), .A2(KEYINPUT14), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n437), .A2(new_n443), .A3(new_n449), .A4(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n444), .A2(new_n446), .A3(KEYINPUT15), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  AOI22_X1  g253(.A1(new_n448), .A2(new_n447), .B1(new_n442), .B2(G36gat), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n455), .A2(new_n452), .A3(new_n437), .A4(new_n450), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n454), .A2(new_n456), .A3(KEYINPUT17), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT86), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n454), .A2(new_n456), .A3(KEYINPUT86), .A4(KEYINPUT17), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  XNOR2_X1  g260(.A(G15gat), .B(G22gat), .ZN(new_n462));
  INV_X1    g261(.A(G1gat), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(KEYINPUT16), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n465), .B1(G1gat), .B2(new_n462), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n466), .B(G8gat), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT17), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n454), .A2(new_n456), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n461), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(G229gat), .A2(G233gat), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n467), .A2(new_n469), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n471), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT18), .ZN(new_n475));
  XNOR2_X1  g274(.A(new_n467), .B(new_n469), .ZN(new_n476));
  XOR2_X1   g275(.A(new_n472), .B(KEYINPUT13), .Z(new_n477));
  AOI22_X1  g276(.A1(new_n474), .A2(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n473), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n479), .B1(new_n461), .B2(new_n470), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n480), .A2(KEYINPUT18), .A3(new_n472), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  XNOR2_X1  g281(.A(G113gat), .B(G141gat), .ZN(new_n483));
  XNOR2_X1  g282(.A(new_n483), .B(G197gat), .ZN(new_n484));
  XOR2_X1   g283(.A(KEYINPUT11), .B(G169gat), .Z(new_n485));
  XNOR2_X1  g284(.A(new_n484), .B(new_n485), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n486), .B(KEYINPUT12), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n474), .A2(new_n475), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT87), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n482), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(KEYINPUT87), .B1(new_n474), .B2(new_n475), .ZN(new_n492));
  OAI211_X1 g291(.A(new_n478), .B(new_n481), .C1(new_n492), .C2(new_n487), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT88), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n491), .A2(KEYINPUT88), .A3(new_n493), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n434), .A2(new_n499), .ZN(new_n500));
  XOR2_X1   g299(.A(G99gat), .B(G106gat), .Z(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(KEYINPUT93), .A2(G85gat), .A3(G92gat), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT7), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g304(.A1(KEYINPUT93), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n506));
  AND2_X1   g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(G99gat), .A2(G106gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(KEYINPUT8), .ZN(new_n509));
  OR2_X1    g308(.A1(KEYINPUT94), .A2(G85gat), .ZN(new_n510));
  INV_X1    g309(.A(G92gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(KEYINPUT94), .A2(G85gat), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n502), .A2(new_n507), .A3(new_n509), .A4(new_n513), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n513), .A2(new_n509), .A3(new_n505), .A4(new_n506), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(new_n501), .ZN(new_n516));
  AND2_X1   g315(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n517), .B1(new_n469), .B2(new_n468), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n461), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(G232gat), .A2(G233gat), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  AOI22_X1  g320(.A1(new_n469), .A2(new_n517), .B1(KEYINPUT41), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(G190gat), .B(G218gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n524), .B(KEYINPUT95), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n523), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n519), .A2(new_n525), .A3(new_n522), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n521), .A2(KEYINPUT41), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n529), .B(KEYINPUT91), .ZN(new_n530));
  XOR2_X1   g329(.A(G134gat), .B(G162gat), .Z(new_n531));
  XNOR2_X1  g330(.A(new_n530), .B(new_n531), .ZN(new_n532));
  AND3_X1   g331(.A1(new_n527), .A2(new_n528), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n528), .A2(KEYINPUT96), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT96), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n519), .A2(new_n535), .A3(new_n525), .A4(new_n522), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n534), .A2(new_n536), .A3(new_n527), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n532), .B(KEYINPUT92), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n533), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  AND2_X1   g340(.A1(G71gat), .A2(G78gat), .ZN(new_n542));
  NOR2_X1   g341(.A1(G71gat), .A2(G78gat), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(G57gat), .B(G64gat), .ZN(new_n545));
  AOI21_X1  g344(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(G57gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(G64gat), .ZN(new_n549));
  INV_X1    g348(.A(G64gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(G57gat), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(G71gat), .B(G78gat), .ZN(new_n553));
  INV_X1    g352(.A(new_n546), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  AND3_X1   g354(.A1(new_n547), .A2(new_n555), .A3(KEYINPUT97), .ZN(new_n556));
  AOI21_X1  g355(.A(KEYINPUT97), .B1(new_n547), .B2(new_n555), .ZN(new_n557));
  OAI211_X1 g356(.A(new_n514), .B(new_n516), .C1(new_n556), .C2(new_n557), .ZN(new_n558));
  AND2_X1   g357(.A1(new_n515), .A2(new_n501), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n515), .A2(new_n501), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT97), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n547), .A2(new_n555), .ZN(new_n562));
  OAI22_X1  g361(.A1(new_n559), .A2(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT10), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n558), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT98), .ZN(new_n566));
  AND3_X1   g365(.A1(new_n547), .A2(new_n555), .A3(KEYINPUT90), .ZN(new_n567));
  AOI21_X1  g366(.A(KEYINPUT90), .B1(new_n547), .B2(new_n555), .ZN(new_n568));
  OAI21_X1  g367(.A(KEYINPUT10), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n514), .A2(new_n516), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n566), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT90), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n562), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n547), .A2(new_n555), .A3(KEYINPUT90), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n575), .A2(new_n517), .A3(KEYINPUT98), .A4(KEYINPUT10), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n565), .A2(new_n571), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(G230gat), .A2(G233gat), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(G120gat), .B(G148gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(G176gat), .B(G204gat), .ZN(new_n581));
  XOR2_X1   g380(.A(new_n580), .B(new_n581), .Z(new_n582));
  NAND2_X1  g381(.A1(new_n558), .A2(new_n563), .ZN(new_n583));
  INV_X1    g382(.A(new_n578), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n579), .A2(new_n582), .A3(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT99), .ZN(new_n587));
  AND3_X1   g386(.A1(new_n577), .A2(new_n587), .A3(new_n578), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n587), .B1(new_n577), .B2(new_n578), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n585), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT100), .ZN(new_n591));
  INV_X1    g390(.A(new_n582), .ZN(new_n592));
  AND3_X1   g391(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n591), .B1(new_n590), .B2(new_n592), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n586), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n467), .B1(KEYINPUT21), .B2(new_n575), .ZN(new_n596));
  AOI21_X1  g395(.A(KEYINPUT21), .B1(new_n547), .B2(new_n555), .ZN(new_n597));
  XOR2_X1   g396(.A(G127gat), .B(G155gat), .Z(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n596), .B(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(G231gat), .A2(G233gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(KEYINPUT89), .ZN(new_n602));
  XOR2_X1   g401(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(G183gat), .B(G211gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n600), .B(new_n606), .ZN(new_n607));
  NOR3_X1   g406(.A1(new_n541), .A2(new_n595), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n500), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n609), .A2(new_n397), .ZN(new_n610));
  XNOR2_X1  g409(.A(KEYINPUT101), .B(G1gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(G1324gat));
  INV_X1    g411(.A(new_n609), .ZN(new_n613));
  XOR2_X1   g412(.A(KEYINPUT16), .B(G8gat), .Z(new_n614));
  NAND4_X1  g413(.A1(new_n613), .A2(KEYINPUT42), .A3(new_n426), .A4(new_n614), .ZN(new_n615));
  OR3_X1    g414(.A1(new_n609), .A2(KEYINPUT102), .A3(new_n391), .ZN(new_n616));
  OAI21_X1  g415(.A(KEYINPUT102), .B1(new_n609), .B2(new_n391), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n616), .A2(G8gat), .A3(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n614), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n619), .B1(new_n616), .B2(new_n617), .ZN(new_n620));
  OAI211_X1 g419(.A(new_n615), .B(new_n618), .C1(new_n620), .C2(KEYINPUT42), .ZN(G1325gat));
  NOR2_X1   g420(.A1(new_n431), .A2(new_n432), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  AND3_X1   g422(.A1(new_n613), .A2(G15gat), .A3(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(G15gat), .B1(new_n613), .B2(new_n401), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT103), .ZN(new_n626));
  OR2_X1    g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n625), .A2(new_n626), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n624), .B1(new_n627), .B2(new_n628), .ZN(G1326gat));
  NOR2_X1   g428(.A1(new_n609), .A2(new_n398), .ZN(new_n630));
  XOR2_X1   g429(.A(KEYINPUT43), .B(G22gat), .Z(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(G1327gat));
  NAND2_X1  g431(.A1(new_n392), .A2(KEYINPUT83), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n399), .A2(KEYINPUT35), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n633), .A2(new_n404), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n433), .A2(new_n428), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n607), .ZN(new_n638));
  NOR3_X1   g437(.A1(new_n595), .A2(new_n638), .A3(new_n540), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n637), .A2(new_n498), .A3(new_n639), .ZN(new_n640));
  NOR3_X1   g439(.A1(new_n640), .A2(new_n397), .A3(new_n442), .ZN(new_n641));
  XOR2_X1   g440(.A(new_n641), .B(KEYINPUT45), .Z(new_n642));
  INV_X1    g441(.A(KEYINPUT44), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n643), .B1(new_n434), .B2(new_n540), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n637), .A2(KEYINPUT44), .A3(new_n541), .ZN(new_n645));
  AND2_X1   g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n494), .ZN(new_n647));
  NOR3_X1   g446(.A1(new_n647), .A2(new_n595), .A3(new_n638), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n442), .B1(new_n649), .B2(new_n397), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n642), .A2(new_n650), .ZN(G1328gat));
  OAI21_X1  g450(.A(G36gat), .B1(new_n649), .B2(new_n391), .ZN(new_n652));
  OR2_X1    g451(.A1(new_n391), .A2(G36gat), .ZN(new_n653));
  OAI22_X1  g452(.A1(new_n640), .A2(new_n653), .B1(KEYINPUT104), .B2(KEYINPUT46), .ZN(new_n654));
  NAND2_X1  g453(.A1(KEYINPUT104), .A2(KEYINPUT46), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  OR2_X1    g455(.A1(new_n654), .A2(new_n655), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n652), .A2(new_n656), .A3(new_n657), .ZN(G1329gat));
  INV_X1    g457(.A(new_n401), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n445), .B1(new_n640), .B2(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n622), .A2(new_n445), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n660), .B1(new_n649), .B2(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g463(.A1(new_n644), .A2(new_n645), .A3(new_n253), .A4(new_n648), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n665), .A2(G50gat), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT105), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n500), .A2(new_n667), .A3(new_n639), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n640), .A2(KEYINPUT105), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n253), .A2(new_n246), .ZN(new_n670));
  XOR2_X1   g469(.A(new_n670), .B(KEYINPUT106), .Z(new_n671));
  NAND3_X1  g470(.A1(new_n668), .A2(new_n669), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n666), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT107), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n666), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n673), .A2(new_n675), .A3(KEYINPUT48), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT48), .ZN(new_n677));
  OAI211_X1 g476(.A(new_n666), .B(new_n672), .C1(new_n674), .C2(new_n677), .ZN(new_n678));
  AND2_X1   g477(.A1(new_n676), .A2(new_n678), .ZN(G1331gat));
  INV_X1    g478(.A(new_n595), .ZN(new_n680));
  NOR4_X1   g479(.A1(new_n680), .A2(new_n541), .A3(new_n494), .A4(new_n607), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n637), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n682), .A2(new_n397), .ZN(new_n683));
  XNOR2_X1  g482(.A(KEYINPUT108), .B(G57gat), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n683), .B(new_n684), .ZN(G1332gat));
  INV_X1    g484(.A(new_n682), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n391), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(KEYINPUT109), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT110), .ZN(new_n690));
  OR2_X1    g489(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n690), .B(new_n691), .ZN(G1333gat));
  NOR3_X1   g491(.A1(new_n682), .A2(G71gat), .A3(new_n659), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n686), .A2(new_n623), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n693), .B1(G71gat), .B2(new_n694), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g495(.A1(new_n682), .A2(new_n398), .ZN(new_n697));
  XNOR2_X1  g496(.A(KEYINPUT111), .B(G78gat), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n697), .B(new_n698), .ZN(G1335gat));
  NAND2_X1  g498(.A1(new_n510), .A2(new_n512), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n397), .A2(new_n700), .A3(new_n680), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT51), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n637), .A2(new_n541), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n494), .A2(new_n638), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n702), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n706), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n703), .A2(new_n702), .A3(new_n705), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n707), .A2(new_n708), .A3(KEYINPUT112), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT112), .ZN(new_n710));
  INV_X1    g509(.A(new_n708), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n710), .B1(new_n711), .B2(new_n706), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n701), .B1(new_n709), .B2(new_n712), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n705), .A2(new_n680), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n646), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n700), .B1(new_n715), .B2(new_n397), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n713), .A2(new_n716), .ZN(G1336gat));
  NOR2_X1   g516(.A1(new_n391), .A2(G92gat), .ZN(new_n718));
  OAI211_X1 g517(.A(new_n595), .B(new_n718), .C1(new_n707), .C2(new_n708), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n644), .A2(new_n645), .A3(new_n426), .A4(new_n714), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(G92gat), .ZN(new_n721));
  XNOR2_X1  g520(.A(KEYINPUT113), .B(KEYINPUT52), .ZN(new_n722));
  AND3_X1   g521(.A1(new_n719), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n722), .B1(new_n719), .B2(new_n721), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n723), .A2(new_n724), .ZN(G1337gat));
  XOR2_X1   g524(.A(KEYINPUT114), .B(G99gat), .Z(new_n726));
  NOR3_X1   g525(.A1(new_n659), .A2(new_n680), .A3(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n727), .B1(new_n709), .B2(new_n712), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n726), .B1(new_n715), .B2(new_n622), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(G1338gat));
  NOR2_X1   g529(.A1(new_n398), .A2(G106gat), .ZN(new_n731));
  OAI211_X1 g530(.A(new_n595), .B(new_n731), .C1(new_n707), .C2(new_n708), .ZN(new_n732));
  NAND4_X1  g531(.A1(new_n644), .A2(new_n645), .A3(new_n253), .A4(new_n714), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(G106gat), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(KEYINPUT53), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT53), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n732), .A2(new_n737), .A3(new_n734), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n736), .A2(new_n738), .ZN(G1339gat));
  NOR2_X1   g538(.A1(new_n647), .A2(G113gat), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n579), .A2(KEYINPUT99), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT54), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n577), .A2(new_n587), .A3(new_n578), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n741), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT115), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n565), .A2(new_n571), .A3(new_n576), .A4(new_n584), .ZN(new_n746));
  AND4_X1   g545(.A1(new_n745), .A2(new_n579), .A3(KEYINPUT54), .A4(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n742), .B1(new_n577), .B2(new_n578), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n745), .B1(new_n748), .B2(new_n746), .ZN(new_n749));
  OAI211_X1 g548(.A(new_n592), .B(new_n744), .C1(new_n747), .C2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT55), .ZN(new_n751));
  OAI21_X1  g550(.A(KEYINPUT116), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(new_n586), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n753), .B1(new_n750), .B2(new_n751), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n588), .A2(new_n589), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n582), .B1(new_n755), .B2(new_n742), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n748), .A2(new_n746), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(KEYINPUT115), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n748), .A2(new_n745), .A3(new_n746), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT116), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n756), .A2(new_n760), .A3(new_n761), .A4(KEYINPUT55), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n752), .A2(new_n754), .A3(new_n494), .A4(new_n762), .ZN(new_n763));
  OAI22_X1  g562(.A1(new_n480), .A2(new_n472), .B1(new_n476), .B2(new_n477), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(new_n486), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n478), .A2(new_n487), .A3(new_n481), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n595), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n541), .B1(new_n763), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n766), .A2(new_n765), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n540), .A2(new_n769), .ZN(new_n770));
  AND4_X1   g569(.A1(new_n762), .A2(new_n770), .A3(new_n752), .A4(new_n754), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n607), .B1(new_n768), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n608), .A2(new_n647), .ZN(new_n773));
  AND3_X1   g572(.A1(new_n772), .A2(KEYINPUT117), .A3(new_n773), .ZN(new_n774));
  AOI21_X1  g573(.A(KEYINPUT117), .B1(new_n772), .B2(new_n773), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(new_n397), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n396), .A2(new_n398), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n778), .A2(new_n426), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n776), .A2(new_n777), .A3(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n781), .A2(KEYINPUT118), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT118), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n780), .A2(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n740), .B1(new_n782), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n772), .A2(new_n773), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT117), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n772), .A2(KEYINPUT117), .A3(new_n773), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n790), .A2(new_n397), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(new_n402), .ZN(new_n792));
  OAI21_X1  g591(.A(G113gat), .B1(new_n792), .B2(new_n499), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n785), .A2(new_n793), .ZN(G1340gat));
  NOR2_X1   g593(.A1(new_n680), .A2(G120gat), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n795), .B1(new_n782), .B2(new_n784), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n791), .A2(new_n402), .A3(new_n595), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT119), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n797), .A2(new_n798), .A3(G120gat), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n798), .B1(new_n797), .B2(G120gat), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n796), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT120), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  OAI211_X1 g603(.A(new_n796), .B(KEYINPUT120), .C1(new_n800), .C2(new_n801), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(G1341gat));
  NAND4_X1  g605(.A1(new_n791), .A2(G127gat), .A3(new_n402), .A4(new_n638), .ZN(new_n807));
  AND2_X1   g606(.A1(new_n807), .A2(KEYINPUT121), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n807), .A2(KEYINPUT121), .ZN(new_n809));
  AOI21_X1  g608(.A(G127gat), .B1(new_n781), .B2(new_n638), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n808), .A2(new_n809), .A3(new_n810), .ZN(G1342gat));
  INV_X1    g610(.A(G134gat), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n781), .A2(new_n812), .A3(new_n541), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n791), .A2(new_n402), .A3(new_n541), .ZN(new_n814));
  AOI22_X1  g613(.A1(new_n813), .A2(KEYINPUT56), .B1(new_n814), .B2(G134gat), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n815), .B1(KEYINPUT56), .B2(new_n813), .ZN(G1343gat));
  INV_X1    g615(.A(KEYINPUT58), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n623), .A2(new_n398), .A3(new_n426), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n776), .A2(new_n777), .A3(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n820), .A2(new_n215), .A3(new_n498), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT57), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n398), .A2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n752), .A2(new_n754), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n498), .A2(new_n825), .A3(new_n762), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n541), .B1(new_n826), .B2(new_n767), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n607), .B1(new_n827), .B2(new_n771), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n824), .B1(new_n828), .B2(new_n773), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n788), .A2(new_n253), .A3(new_n789), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n829), .B1(new_n830), .B2(new_n822), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n622), .A2(new_n777), .A3(new_n391), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n831), .A2(new_n499), .A3(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(G141gat), .B1(new_n833), .B2(KEYINPUT123), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n831), .A2(new_n832), .ZN(new_n835));
  AND3_X1   g634(.A1(new_n835), .A2(KEYINPUT123), .A3(new_n498), .ZN(new_n836));
  OAI211_X1 g635(.A(new_n817), .B(new_n821), .C1(new_n834), .C2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(new_n829), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n774), .A2(new_n775), .A3(new_n398), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n838), .B1(new_n839), .B2(KEYINPUT57), .ZN(new_n840));
  INV_X1    g639(.A(new_n832), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n840), .A2(new_n494), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(G141gat), .ZN(new_n843));
  AOI211_X1 g642(.A(KEYINPUT122), .B(new_n817), .C1(new_n843), .C2(new_n821), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT122), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n831), .A2(new_n647), .A3(new_n832), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n821), .B1(new_n846), .B2(new_n215), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n845), .B1(new_n847), .B2(KEYINPUT58), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n837), .B1(new_n844), .B2(new_n848), .ZN(G1344gat));
  NAND3_X1  g648(.A1(new_n820), .A2(new_n217), .A3(new_n595), .ZN(new_n850));
  AOI211_X1 g649(.A(KEYINPUT59), .B(new_n217), .C1(new_n835), .C2(new_n595), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT59), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n790), .A2(new_n824), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n499), .A2(new_n608), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n828), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g654(.A(KEYINPUT57), .B1(new_n855), .B2(new_n253), .ZN(new_n856));
  OAI211_X1 g655(.A(new_n595), .B(new_n841), .C1(new_n853), .C2(new_n856), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n852), .B1(new_n857), .B2(G148gat), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n850), .B1(new_n851), .B2(new_n858), .ZN(G1345gat));
  NAND3_X1  g658(.A1(new_n820), .A2(new_n221), .A3(new_n638), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n831), .A2(new_n607), .A3(new_n832), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n860), .B1(new_n861), .B2(new_n221), .ZN(G1346gat));
  NAND3_X1  g661(.A1(new_n820), .A2(new_n222), .A3(new_n541), .ZN(new_n863));
  NOR3_X1   g662(.A1(new_n831), .A2(new_n540), .A3(new_n832), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n863), .B1(new_n864), .B2(new_n222), .ZN(G1347gat));
  NOR2_X1   g664(.A1(new_n777), .A2(new_n391), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n776), .A2(new_n325), .A3(new_n866), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n867), .A2(new_n258), .A3(new_n499), .ZN(new_n868));
  INV_X1    g667(.A(new_n778), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n776), .A2(new_n869), .A3(new_n866), .ZN(new_n870));
  INV_X1    g669(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(new_n494), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n868), .B1(new_n872), .B2(new_n258), .ZN(G1348gat));
  OAI21_X1  g672(.A(G176gat), .B1(new_n867), .B2(new_n680), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n595), .A2(new_n259), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n874), .B1(new_n870), .B2(new_n875), .ZN(G1349gat));
  AND2_X1   g675(.A1(new_n638), .A2(new_n277), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n870), .A2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT124), .ZN(new_n880));
  AOI22_X1  g679(.A1(new_n879), .A2(new_n880), .B1(KEYINPUT125), .B2(KEYINPUT60), .ZN(new_n881));
  OAI21_X1  g680(.A(KEYINPUT124), .B1(new_n870), .B2(new_n878), .ZN(new_n882));
  OAI21_X1  g681(.A(G183gat), .B1(new_n867), .B2(new_n607), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  NOR2_X1   g683(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  XNOR2_X1  g685(.A(new_n884), .B(new_n886), .ZN(G1350gat));
  NAND3_X1  g686(.A1(new_n871), .A2(new_n278), .A3(new_n541), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT61), .ZN(new_n889));
  OR2_X1    g688(.A1(new_n867), .A2(new_n540), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n889), .B1(new_n890), .B2(G190gat), .ZN(new_n891));
  OAI211_X1 g690(.A(new_n889), .B(G190gat), .C1(new_n867), .C2(new_n540), .ZN(new_n892));
  INV_X1    g691(.A(new_n892), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n888), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(KEYINPUT126), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT126), .ZN(new_n896));
  OAI211_X1 g695(.A(new_n888), .B(new_n896), .C1(new_n891), .C2(new_n893), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n895), .A2(new_n897), .ZN(G1351gat));
  NOR2_X1   g697(.A1(new_n853), .A2(new_n856), .ZN(new_n899));
  OR2_X1    g698(.A1(new_n899), .A2(KEYINPUT127), .ZN(new_n900));
  INV_X1    g699(.A(new_n866), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n623), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n899), .A2(KEYINPUT127), .ZN(new_n903));
  INV_X1    g702(.A(G197gat), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n499), .A2(new_n904), .ZN(new_n905));
  NAND4_X1  g704(.A1(new_n900), .A2(new_n902), .A3(new_n903), .A4(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n839), .A2(new_n902), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n904), .B1(new_n907), .B2(new_n647), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n906), .A2(new_n908), .ZN(G1352gat));
  NAND3_X1  g708(.A1(new_n900), .A2(new_n902), .A3(new_n903), .ZN(new_n910));
  OAI21_X1  g709(.A(G204gat), .B1(new_n910), .B2(new_n680), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n907), .A2(G204gat), .A3(new_n680), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n912), .B(KEYINPUT62), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n911), .A2(new_n913), .ZN(G1353gat));
  OR3_X1    g713(.A1(new_n907), .A2(G211gat), .A3(new_n607), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n902), .A2(new_n638), .ZN(new_n916));
  OAI21_X1  g715(.A(G211gat), .B1(new_n899), .B2(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT63), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n917), .A2(new_n918), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n915), .B1(new_n919), .B2(new_n920), .ZN(G1354gat));
  INV_X1    g720(.A(G218gat), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n540), .A2(new_n922), .ZN(new_n923));
  NAND4_X1  g722(.A1(new_n900), .A2(new_n902), .A3(new_n903), .A4(new_n923), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n922), .B1(new_n907), .B2(new_n540), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n924), .A2(new_n925), .ZN(G1355gat));
endmodule


