//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 1 0 0 0 0 1 1 1 1 0 1 1 0 1 0 1 0 0 0 1 0 1 1 0 0 1 1 0 0 1 1 1 1 0 0 1 0 1 1 1 0 1 1 1 1 0 0 1 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:24 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n817, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n984, new_n985, new_n986, new_n987, new_n988, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061;
  INV_X1    g000(.A(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G217), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT25), .ZN(new_n189));
  AOI21_X1  g003(.A(G902), .B1(new_n189), .B2(KEYINPUT75), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT22), .B(G137), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n191), .B(KEYINPUT74), .ZN(new_n192));
  AND2_X1   g006(.A1(KEYINPUT68), .A2(G953), .ZN(new_n193));
  NOR2_X1   g007(.A1(KEYINPUT68), .A2(G953), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n195), .A2(G221), .A3(G234), .ZN(new_n196));
  XNOR2_X1  g010(.A(new_n192), .B(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT73), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT23), .ZN(new_n200));
  INV_X1    g014(.A(G119), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n200), .B1(new_n201), .B2(G128), .ZN(new_n202));
  INV_X1    g016(.A(G128), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n203), .A2(KEYINPUT23), .A3(G119), .ZN(new_n204));
  OAI211_X1 g018(.A(new_n202), .B(new_n204), .C1(G119), .C2(new_n203), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G110), .ZN(new_n206));
  XOR2_X1   g020(.A(KEYINPUT24), .B(G110), .Z(new_n207));
  XNOR2_X1  g021(.A(G119), .B(G128), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n206), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G140), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G125), .ZN(new_n212));
  INV_X1    g026(.A(G125), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G140), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n212), .A2(new_n214), .A3(KEYINPUT71), .ZN(new_n215));
  OR3_X1    g029(.A1(new_n213), .A2(KEYINPUT71), .A3(G140), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n215), .A2(new_n216), .A3(KEYINPUT16), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT16), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n212), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G146), .ZN(new_n221));
  INV_X1    g035(.A(G146), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n217), .A2(new_n222), .A3(new_n219), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n210), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  XOR2_X1   g038(.A(KEYINPUT72), .B(G110), .Z(new_n225));
  OAI22_X1  g039(.A1(new_n205), .A2(new_n225), .B1(new_n208), .B2(new_n207), .ZN(new_n226));
  AND2_X1   g040(.A1(new_n212), .A2(new_n214), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(new_n222), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n222), .B1(new_n217), .B2(new_n219), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n199), .B1(new_n224), .B2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n223), .ZN(new_n233));
  OAI211_X1 g047(.A(new_n209), .B(new_n206), .C1(new_n233), .C2(new_n230), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n221), .A2(new_n228), .A3(new_n226), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n234), .A2(KEYINPUT73), .A3(new_n235), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n198), .B1(new_n232), .B2(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n197), .B1(new_n234), .B2(new_n235), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n190), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n189), .A2(KEYINPUT75), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n188), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  OAI221_X1 g055(.A(new_n190), .B1(KEYINPUT75), .B2(new_n189), .C1(new_n237), .C2(new_n238), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  OR3_X1    g057(.A1(new_n237), .A2(KEYINPUT76), .A3(new_n238), .ZN(new_n244));
  INV_X1    g058(.A(G902), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n188), .A2(new_n245), .ZN(new_n246));
  XOR2_X1   g060(.A(new_n246), .B(KEYINPUT77), .Z(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  OAI21_X1  g062(.A(KEYINPUT76), .B1(new_n237), .B2(new_n238), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n244), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n243), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G113), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(KEYINPUT2), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT2), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G113), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g070(.A(G116), .B(G119), .ZN(new_n257));
  XNOR2_X1  g071(.A(new_n256), .B(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT11), .ZN(new_n259));
  INV_X1    g073(.A(G134), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n259), .B1(new_n260), .B2(G137), .ZN(new_n261));
  INV_X1    g075(.A(G137), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n262), .A2(KEYINPUT11), .A3(G134), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n260), .A2(G137), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n261), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G131), .ZN(new_n266));
  INV_X1    g080(.A(G131), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n261), .A2(new_n263), .A3(new_n267), .A4(new_n264), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(KEYINPUT0), .A2(G128), .ZN(new_n270));
  OR2_X1    g084(.A1(KEYINPUT0), .A2(G128), .ZN(new_n271));
  INV_X1    g085(.A(G143), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n272), .A2(G146), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n222), .A2(G143), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n270), .B(new_n271), .C1(new_n273), .C2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n222), .A2(G143), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n272), .A2(G146), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n276), .A2(new_n277), .A3(KEYINPUT0), .A4(G128), .ZN(new_n278));
  AND2_X1   g092(.A1(new_n275), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n258), .B1(new_n269), .B2(new_n279), .ZN(new_n280));
  XNOR2_X1  g094(.A(G143), .B(G146), .ZN(new_n281));
  XNOR2_X1  g095(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n281), .A2(new_n282), .A3(G128), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n222), .A2(G143), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT1), .ZN(new_n285));
  AND2_X1   g099(.A1(new_n285), .A2(KEYINPUT66), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n285), .A2(KEYINPUT66), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n284), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n203), .B1(new_n273), .B2(new_n274), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n283), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT64), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n291), .A2(new_n262), .A3(G134), .ZN(new_n292));
  OAI21_X1  g106(.A(KEYINPUT64), .B1(new_n260), .B2(G137), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n262), .A2(G134), .ZN(new_n294));
  OAI211_X1 g108(.A(G131), .B(new_n292), .C1(new_n293), .C2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n290), .A2(new_n268), .A3(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(KEYINPUT28), .B1(new_n280), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n295), .A2(new_n268), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT65), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n295), .A2(KEYINPUT65), .A3(new_n268), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n300), .A2(new_n301), .A3(new_n290), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n279), .A2(new_n269), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(new_n258), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT67), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n303), .A2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(new_n258), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n279), .A2(new_n269), .A3(KEYINPUT67), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n307), .A2(new_n308), .A3(new_n309), .A4(new_n296), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n305), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n297), .B1(new_n311), .B2(KEYINPUT28), .ZN(new_n312));
  INV_X1    g126(.A(G237), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n195), .A2(G210), .A3(new_n313), .ZN(new_n314));
  XNOR2_X1  g128(.A(new_n314), .B(KEYINPUT27), .ZN(new_n315));
  XNOR2_X1  g129(.A(KEYINPUT26), .B(G101), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n315), .B(new_n316), .ZN(new_n317));
  OR2_X1    g131(.A1(new_n312), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n309), .A2(new_n296), .ZN(new_n319));
  AOI21_X1  g133(.A(KEYINPUT67), .B1(new_n279), .B2(new_n269), .ZN(new_n320));
  NOR3_X1   g134(.A1(new_n319), .A2(new_n258), .A3(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(KEYINPUT30), .B1(new_n319), .B2(new_n320), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT30), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n302), .A2(new_n323), .A3(new_n303), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n321), .B1(new_n325), .B2(new_n258), .ZN(new_n326));
  AOI21_X1  g140(.A(KEYINPUT31), .B1(new_n326), .B2(new_n317), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n308), .B1(new_n322), .B2(new_n324), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT31), .ZN(new_n329));
  INV_X1    g143(.A(new_n317), .ZN(new_n330));
  NOR4_X1   g144(.A1(new_n328), .A2(new_n329), .A3(new_n330), .A4(new_n321), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n318), .B1(new_n327), .B2(new_n331), .ZN(new_n332));
  NOR2_X1   g146(.A1(G472), .A2(G902), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n332), .A2(KEYINPUT32), .A3(new_n333), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n330), .B1(new_n328), .B2(new_n321), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n308), .B1(new_n302), .B2(new_n303), .ZN(new_n336));
  OAI21_X1  g150(.A(KEYINPUT28), .B1(new_n321), .B2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(new_n297), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n337), .A2(new_n338), .A3(new_n317), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT29), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n335), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n258), .B1(new_n319), .B2(new_n320), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(new_n310), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n297), .B1(new_n343), .B2(KEYINPUT28), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n330), .A2(new_n340), .ZN(new_n345));
  AOI21_X1  g159(.A(G902), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n341), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n347), .A2(KEYINPUT70), .A3(G472), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n334), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(KEYINPUT70), .B1(new_n347), .B2(G472), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT69), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n312), .A2(new_n317), .ZN(new_n353));
  AND3_X1   g167(.A1(new_n302), .A2(new_n323), .A3(new_n303), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n307), .A2(new_n309), .A3(new_n296), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n354), .B1(KEYINPUT30), .B2(new_n355), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n310), .B(new_n317), .C1(new_n356), .C2(new_n308), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(new_n329), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n326), .A2(KEYINPUT31), .A3(new_n317), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n353), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n333), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n352), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n332), .A2(KEYINPUT69), .A3(new_n333), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT32), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n362), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n251), .B1(new_n351), .B2(new_n365), .ZN(new_n366));
  XNOR2_X1  g180(.A(KEYINPUT9), .B(G234), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT78), .ZN(new_n368));
  XNOR2_X1  g182(.A(new_n367), .B(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(new_n245), .ZN(new_n370));
  AND2_X1   g184(.A1(new_n370), .A2(G221), .ZN(new_n371));
  INV_X1    g185(.A(G469), .ZN(new_n372));
  XOR2_X1   g186(.A(KEYINPUT83), .B(G101), .Z(new_n373));
  INV_X1    g187(.A(G104), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n374), .A2(KEYINPUT3), .ZN(new_n375));
  OR2_X1    g189(.A1(KEYINPUT80), .A2(G107), .ZN(new_n376));
  NAND2_X1  g190(.A1(KEYINPUT80), .A2(G107), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n375), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(G107), .ZN(new_n379));
  OAI21_X1  g193(.A(KEYINPUT81), .B1(new_n379), .B2(G104), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT81), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n381), .A2(new_n374), .A3(G107), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n379), .A2(G104), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(KEYINPUT3), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n373), .A2(new_n378), .A3(new_n383), .A4(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(G104), .B1(new_n376), .B2(new_n377), .ZN(new_n387));
  INV_X1    g201(.A(new_n384), .ZN(new_n388));
  OAI21_X1  g202(.A(G101), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  AND2_X1   g203(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT84), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n390), .A2(new_n391), .A3(KEYINPUT10), .A4(new_n290), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n290), .A2(KEYINPUT10), .A3(new_n386), .A4(new_n389), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(KEYINPUT84), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n269), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n275), .A2(new_n278), .ZN(new_n397));
  INV_X1    g211(.A(G101), .ZN(new_n398));
  AOI22_X1  g212(.A1(new_n380), .A2(new_n382), .B1(new_n384), .B2(KEYINPUT3), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n398), .B1(new_n399), .B2(new_n378), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT4), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n397), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT82), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n381), .B1(new_n374), .B2(G107), .ZN(new_n404));
  NOR3_X1   g218(.A1(new_n379), .A2(KEYINPUT81), .A3(G104), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n385), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  AND3_X1   g220(.A1(new_n375), .A2(new_n376), .A3(new_n377), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n403), .B(G101), .C1(new_n406), .C2(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n408), .A2(KEYINPUT4), .A3(new_n386), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n400), .A2(new_n403), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n402), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(G128), .B1(new_n276), .B2(new_n277), .ZN(new_n412));
  NOR3_X1   g226(.A1(new_n273), .A2(new_n274), .A3(new_n203), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n412), .B1(new_n413), .B2(new_n282), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n274), .A2(KEYINPUT1), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n390), .A2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT10), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n395), .A2(new_n396), .A3(new_n411), .A4(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n195), .A2(G227), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n421), .B(KEYINPUT79), .ZN(new_n422));
  XNOR2_X1  g236(.A(G110), .B(G140), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n422), .B(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n420), .A2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT85), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT12), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n386), .A2(new_n389), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n429), .B1(new_n414), .B2(new_n415), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n290), .B1(new_n386), .B2(new_n389), .ZN(new_n431));
  OAI211_X1 g245(.A(new_n427), .B(new_n428), .C1(new_n430), .C2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(KEYINPUT86), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n417), .B1(new_n290), .B2(new_n390), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT86), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n396), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n427), .B(new_n269), .C1(new_n430), .C2(new_n431), .ZN(new_n437));
  AOI22_X1  g251(.A1(new_n433), .A2(new_n436), .B1(KEYINPUT12), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n426), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT88), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n411), .A2(new_n419), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n393), .B(new_n391), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n440), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND4_X1  g257(.A1(new_n395), .A2(KEYINPUT88), .A3(new_n411), .A4(new_n419), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n443), .A2(new_n269), .A3(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n424), .B1(new_n445), .B2(new_n420), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT89), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n439), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(new_n420), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n395), .A2(new_n411), .A3(new_n419), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n396), .B1(new_n450), .B2(new_n440), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n449), .B1(new_n451), .B2(new_n444), .ZN(new_n452));
  NOR3_X1   g266(.A1(new_n452), .A2(KEYINPUT89), .A3(new_n424), .ZN(new_n453));
  OAI211_X1 g267(.A(new_n372), .B(new_n245), .C1(new_n448), .C2(new_n453), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n372), .A2(new_n245), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n424), .B1(new_n438), .B2(new_n420), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT87), .ZN(new_n457));
  AOI22_X1  g271(.A1(new_n451), .A2(new_n444), .B1(new_n425), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n426), .A2(KEYINPUT87), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n456), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n455), .B1(new_n460), .B2(G469), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n371), .B1(new_n454), .B2(new_n461), .ZN(new_n462));
  XNOR2_X1  g276(.A(G110), .B(G122), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n463), .B(KEYINPUT8), .ZN(new_n464));
  INV_X1    g278(.A(G116), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n465), .A2(G119), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT5), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n252), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n201), .A2(G116), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n465), .A2(G119), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n469), .A2(new_n470), .A3(KEYINPUT5), .ZN(new_n471));
  AOI22_X1  g285(.A1(new_n468), .A2(new_n471), .B1(new_n257), .B2(new_n256), .ZN(new_n472));
  AND3_X1   g286(.A1(new_n472), .A2(new_n386), .A3(new_n389), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n256), .A2(new_n257), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n468), .A2(new_n471), .ZN(new_n475));
  AOI22_X1  g289(.A1(new_n386), .A2(new_n389), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n464), .B1(new_n473), .B2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT91), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  OAI211_X1 g293(.A(KEYINPUT91), .B(new_n464), .C1(new_n473), .C2(new_n476), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n290), .A2(new_n213), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n275), .A2(G125), .A3(new_n278), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT7), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n485), .A2(KEYINPUT92), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(G953), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(G224), .ZN(new_n489));
  AOI22_X1  g303(.A1(new_n484), .A2(new_n487), .B1(KEYINPUT7), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(KEYINPUT7), .ZN(new_n491));
  AOI211_X1 g305(.A(new_n491), .B(new_n486), .C1(new_n482), .C2(new_n483), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n473), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n409), .A2(new_n410), .ZN(new_n495));
  OAI211_X1 g309(.A(new_n401), .B(G101), .C1(new_n406), .C2(new_n407), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n258), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n494), .B(new_n463), .C1(new_n495), .C2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n481), .A2(new_n493), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(new_n245), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT93), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(G210), .B1(G237), .B2(G902), .ZN(new_n503));
  INV_X1    g317(.A(new_n463), .ZN(new_n504));
  AOI211_X1 g318(.A(KEYINPUT82), .B(new_n398), .C1(new_n399), .C2(new_n378), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n386), .A2(KEYINPUT4), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n410), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n497), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n504), .B1(new_n509), .B2(new_n473), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n510), .A2(KEYINPUT6), .A3(new_n498), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT6), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n512), .B(new_n504), .C1(new_n509), .C2(new_n473), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n484), .B(new_n489), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n511), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n499), .A2(KEYINPUT93), .A3(new_n245), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n502), .A2(new_n503), .A3(new_n515), .A4(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT94), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AND2_X1   g333(.A1(new_n515), .A2(new_n516), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n520), .A2(KEYINPUT94), .A3(new_n503), .A4(new_n502), .ZN(new_n521));
  INV_X1    g335(.A(new_n503), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n515), .A2(new_n516), .ZN(new_n523));
  AOI21_X1  g337(.A(KEYINPUT93), .B1(new_n499), .B2(new_n245), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n519), .A2(new_n521), .A3(new_n525), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n233), .A2(new_n230), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT68), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(new_n488), .ZN(new_n529));
  NAND2_X1  g343(.A1(KEYINPUT68), .A2(G953), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n529), .A2(G214), .A3(new_n313), .A4(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(new_n272), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n195), .A2(G143), .A3(G214), .A4(new_n313), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n267), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(KEYINPUT17), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n532), .A2(new_n533), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(G131), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n532), .A2(new_n533), .A3(new_n267), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  OAI211_X1 g353(.A(new_n527), .B(new_n535), .C1(new_n539), .C2(KEYINPUT17), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT18), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n532), .B(new_n533), .C1(new_n541), .C2(new_n267), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n215), .A2(new_n216), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n228), .B1(new_n543), .B2(new_n222), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT95), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n541), .A2(new_n267), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n536), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n547), .B1(new_n536), .B2(new_n548), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n546), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  XNOR2_X1  g366(.A(G113), .B(G122), .ZN(new_n553));
  XNOR2_X1  g367(.A(KEYINPUT96), .B(G104), .ZN(new_n554));
  XOR2_X1   g368(.A(new_n553), .B(new_n554), .Z(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n540), .A2(new_n552), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(KEYINPUT98), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n556), .B1(new_n540), .B2(new_n552), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n540), .A2(new_n552), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT98), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n561), .A2(new_n562), .A3(new_n555), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(new_n245), .ZN(new_n564));
  OAI21_X1  g378(.A(G475), .B1(new_n560), .B2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT99), .ZN(new_n566));
  INV_X1    g380(.A(G122), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(G116), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n465), .A2(G122), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n376), .A2(new_n568), .A3(new_n569), .A4(new_n377), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  AOI22_X1  g385(.A1(new_n568), .A2(new_n569), .B1(new_n376), .B2(new_n377), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n566), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n272), .A2(G128), .ZN(new_n574));
  OAI21_X1  g388(.A(G134), .B1(new_n574), .B2(KEYINPUT13), .ZN(new_n575));
  XOR2_X1   g389(.A(G128), .B(G143), .Z(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(G128), .B(G143), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n578), .B(G134), .C1(KEYINPUT13), .C2(new_n574), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n568), .A2(new_n569), .ZN(new_n581));
  XNOR2_X1  g395(.A(KEYINPUT80), .B(G107), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n583), .A2(KEYINPUT99), .A3(new_n570), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n573), .A2(new_n580), .A3(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n465), .A2(KEYINPUT14), .A3(G122), .ZN(new_n586));
  OAI211_X1 g400(.A(G107), .B(new_n586), .C1(new_n581), .C2(KEYINPUT14), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n576), .A2(new_n260), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n578), .A2(G134), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n587), .A2(new_n570), .A3(new_n588), .A4(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n585), .A2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(G217), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n592), .A2(G953), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n369), .A2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n585), .A2(new_n594), .A3(new_n590), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n596), .A2(new_n245), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(KEYINPUT100), .ZN(new_n599));
  INV_X1    g413(.A(G478), .ZN(new_n600));
  NOR2_X1   g414(.A1(KEYINPUT101), .A2(KEYINPUT15), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(KEYINPUT101), .A2(KEYINPUT15), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n600), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT100), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n596), .A2(new_n605), .A3(new_n245), .A4(new_n597), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n599), .A2(new_n604), .A3(new_n606), .ZN(new_n607));
  OR2_X1    g421(.A1(new_n598), .A2(new_n604), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT20), .ZN(new_n611));
  NOR2_X1   g425(.A1(G475), .A2(G902), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT97), .ZN(new_n613));
  AND2_X1   g427(.A1(new_n531), .A2(new_n272), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n531), .A2(new_n272), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n548), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(KEYINPUT95), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n545), .B1(new_n617), .B2(new_n549), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT19), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n619), .B1(new_n215), .B2(new_n216), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n227), .A2(KEYINPUT19), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n222), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  AND3_X1   g436(.A1(new_n532), .A2(new_n533), .A3(new_n267), .ZN(new_n623));
  OAI211_X1 g437(.A(new_n221), .B(new_n622), .C1(new_n623), .C2(new_n534), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  OAI211_X1 g439(.A(new_n613), .B(new_n555), .C1(new_n618), .C2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(new_n557), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n552), .A2(new_n624), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n613), .B1(new_n628), .B2(new_n555), .ZN(new_n629));
  OAI211_X1 g443(.A(new_n611), .B(new_n612), .C1(new_n627), .C2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n617), .A2(new_n549), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n543), .A2(KEYINPUT19), .ZN(new_n633));
  OR2_X1    g447(.A1(new_n227), .A2(KEYINPUT19), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n230), .B1(new_n635), .B2(new_n222), .ZN(new_n636));
  AOI22_X1  g450(.A1(new_n632), .A2(new_n546), .B1(new_n539), .B2(new_n636), .ZN(new_n637));
  OAI21_X1  g451(.A(KEYINPUT97), .B1(new_n637), .B2(new_n556), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n638), .A2(new_n557), .A3(new_n626), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n611), .B1(new_n639), .B2(new_n612), .ZN(new_n640));
  OAI211_X1 g454(.A(new_n565), .B(new_n610), .C1(new_n631), .C2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(G952), .ZN(new_n642));
  AOI211_X1 g456(.A(G953), .B(new_n642), .C1(G234), .C2(G237), .ZN(new_n643));
  AOI211_X1 g457(.A(new_n245), .B(new_n195), .C1(G234), .C2(G237), .ZN(new_n644));
  XNOR2_X1  g458(.A(KEYINPUT21), .B(G898), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n643), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n641), .A2(new_n646), .ZN(new_n647));
  OAI21_X1  g461(.A(G214), .B1(G237), .B2(G902), .ZN(new_n648));
  XOR2_X1   g462(.A(new_n648), .B(KEYINPUT90), .Z(new_n649));
  AND3_X1   g463(.A1(new_n526), .A2(new_n647), .A3(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n366), .A2(new_n462), .A3(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(new_n651), .B(new_n373), .Z(G3));
  NAND2_X1  g466(.A1(new_n525), .A2(new_n517), .ZN(new_n653));
  INV_X1    g467(.A(new_n646), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n653), .A2(new_n648), .A3(new_n654), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n565), .B1(new_n631), .B2(new_n640), .ZN(new_n656));
  AND2_X1   g470(.A1(new_n594), .A2(KEYINPUT103), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n591), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n594), .A2(KEYINPUT103), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n659), .A2(new_n585), .A3(new_n590), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n658), .A2(KEYINPUT33), .A3(new_n660), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT102), .B(KEYINPUT33), .Z(new_n662));
  NAND3_X1  g476(.A1(new_n596), .A2(new_n597), .A3(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n600), .A2(G902), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n661), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT104), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n599), .A2(new_n600), .A3(new_n606), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n661), .A2(new_n663), .A3(KEYINPUT104), .A4(new_n664), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(KEYINPUT105), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT105), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n667), .A2(new_n668), .A3(new_n672), .A4(new_n669), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n656), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(KEYINPUT106), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n612), .B1(new_n627), .B2(new_n629), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(KEYINPUT20), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(new_n630), .ZN(new_n679));
  AOI22_X1  g493(.A1(new_n679), .A2(new_n565), .B1(new_n671), .B2(new_n673), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT106), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n655), .B1(new_n676), .B2(new_n682), .ZN(new_n683));
  OAI21_X1  g497(.A(G472), .B1(new_n360), .B2(G902), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n362), .A2(new_n684), .A3(new_n363), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n685), .A2(new_n251), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n683), .A2(new_n462), .A3(new_n686), .ZN(new_n687));
  XOR2_X1   g501(.A(KEYINPUT34), .B(G104), .Z(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G6));
  OR2_X1    g503(.A1(new_n558), .A2(new_n559), .ZN(new_n690));
  AOI21_X1  g504(.A(G902), .B1(new_n558), .B2(new_n559), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AOI22_X1  g506(.A1(new_n678), .A2(new_n630), .B1(new_n692), .B2(G475), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n609), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n655), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n686), .A2(new_n695), .A3(new_n462), .ZN(new_n696));
  XOR2_X1   g510(.A(KEYINPUT35), .B(G107), .Z(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(G9));
  NAND2_X1  g512(.A1(new_n232), .A2(new_n236), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT36), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n699), .A2(new_n700), .A3(new_n198), .ZN(new_n701));
  OAI211_X1 g515(.A(new_n232), .B(new_n236), .C1(KEYINPUT36), .C2(new_n197), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  AOI22_X1  g518(.A1(new_n241), .A2(new_n242), .B1(new_n704), .B2(new_n248), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n685), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n650), .A2(new_n462), .A3(new_n706), .ZN(new_n707));
  XOR2_X1   g521(.A(KEYINPUT37), .B(G110), .Z(new_n708));
  XNOR2_X1  g522(.A(new_n707), .B(new_n708), .ZN(G12));
  INV_X1    g523(.A(new_n648), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n710), .B1(new_n525), .B2(new_n517), .ZN(new_n711));
  INV_X1    g525(.A(new_n705), .ZN(new_n712));
  AND3_X1   g526(.A1(new_n362), .A2(new_n364), .A3(new_n363), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n347), .A2(G472), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT70), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n716), .A2(new_n334), .A3(new_n348), .ZN(new_n717));
  OAI211_X1 g531(.A(new_n711), .B(new_n712), .C1(new_n713), .C2(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(G900), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n644), .A2(new_n719), .ZN(new_n720));
  OR2_X1    g534(.A1(new_n720), .A2(KEYINPUT107), .ZN(new_n721));
  INV_X1    g535(.A(new_n643), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n720), .A2(KEYINPUT107), .ZN(new_n723));
  AND3_X1   g537(.A1(new_n721), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n694), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n462), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n718), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(new_n203), .ZN(G30));
  OAI21_X1  g542(.A(new_n317), .B1(new_n328), .B2(new_n321), .ZN(new_n729));
  INV_X1    g543(.A(new_n729), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n245), .B1(new_n343), .B2(new_n317), .ZN(new_n731));
  OAI21_X1  g545(.A(G472), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  AND2_X1   g546(.A1(new_n334), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n365), .A2(new_n733), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n610), .B1(new_n679), .B2(new_n565), .ZN(new_n735));
  AND4_X1   g549(.A1(new_n648), .A2(new_n734), .A3(new_n705), .A4(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n526), .B(KEYINPUT38), .ZN(new_n737));
  XOR2_X1   g551(.A(new_n724), .B(KEYINPUT39), .Z(new_n738));
  NAND2_X1  g552(.A1(new_n462), .A2(new_n738), .ZN(new_n739));
  OAI211_X1 g553(.A(new_n736), .B(new_n737), .C1(KEYINPUT40), .C2(new_n739), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n740), .B1(KEYINPUT40), .B2(new_n739), .ZN(new_n741));
  XOR2_X1   g555(.A(KEYINPUT108), .B(G143), .Z(new_n742));
  XNOR2_X1  g556(.A(new_n741), .B(new_n742), .ZN(G45));
  NAND2_X1  g557(.A1(new_n653), .A2(new_n648), .ZN(new_n744));
  AOI211_X1 g558(.A(new_n744), .B(new_n705), .C1(new_n351), .C2(new_n365), .ZN(new_n745));
  INV_X1    g559(.A(new_n724), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n656), .A2(new_n674), .A3(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT109), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n680), .A2(KEYINPUT109), .A3(new_n746), .ZN(new_n750));
  AND3_X1   g564(.A1(new_n462), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n745), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G146), .ZN(G48));
  INV_X1    g567(.A(new_n454), .ZN(new_n754));
  OAI21_X1  g568(.A(KEYINPUT89), .B1(new_n452), .B2(new_n424), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n445), .A2(new_n420), .ZN(new_n756));
  INV_X1    g570(.A(new_n424), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n756), .A2(new_n447), .A3(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n755), .A2(new_n758), .A3(new_n439), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n372), .B1(new_n759), .B2(new_n245), .ZN(new_n760));
  NOR3_X1   g574(.A1(new_n754), .A2(new_n760), .A3(new_n371), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n366), .A2(new_n761), .A3(new_n683), .ZN(new_n762));
  XNOR2_X1  g576(.A(KEYINPUT41), .B(G113), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n762), .B(new_n763), .ZN(G15));
  NAND3_X1  g578(.A1(new_n366), .A2(new_n761), .A3(new_n695), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G116), .ZN(G18));
  AOI21_X1  g580(.A(new_n705), .B1(new_n351), .B2(new_n365), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n767), .A2(new_n761), .A3(new_n647), .A4(new_n711), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G119), .ZN(G21));
  NAND2_X1  g583(.A1(new_n358), .A2(new_n359), .ZN(new_n770));
  OR2_X1    g584(.A1(new_n344), .A2(new_n317), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n361), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n243), .A2(KEYINPUT110), .A3(new_n250), .ZN(new_n774));
  INV_X1    g588(.A(new_n774), .ZN(new_n775));
  AOI21_X1  g589(.A(KEYINPUT110), .B1(new_n243), .B2(new_n250), .ZN(new_n776));
  OAI211_X1 g590(.A(new_n684), .B(new_n773), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n711), .A2(new_n735), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n779), .A2(new_n646), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n761), .A2(new_n778), .A3(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G122), .ZN(G24));
  NAND2_X1  g596(.A1(new_n759), .A2(new_n245), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(G469), .ZN(new_n784));
  INV_X1    g598(.A(new_n371), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n784), .A2(new_n785), .A3(new_n454), .A4(new_n711), .ZN(new_n786));
  INV_X1    g600(.A(G472), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n787), .B1(new_n332), .B2(new_n245), .ZN(new_n788));
  NOR3_X1   g602(.A1(new_n788), .A2(new_n772), .A3(new_n705), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n749), .A2(new_n750), .A3(new_n789), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n786), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(new_n213), .ZN(G27));
  INV_X1    g606(.A(new_n776), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(new_n774), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n364), .B1(new_n360), .B2(new_n361), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n716), .A2(new_n795), .A3(new_n334), .A4(new_n348), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n749), .A2(new_n794), .A3(new_n750), .A4(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n502), .A2(new_n515), .A3(new_n516), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n710), .B1(new_n798), .B2(new_n522), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n799), .A2(new_n519), .A3(new_n521), .ZN(new_n800));
  INV_X1    g614(.A(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n454), .A2(new_n461), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n801), .A2(new_n802), .A3(new_n785), .ZN(new_n803));
  OAI21_X1  g617(.A(KEYINPUT42), .B1(new_n797), .B2(new_n803), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n799), .A2(new_n519), .A3(new_n521), .A4(new_n785), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n805), .B1(new_n454), .B2(new_n461), .ZN(new_n806));
  AOI21_X1  g620(.A(KEYINPUT109), .B1(new_n680), .B2(new_n746), .ZN(new_n807));
  AND4_X1   g621(.A1(KEYINPUT109), .A2(new_n656), .A3(new_n674), .A4(new_n746), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT42), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n366), .A2(new_n806), .A3(new_n809), .A4(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT111), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n804), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n812), .B1(new_n804), .B2(new_n811), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(G131), .ZN(G33));
  NAND3_X1  g630(.A1(new_n366), .A2(new_n806), .A3(new_n725), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(G134), .ZN(G36));
  NAND2_X1  g632(.A1(new_n685), .A2(new_n712), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(KEYINPUT113), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n656), .B1(new_n673), .B2(new_n671), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n821), .B1(KEYINPUT112), .B2(KEYINPUT43), .ZN(new_n822));
  XNOR2_X1  g636(.A(KEYINPUT112), .B(KEYINPUT43), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  OR2_X1    g638(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n820), .A2(KEYINPUT44), .A3(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(new_n826), .ZN(new_n827));
  OAI21_X1  g641(.A(KEYINPUT114), .B1(new_n827), .B2(new_n800), .ZN(new_n828));
  AOI21_X1  g642(.A(KEYINPUT44), .B1(new_n820), .B2(new_n825), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n460), .A2(KEYINPUT45), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n830), .A2(new_n372), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n460), .A2(KEYINPUT45), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n455), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n833), .A2(KEYINPUT46), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n454), .B1(new_n833), .B2(KEYINPUT46), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n785), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(new_n738), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n829), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT114), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n826), .A2(new_n839), .A3(new_n801), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n828), .A2(new_n838), .A3(new_n840), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n841), .B(G137), .ZN(G39));
  NAND4_X1  g656(.A1(new_n365), .A2(new_n716), .A3(new_n334), .A4(new_n348), .ZN(new_n843));
  INV_X1    g657(.A(new_n843), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n809), .A2(new_n844), .A3(new_n251), .A4(new_n801), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT47), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n836), .A2(new_n846), .ZN(new_n847));
  OAI211_X1 g661(.A(KEYINPUT47), .B(new_n785), .C1(new_n834), .C2(new_n835), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n845), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n849), .B(new_n211), .ZN(G42));
  INV_X1    g664(.A(KEYINPUT52), .ZN(new_n851));
  INV_X1    g665(.A(new_n726), .ZN(new_n852));
  INV_X1    g666(.A(new_n786), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n749), .A2(new_n750), .A3(new_n789), .ZN(new_n854));
  AOI22_X1  g668(.A1(new_n745), .A2(new_n852), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n704), .A2(new_n248), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n243), .A2(new_n856), .A3(new_n746), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n711), .A2(new_n735), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n858), .B1(new_n365), .B2(new_n733), .ZN(new_n859));
  AOI22_X1  g673(.A1(new_n745), .A2(new_n751), .B1(new_n462), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(KEYINPUT116), .B1(new_n855), .B2(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n462), .A2(new_n749), .A3(new_n750), .ZN(new_n862));
  INV_X1    g676(.A(new_n858), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(new_n734), .ZN(new_n864));
  INV_X1    g678(.A(new_n462), .ZN(new_n865));
  OAI22_X1  g679(.A1(new_n718), .A2(new_n862), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  OAI22_X1  g680(.A1(new_n718), .A2(new_n726), .B1(new_n786), .B2(new_n790), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT116), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n851), .B1(new_n861), .B2(new_n869), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n693), .A2(KEYINPUT115), .A3(new_n610), .A4(new_n746), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT115), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n872), .B1(new_n641), .B2(new_n724), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  AOI22_X1  g688(.A1(new_n767), .A2(new_n874), .B1(new_n809), .B2(new_n789), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n817), .B1(new_n875), .B2(new_n803), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n768), .A2(new_n762), .A3(new_n765), .A4(new_n781), .ZN(new_n877));
  AND2_X1   g691(.A1(new_n526), .A2(new_n649), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n646), .B1(new_n694), .B2(new_n675), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n686), .A2(new_n878), .A3(new_n462), .A4(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n651), .A2(new_n707), .A3(new_n880), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n876), .A2(new_n877), .A3(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n855), .A2(new_n860), .A3(KEYINPUT116), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n868), .B1(new_n866), .B2(new_n867), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n883), .A2(new_n884), .A3(KEYINPUT52), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n870), .A2(new_n815), .A3(new_n882), .A4(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(KEYINPUT53), .ZN(new_n887));
  AOI21_X1  g701(.A(KEYINPUT52), .B1(new_n883), .B2(new_n884), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n851), .B1(new_n855), .B2(new_n860), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n843), .A2(new_n874), .A3(new_n712), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n803), .B1(new_n891), .B2(new_n790), .ZN(new_n892));
  INV_X1    g706(.A(new_n817), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n881), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  AND4_X1   g708(.A1(new_n762), .A2(new_n768), .A3(new_n765), .A4(new_n781), .ZN(new_n895));
  AND3_X1   g709(.A1(new_n815), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT53), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n890), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n887), .A2(new_n898), .A3(KEYINPUT54), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n885), .A2(new_n882), .A3(new_n815), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n897), .B1(new_n900), .B2(new_n888), .ZN(new_n901));
  AND3_X1   g715(.A1(new_n804), .A2(new_n811), .A3(KEYINPUT53), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n894), .A2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n895), .A2(KEYINPUT117), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT117), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n877), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(new_n889), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n904), .A2(new_n908), .A3(new_n870), .A4(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n901), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n899), .B1(KEYINPUT54), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n825), .A2(new_n643), .ZN(new_n913));
  INV_X1    g727(.A(new_n761), .ZN(new_n914));
  NOR3_X1   g728(.A1(new_n913), .A2(new_n914), .A3(new_n777), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n737), .A2(new_n648), .ZN(new_n916));
  AOI21_X1  g730(.A(KEYINPUT50), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n915), .A2(KEYINPUT50), .A3(new_n916), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n761), .A2(new_n801), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n913), .A2(new_n920), .ZN(new_n921));
  AOI22_X1  g735(.A1(new_n918), .A2(new_n919), .B1(new_n789), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n847), .A2(new_n848), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n784), .A2(new_n454), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n924), .A2(new_n785), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n913), .A2(new_n777), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(new_n801), .ZN(new_n928));
  OR2_X1    g742(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n251), .A2(new_n722), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n365), .A2(new_n733), .A3(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT118), .ZN(new_n932));
  OR3_X1    g746(.A1(new_n920), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n932), .B1(new_n920), .B2(new_n931), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n656), .A2(new_n674), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n922), .A2(new_n929), .A3(KEYINPUT51), .A4(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT51), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n921), .A2(new_n789), .ZN(new_n939));
  INV_X1    g753(.A(new_n919), .ZN(new_n940));
  OAI211_X1 g754(.A(new_n936), .B(new_n939), .C1(new_n940), .C2(new_n917), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n926), .A2(new_n928), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n938), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  AOI211_X1 g757(.A(new_n642), .B(G953), .C1(new_n927), .C2(new_n853), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n676), .A2(new_n682), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n933), .A2(new_n945), .A3(new_n934), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n794), .A2(new_n796), .ZN(new_n947));
  NOR3_X1   g761(.A1(new_n913), .A2(new_n920), .A3(new_n947), .ZN(new_n948));
  XNOR2_X1  g762(.A(KEYINPUT119), .B(KEYINPUT48), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n948), .A2(new_n949), .ZN(new_n951));
  OAI211_X1 g765(.A(new_n944), .B(new_n946), .C1(new_n950), .C2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n937), .A2(new_n943), .A3(new_n953), .ZN(new_n954));
  OAI22_X1  g768(.A1(new_n912), .A2(new_n954), .B1(G952), .B2(G953), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n924), .B(KEYINPUT49), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n794), .A2(new_n821), .A3(new_n785), .A4(new_n649), .ZN(new_n957));
  OR4_X1    g771(.A1(new_n737), .A2(new_n956), .A3(new_n734), .A4(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n955), .A2(new_n958), .ZN(G75));
  NAND2_X1  g773(.A1(new_n511), .A2(new_n513), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(new_n514), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n961), .B(KEYINPUT55), .Z(new_n962));
  INV_X1    g776(.A(G210), .ZN(new_n963));
  AOI211_X1 g777(.A(new_n963), .B(new_n245), .C1(new_n901), .C2(new_n910), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n962), .B1(new_n964), .B2(KEYINPUT56), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT56), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n962), .B(KEYINPUT120), .Z(new_n967));
  NAND2_X1  g781(.A1(new_n911), .A2(G902), .ZN(new_n968));
  OAI211_X1 g782(.A(new_n966), .B(new_n967), .C1(new_n968), .C2(new_n963), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n195), .A2(G952), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(KEYINPUT121), .ZN(new_n971));
  AND3_X1   g785(.A1(new_n965), .A2(new_n969), .A3(new_n971), .ZN(G51));
  XNOR2_X1  g786(.A(new_n455), .B(KEYINPUT57), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT54), .ZN(new_n974));
  AND3_X1   g788(.A1(new_n901), .A2(new_n974), .A3(new_n910), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n974), .B1(new_n901), .B2(new_n910), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n973), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(new_n759), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n903), .B1(new_n907), .B2(new_n905), .ZN(new_n979));
  AOI22_X1  g793(.A1(new_n886), .A2(new_n897), .B1(new_n979), .B2(new_n890), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n980), .A2(new_n245), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n981), .A2(new_n832), .A3(new_n831), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n970), .B1(new_n978), .B2(new_n982), .ZN(G54));
  NAND2_X1  g797(.A1(KEYINPUT58), .A2(G475), .ZN(new_n984));
  INV_X1    g798(.A(new_n984), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n639), .B1(new_n981), .B2(new_n985), .ZN(new_n986));
  INV_X1    g800(.A(new_n639), .ZN(new_n987));
  NOR3_X1   g801(.A1(new_n968), .A2(new_n987), .A3(new_n984), .ZN(new_n988));
  NOR3_X1   g802(.A1(new_n986), .A2(new_n988), .A3(new_n970), .ZN(G60));
  AND2_X1   g803(.A1(new_n661), .A2(new_n663), .ZN(new_n990));
  XNOR2_X1  g804(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n600), .A2(new_n245), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n991), .B(new_n992), .ZN(new_n993));
  OAI211_X1 g807(.A(new_n990), .B(new_n993), .C1(new_n975), .C2(new_n976), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n994), .A2(new_n971), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n990), .B1(new_n912), .B2(new_n993), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n995), .A2(new_n996), .ZN(G63));
  INV_X1    g811(.A(KEYINPUT61), .ZN(new_n998));
  XNOR2_X1  g812(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n592), .A2(new_n245), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n999), .B(new_n1000), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n911), .A2(new_n704), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1002), .A2(new_n971), .ZN(new_n1003));
  INV_X1    g817(.A(new_n1001), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n1004), .B1(new_n901), .B2(new_n910), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n244), .A2(new_n249), .ZN(new_n1006));
  INV_X1    g820(.A(new_n1006), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n998), .B1(new_n1003), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g823(.A(KEYINPUT124), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n1010), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1011));
  INV_X1    g825(.A(new_n971), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1012), .B1(new_n1005), .B2(new_n704), .ZN(new_n1013));
  OAI211_X1 g827(.A(KEYINPUT124), .B(new_n1006), .C1(new_n980), .C2(new_n1004), .ZN(new_n1014));
  NAND4_X1  g828(.A1(new_n1011), .A2(new_n1013), .A3(KEYINPUT61), .A4(new_n1014), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1009), .A2(new_n1015), .ZN(G66));
  OR2_X1    g830(.A1(new_n877), .A2(new_n881), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1017), .A2(new_n195), .ZN(new_n1018));
  INV_X1    g832(.A(G224), .ZN(new_n1019));
  OAI21_X1  g833(.A(G953), .B1(new_n645), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n960), .B1(G898), .B2(new_n195), .ZN(new_n1022));
  XOR2_X1   g836(.A(new_n1022), .B(KEYINPUT125), .Z(new_n1023));
  XNOR2_X1  g837(.A(new_n1021), .B(new_n1023), .ZN(G69));
  NAND2_X1  g838(.A1(new_n855), .A2(new_n752), .ZN(new_n1025));
  OR3_X1    g839(.A1(new_n741), .A2(KEYINPUT62), .A3(new_n1025), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n800), .B1(new_n675), .B2(new_n694), .ZN(new_n1027));
  AND4_X1   g841(.A1(new_n366), .A2(new_n462), .A3(new_n738), .A4(new_n1027), .ZN(new_n1028));
  NOR2_X1   g842(.A1(new_n849), .A2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g843(.A(KEYINPUT62), .B1(new_n741), .B2(new_n1025), .ZN(new_n1030));
  NAND4_X1  g844(.A1(new_n1026), .A2(new_n1029), .A3(new_n841), .A4(new_n1030), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1031), .A2(new_n195), .ZN(new_n1032));
  XNOR2_X1  g846(.A(new_n356), .B(new_n635), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g848(.A(new_n195), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n1033), .B1(G900), .B2(new_n1035), .ZN(new_n1036));
  NOR4_X1   g850(.A1(new_n836), .A2(new_n837), .A3(new_n779), .A4(new_n947), .ZN(new_n1037));
  NAND3_X1  g851(.A1(new_n855), .A2(new_n752), .A3(new_n817), .ZN(new_n1038));
  NOR3_X1   g852(.A1(new_n849), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  NAND3_X1  g853(.A1(new_n1039), .A2(new_n815), .A3(new_n841), .ZN(new_n1040));
  OAI21_X1  g854(.A(new_n1036), .B1(new_n1040), .B2(new_n1035), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n1034), .A2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g856(.A(new_n195), .B1(G227), .B2(G900), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g858(.A(new_n1043), .ZN(new_n1045));
  NAND3_X1  g859(.A1(new_n1034), .A2(new_n1045), .A3(new_n1041), .ZN(new_n1046));
  NAND2_X1  g860(.A1(new_n1044), .A2(new_n1046), .ZN(G72));
  XNOR2_X1  g861(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1048));
  NOR2_X1   g862(.A1(new_n787), .A2(new_n245), .ZN(new_n1049));
  XNOR2_X1  g863(.A(new_n1048), .B(new_n1049), .ZN(new_n1050));
  OAI21_X1  g864(.A(new_n1050), .B1(new_n1031), .B2(new_n1017), .ZN(new_n1051));
  AOI21_X1  g865(.A(new_n970), .B1(new_n1051), .B2(new_n730), .ZN(new_n1052));
  NAND2_X1  g866(.A1(new_n357), .A2(new_n335), .ZN(new_n1053));
  NAND4_X1  g867(.A1(new_n887), .A2(new_n898), .A3(new_n1050), .A4(new_n1053), .ZN(new_n1054));
  NAND2_X1  g868(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g869(.A1(new_n326), .A2(new_n330), .ZN(new_n1056));
  OAI21_X1  g870(.A(new_n1050), .B1(new_n1040), .B2(new_n1017), .ZN(new_n1057));
  INV_X1    g871(.A(KEYINPUT127), .ZN(new_n1058));
  NAND2_X1  g872(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  OAI211_X1 g873(.A(KEYINPUT127), .B(new_n1050), .C1(new_n1040), .C2(new_n1017), .ZN(new_n1060));
  AOI21_X1  g874(.A(new_n1056), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NOR2_X1   g875(.A1(new_n1055), .A2(new_n1061), .ZN(G57));
endmodule


