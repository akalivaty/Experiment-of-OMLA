

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U549 ( .A(G2105), .ZN(n551) );
  NOR2_X1 U550 ( .A1(G2104), .A2(n551), .ZN(n1011) );
  BUF_X1 U551 ( .A(n1016), .Z(n519) );
  XNOR2_X1 U552 ( .A(n549), .B(KEYINPUT65), .ZN(n1016) );
  AND2_X1 U553 ( .A1(n727), .A2(n726), .ZN(n728) );
  NOR2_X1 U554 ( .A1(n705), .A2(n995), .ZN(n694) );
  INV_X1 U555 ( .A(n695), .ZN(n741) );
  AND2_X2 U556 ( .A1(G160), .A2(n687), .ZN(n695) );
  NOR2_X1 U557 ( .A1(n709), .A2(n708), .ZN(n711) );
  INV_X1 U558 ( .A(KEYINPUT95), .ZN(n710) );
  INV_X1 U559 ( .A(G2104), .ZN(n541) );
  XNOR2_X1 U560 ( .A(KEYINPUT96), .B(KEYINPUT30), .ZN(n520) );
  NAND2_X1 U561 ( .A1(n895), .A2(n794), .ZN(n521) );
  AND2_X1 U562 ( .A1(G125), .A2(n1011), .ZN(n522) );
  NOR2_X1 U563 ( .A1(n761), .A2(n804), .ZN(n523) );
  XOR2_X1 U564 ( .A(n764), .B(KEYINPUT100), .Z(n524) );
  AND2_X1 U565 ( .A1(G1996), .A2(n695), .ZN(n689) );
  NAND2_X1 U566 ( .A1(n731), .A2(n730), .ZN(n733) );
  INV_X1 U567 ( .A(KEYINPUT98), .ZN(n739) );
  XNOR2_X1 U568 ( .A(n748), .B(KEYINPUT32), .ZN(n755) );
  NAND2_X1 U569 ( .A1(n741), .A2(G8), .ZN(n804) );
  NOR2_X1 U570 ( .A1(n521), .A2(n796), .ZN(n797) );
  NAND2_X1 U571 ( .A1(n541), .A2(n551), .ZN(n542) );
  NOR2_X1 U572 ( .A1(n552), .A2(n522), .ZN(n553) );
  NOR2_X1 U573 ( .A1(n539), .A2(n538), .ZN(n540) );
  AND2_X1 U574 ( .A1(n554), .A2(n553), .ZN(n555) );
  INV_X1 U575 ( .A(G651), .ZN(n529) );
  NOR2_X1 U576 ( .A1(G543), .A2(n529), .ZN(n525) );
  XOR2_X1 U577 ( .A(KEYINPUT1), .B(n525), .Z(n653) );
  NAND2_X1 U578 ( .A1(G63), .A2(n653), .ZN(n527) );
  XOR2_X1 U579 ( .A(KEYINPUT0), .B(G543), .Z(n530) );
  NOR2_X2 U580 ( .A1(G651), .A2(n530), .ZN(n654) );
  NAND2_X1 U581 ( .A1(G51), .A2(n654), .ZN(n526) );
  NAND2_X1 U582 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U583 ( .A(KEYINPUT6), .B(n528), .ZN(n539) );
  NOR2_X1 U584 ( .A1(n530), .A2(n529), .ZN(n650) );
  NAND2_X1 U585 ( .A1(n650), .A2(G76), .ZN(n531) );
  XNOR2_X1 U586 ( .A(n531), .B(KEYINPUT76), .ZN(n535) );
  XOR2_X1 U587 ( .A(KEYINPUT4), .B(KEYINPUT75), .Z(n533) );
  NOR2_X1 U588 ( .A1(G651), .A2(G543), .ZN(n649) );
  NAND2_X1 U589 ( .A1(G89), .A2(n649), .ZN(n532) );
  XNOR2_X1 U590 ( .A(n533), .B(n532), .ZN(n534) );
  NAND2_X1 U591 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U592 ( .A(KEYINPUT77), .B(n536), .ZN(n537) );
  XNOR2_X1 U593 ( .A(KEYINPUT5), .B(n537), .ZN(n538) );
  XOR2_X1 U594 ( .A(KEYINPUT7), .B(n540), .Z(G168) );
  XNOR2_X2 U595 ( .A(n542), .B(KEYINPUT17), .ZN(n1015) );
  NAND2_X1 U596 ( .A1(G137), .A2(n1015), .ZN(n545) );
  NAND2_X1 U597 ( .A1(G2104), .A2(G2105), .ZN(n543) );
  XOR2_X2 U598 ( .A(KEYINPUT66), .B(n543), .Z(n1012) );
  NAND2_X1 U599 ( .A1(G113), .A2(n1012), .ZN(n544) );
  NAND2_X1 U600 ( .A1(n545), .A2(n544), .ZN(n546) );
  OR2_X1 U601 ( .A1(n546), .A2(KEYINPUT67), .ZN(n548) );
  NAND2_X1 U602 ( .A1(n546), .A2(KEYINPUT67), .ZN(n547) );
  NAND2_X1 U603 ( .A1(n548), .A2(n547), .ZN(n554) );
  NAND2_X1 U604 ( .A1(n551), .A2(G2104), .ZN(n549) );
  NAND2_X1 U605 ( .A1(G101), .A2(n1016), .ZN(n550) );
  XNOR2_X1 U606 ( .A(KEYINPUT23), .B(n550), .ZN(n552) );
  XNOR2_X2 U607 ( .A(n555), .B(KEYINPUT64), .ZN(G160) );
  XOR2_X1 U608 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U609 ( .A1(G138), .A2(n1015), .ZN(n557) );
  NAND2_X1 U610 ( .A1(G102), .A2(n1016), .ZN(n556) );
  NAND2_X1 U611 ( .A1(n557), .A2(n556), .ZN(n561) );
  NAND2_X1 U612 ( .A1(n1011), .A2(G126), .ZN(n559) );
  NAND2_X1 U613 ( .A1(G114), .A2(n1012), .ZN(n558) );
  NAND2_X1 U614 ( .A1(n559), .A2(n558), .ZN(n560) );
  NOR2_X1 U615 ( .A1(n561), .A2(n560), .ZN(G164) );
  AND2_X1 U616 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U617 ( .A(G57), .ZN(G237) );
  INV_X1 U618 ( .A(G132), .ZN(G219) );
  INV_X1 U619 ( .A(G82), .ZN(G220) );
  NAND2_X1 U620 ( .A1(G7), .A2(G661), .ZN(n562) );
  XNOR2_X1 U621 ( .A(n562), .B(KEYINPUT10), .ZN(G223) );
  XNOR2_X1 U622 ( .A(G223), .B(KEYINPUT69), .ZN(n830) );
  NAND2_X1 U623 ( .A1(n830), .A2(G567), .ZN(n563) );
  XOR2_X1 U624 ( .A(KEYINPUT11), .B(n563), .Z(G234) );
  INV_X1 U625 ( .A(G860), .ZN(n603) );
  NAND2_X1 U626 ( .A1(n649), .A2(G81), .ZN(n564) );
  XNOR2_X1 U627 ( .A(n564), .B(KEYINPUT12), .ZN(n566) );
  NAND2_X1 U628 ( .A1(G68), .A2(n650), .ZN(n565) );
  NAND2_X1 U629 ( .A1(n566), .A2(n565), .ZN(n568) );
  XOR2_X1 U630 ( .A(KEYINPUT70), .B(KEYINPUT13), .Z(n567) );
  XNOR2_X1 U631 ( .A(n568), .B(n567), .ZN(n571) );
  NAND2_X1 U632 ( .A1(n653), .A2(G56), .ZN(n569) );
  XOR2_X1 U633 ( .A(KEYINPUT14), .B(n569), .Z(n570) );
  NOR2_X1 U634 ( .A1(n571), .A2(n570), .ZN(n573) );
  NAND2_X1 U635 ( .A1(n654), .A2(G43), .ZN(n572) );
  NAND2_X1 U636 ( .A1(n573), .A2(n572), .ZN(n994) );
  NOR2_X1 U637 ( .A1(n603), .A2(n994), .ZN(n574) );
  XNOR2_X1 U638 ( .A(n574), .B(KEYINPUT71), .ZN(G153) );
  NAND2_X1 U639 ( .A1(G64), .A2(n653), .ZN(n576) );
  NAND2_X1 U640 ( .A1(G52), .A2(n654), .ZN(n575) );
  NAND2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n581) );
  NAND2_X1 U642 ( .A1(G90), .A2(n649), .ZN(n578) );
  NAND2_X1 U643 ( .A1(G77), .A2(n650), .ZN(n577) );
  NAND2_X1 U644 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U645 ( .A(KEYINPUT9), .B(n579), .Z(n580) );
  NOR2_X1 U646 ( .A1(n581), .A2(n580), .ZN(G171) );
  INV_X1 U647 ( .A(G171), .ZN(G301) );
  NAND2_X1 U648 ( .A1(G66), .A2(n653), .ZN(n582) );
  XNOR2_X1 U649 ( .A(n582), .B(KEYINPUT72), .ZN(n589) );
  NAND2_X1 U650 ( .A1(G92), .A2(n649), .ZN(n584) );
  NAND2_X1 U651 ( .A1(G79), .A2(n650), .ZN(n583) );
  NAND2_X1 U652 ( .A1(n584), .A2(n583), .ZN(n587) );
  NAND2_X1 U653 ( .A1(G54), .A2(n654), .ZN(n585) );
  XNOR2_X1 U654 ( .A(KEYINPUT73), .B(n585), .ZN(n586) );
  NOR2_X1 U655 ( .A1(n587), .A2(n586), .ZN(n588) );
  NAND2_X1 U656 ( .A1(n589), .A2(n588), .ZN(n591) );
  XOR2_X1 U657 ( .A(KEYINPUT74), .B(KEYINPUT15), .Z(n590) );
  XOR2_X1 U658 ( .A(n591), .B(n590), .Z(n904) );
  INV_X1 U659 ( .A(n904), .ZN(n995) );
  NOR2_X1 U660 ( .A1(n995), .A2(G868), .ZN(n593) );
  INV_X1 U661 ( .A(G868), .ZN(n607) );
  NOR2_X1 U662 ( .A1(n607), .A2(G301), .ZN(n592) );
  NOR2_X1 U663 ( .A1(n593), .A2(n592), .ZN(G284) );
  NAND2_X1 U664 ( .A1(G65), .A2(n653), .ZN(n595) );
  NAND2_X1 U665 ( .A1(G53), .A2(n654), .ZN(n594) );
  NAND2_X1 U666 ( .A1(n595), .A2(n594), .ZN(n599) );
  NAND2_X1 U667 ( .A1(G91), .A2(n649), .ZN(n597) );
  NAND2_X1 U668 ( .A1(G78), .A2(n650), .ZN(n596) );
  NAND2_X1 U669 ( .A1(n597), .A2(n596), .ZN(n598) );
  NOR2_X1 U670 ( .A1(n599), .A2(n598), .ZN(n713) );
  INV_X1 U671 ( .A(n713), .ZN(G299) );
  NOR2_X1 U672 ( .A1(G286), .A2(n607), .ZN(n600) );
  XNOR2_X1 U673 ( .A(n600), .B(KEYINPUT78), .ZN(n602) );
  NOR2_X1 U674 ( .A1(G299), .A2(G868), .ZN(n601) );
  NOR2_X1 U675 ( .A1(n602), .A2(n601), .ZN(G297) );
  NAND2_X1 U676 ( .A1(n603), .A2(G559), .ZN(n604) );
  NAND2_X1 U677 ( .A1(n604), .A2(n904), .ZN(n605) );
  XNOR2_X1 U678 ( .A(n605), .B(KEYINPUT16), .ZN(n606) );
  XOR2_X1 U679 ( .A(KEYINPUT79), .B(n606), .Z(G148) );
  NOR2_X1 U680 ( .A1(n995), .A2(n607), .ZN(n608) );
  XOR2_X1 U681 ( .A(KEYINPUT80), .B(n608), .Z(n609) );
  NOR2_X1 U682 ( .A1(G559), .A2(n609), .ZN(n611) );
  NOR2_X1 U683 ( .A1(G868), .A2(n994), .ZN(n610) );
  NOR2_X1 U684 ( .A1(n611), .A2(n610), .ZN(G282) );
  NAND2_X1 U685 ( .A1(G135), .A2(n1015), .ZN(n613) );
  NAND2_X1 U686 ( .A1(G111), .A2(n1012), .ZN(n612) );
  NAND2_X1 U687 ( .A1(n613), .A2(n612), .ZN(n620) );
  NAND2_X1 U688 ( .A1(G99), .A2(n519), .ZN(n614) );
  XNOR2_X1 U689 ( .A(n614), .B(KEYINPUT82), .ZN(n618) );
  XOR2_X1 U690 ( .A(KEYINPUT81), .B(KEYINPUT18), .Z(n616) );
  NAND2_X1 U691 ( .A1(G123), .A2(n1011), .ZN(n615) );
  XNOR2_X1 U692 ( .A(n616), .B(n615), .ZN(n617) );
  NAND2_X1 U693 ( .A1(n618), .A2(n617), .ZN(n619) );
  NOR2_X1 U694 ( .A1(n620), .A2(n619), .ZN(n1025) );
  XNOR2_X1 U695 ( .A(n1025), .B(G2096), .ZN(n621) );
  INV_X1 U696 ( .A(G2100), .ZN(n988) );
  NAND2_X1 U697 ( .A1(n621), .A2(n988), .ZN(G156) );
  NAND2_X1 U698 ( .A1(G88), .A2(n649), .ZN(n623) );
  NAND2_X1 U699 ( .A1(G75), .A2(n650), .ZN(n622) );
  NAND2_X1 U700 ( .A1(n623), .A2(n622), .ZN(n628) );
  NAND2_X1 U701 ( .A1(G62), .A2(n653), .ZN(n625) );
  NAND2_X1 U702 ( .A1(G50), .A2(n654), .ZN(n624) );
  NAND2_X1 U703 ( .A1(n625), .A2(n624), .ZN(n626) );
  XOR2_X1 U704 ( .A(KEYINPUT85), .B(n626), .Z(n627) );
  NOR2_X1 U705 ( .A1(n628), .A2(n627), .ZN(G166) );
  NAND2_X1 U706 ( .A1(G74), .A2(G651), .ZN(n633) );
  NAND2_X1 U707 ( .A1(G49), .A2(n654), .ZN(n630) );
  NAND2_X1 U708 ( .A1(G87), .A2(n530), .ZN(n629) );
  NAND2_X1 U709 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U710 ( .A1(n653), .A2(n631), .ZN(n632) );
  NAND2_X1 U711 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U712 ( .A(n634), .B(KEYINPUT84), .ZN(G288) );
  NAND2_X1 U713 ( .A1(G60), .A2(n653), .ZN(n636) );
  NAND2_X1 U714 ( .A1(G47), .A2(n654), .ZN(n635) );
  NAND2_X1 U715 ( .A1(n636), .A2(n635), .ZN(n639) );
  NAND2_X1 U716 ( .A1(G85), .A2(n649), .ZN(n637) );
  XOR2_X1 U717 ( .A(KEYINPUT68), .B(n637), .Z(n638) );
  NOR2_X1 U718 ( .A1(n639), .A2(n638), .ZN(n641) );
  NAND2_X1 U719 ( .A1(n650), .A2(G72), .ZN(n640) );
  NAND2_X1 U720 ( .A1(n641), .A2(n640), .ZN(G290) );
  NAND2_X1 U721 ( .A1(G86), .A2(n649), .ZN(n643) );
  NAND2_X1 U722 ( .A1(G61), .A2(n653), .ZN(n642) );
  NAND2_X1 U723 ( .A1(n643), .A2(n642), .ZN(n646) );
  NAND2_X1 U724 ( .A1(n650), .A2(G73), .ZN(n644) );
  XOR2_X1 U725 ( .A(KEYINPUT2), .B(n644), .Z(n645) );
  NOR2_X1 U726 ( .A1(n646), .A2(n645), .ZN(n648) );
  NAND2_X1 U727 ( .A1(n654), .A2(G48), .ZN(n647) );
  NAND2_X1 U728 ( .A1(n648), .A2(n647), .ZN(G305) );
  XNOR2_X1 U729 ( .A(G166), .B(G288), .ZN(n660) );
  NAND2_X1 U730 ( .A1(G93), .A2(n649), .ZN(n652) );
  NAND2_X1 U731 ( .A1(G80), .A2(n650), .ZN(n651) );
  NAND2_X1 U732 ( .A1(n652), .A2(n651), .ZN(n658) );
  NAND2_X1 U733 ( .A1(G67), .A2(n653), .ZN(n656) );
  NAND2_X1 U734 ( .A1(G55), .A2(n654), .ZN(n655) );
  NAND2_X1 U735 ( .A1(n656), .A2(n655), .ZN(n657) );
  NOR2_X1 U736 ( .A1(n658), .A2(n657), .ZN(n659) );
  XOR2_X1 U737 ( .A(KEYINPUT83), .B(n659), .Z(n958) );
  XNOR2_X1 U738 ( .A(n660), .B(n958), .ZN(n661) );
  XOR2_X1 U739 ( .A(n661), .B(KEYINPUT19), .Z(n663) );
  XOR2_X1 U740 ( .A(G299), .B(KEYINPUT86), .Z(n662) );
  XNOR2_X1 U741 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U742 ( .A(n664), .B(G290), .ZN(n665) );
  XNOR2_X1 U743 ( .A(n665), .B(G305), .ZN(n993) );
  NAND2_X1 U744 ( .A1(n904), .A2(G559), .ZN(n666) );
  XNOR2_X1 U745 ( .A(n994), .B(n666), .ZN(n957) );
  XOR2_X1 U746 ( .A(n993), .B(n957), .Z(n667) );
  NAND2_X1 U747 ( .A1(n667), .A2(G868), .ZN(n668) );
  XNOR2_X1 U748 ( .A(n668), .B(KEYINPUT87), .ZN(n670) );
  NOR2_X1 U749 ( .A1(n958), .A2(G868), .ZN(n669) );
  NOR2_X1 U750 ( .A1(n670), .A2(n669), .ZN(n671) );
  XOR2_X1 U751 ( .A(KEYINPUT88), .B(n671), .Z(G295) );
  NAND2_X1 U752 ( .A1(G2078), .A2(G2084), .ZN(n672) );
  XOR2_X1 U753 ( .A(KEYINPUT20), .B(n672), .Z(n673) );
  NAND2_X1 U754 ( .A1(G2090), .A2(n673), .ZN(n674) );
  XNOR2_X1 U755 ( .A(KEYINPUT21), .B(n674), .ZN(n675) );
  NAND2_X1 U756 ( .A1(n675), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U757 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U758 ( .A1(G220), .A2(G219), .ZN(n676) );
  XNOR2_X1 U759 ( .A(KEYINPUT22), .B(n676), .ZN(n677) );
  NAND2_X1 U760 ( .A1(n677), .A2(G96), .ZN(n678) );
  NOR2_X1 U761 ( .A1(n678), .A2(G218), .ZN(n679) );
  XNOR2_X1 U762 ( .A(n679), .B(KEYINPUT89), .ZN(n955) );
  NAND2_X1 U763 ( .A1(n955), .A2(G2106), .ZN(n683) );
  NAND2_X1 U764 ( .A1(G120), .A2(G69), .ZN(n680) );
  NOR2_X1 U765 ( .A1(G237), .A2(n680), .ZN(n681) );
  NAND2_X1 U766 ( .A1(G108), .A2(n681), .ZN(n956) );
  NAND2_X1 U767 ( .A1(n956), .A2(G567), .ZN(n682) );
  NAND2_X1 U768 ( .A1(n683), .A2(n682), .ZN(n1035) );
  NAND2_X1 U769 ( .A1(G483), .A2(G661), .ZN(n684) );
  NOR2_X1 U770 ( .A1(n1035), .A2(n684), .ZN(n833) );
  NAND2_X1 U771 ( .A1(n833), .A2(G36), .ZN(G176) );
  XOR2_X1 U772 ( .A(G166), .B(KEYINPUT90), .Z(G303) );
  INV_X1 U773 ( .A(G40), .ZN(n686) );
  NOR2_X1 U774 ( .A1(G164), .A2(G1384), .ZN(n766) );
  INV_X1 U775 ( .A(n766), .ZN(n685) );
  NOR2_X1 U776 ( .A1(n686), .A2(n685), .ZN(n687) );
  INV_X1 U777 ( .A(KEYINPUT26), .ZN(n688) );
  XNOR2_X1 U778 ( .A(n689), .B(n688), .ZN(n693) );
  INV_X1 U779 ( .A(G1341), .ZN(n690) );
  NOR2_X1 U780 ( .A1(n690), .A2(n695), .ZN(n691) );
  NOR2_X1 U781 ( .A1(n691), .A2(n994), .ZN(n692) );
  NAND2_X1 U782 ( .A1(n693), .A2(n692), .ZN(n705) );
  XNOR2_X1 U783 ( .A(KEYINPUT94), .B(n694), .ZN(n703) );
  NOR2_X1 U784 ( .A1(n695), .A2(G1348), .ZN(n697) );
  NOR2_X1 U785 ( .A1(G2067), .A2(n741), .ZN(n696) );
  NOR2_X1 U786 ( .A1(n697), .A2(n696), .ZN(n701) );
  NAND2_X1 U787 ( .A1(n695), .A2(G2072), .ZN(n698) );
  XNOR2_X1 U788 ( .A(n698), .B(KEYINPUT27), .ZN(n700) );
  INV_X1 U789 ( .A(G1956), .ZN(n975) );
  NOR2_X1 U790 ( .A1(n975), .A2(n695), .ZN(n699) );
  NOR2_X1 U791 ( .A1(n700), .A2(n699), .ZN(n712) );
  NAND2_X1 U792 ( .A1(n713), .A2(n712), .ZN(n704) );
  NAND2_X1 U793 ( .A1(n701), .A2(n704), .ZN(n702) );
  NOR2_X1 U794 ( .A1(n703), .A2(n702), .ZN(n709) );
  INV_X1 U795 ( .A(n704), .ZN(n707) );
  NAND2_X1 U796 ( .A1(n995), .A2(n705), .ZN(n706) );
  NOR2_X1 U797 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U798 ( .A(n711), .B(n710), .ZN(n716) );
  OR2_X1 U799 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U800 ( .A(KEYINPUT28), .B(n714), .ZN(n715) );
  NAND2_X1 U801 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U802 ( .A(n717), .B(KEYINPUT29), .ZN(n721) );
  XOR2_X1 U803 ( .A(G2078), .B(KEYINPUT25), .Z(n877) );
  NOR2_X1 U804 ( .A1(n877), .A2(n741), .ZN(n719) );
  NOR2_X1 U805 ( .A1(n695), .A2(G1961), .ZN(n718) );
  NOR2_X1 U806 ( .A1(n719), .A2(n718), .ZN(n729) );
  NOR2_X1 U807 ( .A1(G301), .A2(n729), .ZN(n720) );
  NOR2_X1 U808 ( .A1(n721), .A2(n720), .ZN(n738) );
  NOR2_X1 U809 ( .A1(n804), .A2(G1966), .ZN(n722) );
  XNOR2_X1 U810 ( .A(n722), .B(KEYINPUT93), .ZN(n750) );
  INV_X1 U811 ( .A(G8), .ZN(n723) );
  NOR2_X1 U812 ( .A1(G2084), .A2(n741), .ZN(n749) );
  NOR2_X1 U813 ( .A1(n723), .A2(n749), .ZN(n724) );
  AND2_X1 U814 ( .A1(n750), .A2(n724), .ZN(n725) );
  XNOR2_X1 U815 ( .A(n725), .B(n520), .ZN(n727) );
  INV_X1 U816 ( .A(G168), .ZN(n726) );
  XNOR2_X1 U817 ( .A(n728), .B(KEYINPUT97), .ZN(n731) );
  NAND2_X1 U818 ( .A1(n729), .A2(G301), .ZN(n730) );
  INV_X1 U819 ( .A(KEYINPUT31), .ZN(n732) );
  NAND2_X1 U820 ( .A1(n733), .A2(n732), .ZN(n736) );
  INV_X1 U821 ( .A(n733), .ZN(n734) );
  NAND2_X1 U822 ( .A1(n734), .A2(KEYINPUT31), .ZN(n735) );
  NAND2_X1 U823 ( .A1(n736), .A2(n735), .ZN(n737) );
  NOR2_X1 U824 ( .A1(n738), .A2(n737), .ZN(n740) );
  XNOR2_X1 U825 ( .A(n740), .B(n739), .ZN(n751) );
  NAND2_X1 U826 ( .A1(n751), .A2(G286), .ZN(n746) );
  NOR2_X1 U827 ( .A1(G1971), .A2(n804), .ZN(n743) );
  NOR2_X1 U828 ( .A1(G2090), .A2(n741), .ZN(n742) );
  NOR2_X1 U829 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U830 ( .A1(n744), .A2(G303), .ZN(n745) );
  NAND2_X1 U831 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U832 ( .A1(n747), .A2(G8), .ZN(n748) );
  NAND2_X1 U833 ( .A1(G8), .A2(n749), .ZN(n753) );
  AND2_X1 U834 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U835 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U836 ( .A1(n755), .A2(n754), .ZN(n800) );
  NOR2_X1 U837 ( .A1(G1976), .A2(G288), .ZN(n908) );
  NOR2_X1 U838 ( .A1(G303), .A2(G1971), .ZN(n756) );
  NOR2_X1 U839 ( .A1(n908), .A2(n756), .ZN(n757) );
  XOR2_X1 U840 ( .A(KEYINPUT99), .B(n757), .Z(n759) );
  INV_X1 U841 ( .A(KEYINPUT33), .ZN(n758) );
  AND2_X1 U842 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U843 ( .A1(n800), .A2(n760), .ZN(n763) );
  NAND2_X1 U844 ( .A1(G1976), .A2(G288), .ZN(n902) );
  INV_X1 U845 ( .A(n902), .ZN(n761) );
  OR2_X1 U846 ( .A1(KEYINPUT33), .A2(n523), .ZN(n762) );
  NAND2_X1 U847 ( .A1(n763), .A2(n762), .ZN(n764) );
  XOR2_X1 U848 ( .A(G1981), .B(G305), .Z(n895) );
  NAND2_X1 U849 ( .A1(G40), .A2(G160), .ZN(n765) );
  NOR2_X1 U850 ( .A1(n766), .A2(n765), .ZN(n825) );
  NAND2_X1 U851 ( .A1(G140), .A2(n1015), .ZN(n768) );
  NAND2_X1 U852 ( .A1(G104), .A2(n519), .ZN(n767) );
  NAND2_X1 U853 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U854 ( .A(KEYINPUT34), .B(n769), .ZN(n775) );
  NAND2_X1 U855 ( .A1(n1011), .A2(G128), .ZN(n770) );
  XOR2_X1 U856 ( .A(KEYINPUT91), .B(n770), .Z(n772) );
  NAND2_X1 U857 ( .A1(G116), .A2(n1012), .ZN(n771) );
  NAND2_X1 U858 ( .A1(n772), .A2(n771), .ZN(n773) );
  XOR2_X1 U859 ( .A(KEYINPUT35), .B(n773), .Z(n774) );
  NOR2_X1 U860 ( .A1(n775), .A2(n774), .ZN(n776) );
  XOR2_X1 U861 ( .A(KEYINPUT36), .B(n776), .Z(n1001) );
  XOR2_X1 U862 ( .A(G2067), .B(KEYINPUT37), .Z(n821) );
  AND2_X1 U863 ( .A1(n1001), .A2(n821), .ZN(n856) );
  NAND2_X1 U864 ( .A1(n825), .A2(n856), .ZN(n819) );
  NAND2_X1 U865 ( .A1(G131), .A2(n1015), .ZN(n778) );
  NAND2_X1 U866 ( .A1(G107), .A2(n1012), .ZN(n777) );
  NAND2_X1 U867 ( .A1(n778), .A2(n777), .ZN(n782) );
  NAND2_X1 U868 ( .A1(G95), .A2(n519), .ZN(n780) );
  NAND2_X1 U869 ( .A1(G119), .A2(n1011), .ZN(n779) );
  NAND2_X1 U870 ( .A1(n780), .A2(n779), .ZN(n781) );
  OR2_X1 U871 ( .A1(n782), .A2(n781), .ZN(n1022) );
  NAND2_X1 U872 ( .A1(G1991), .A2(n1022), .ZN(n783) );
  XOR2_X1 U873 ( .A(KEYINPUT92), .B(n783), .Z(n792) );
  NAND2_X1 U874 ( .A1(G141), .A2(n1015), .ZN(n785) );
  NAND2_X1 U875 ( .A1(G129), .A2(n1011), .ZN(n784) );
  NAND2_X1 U876 ( .A1(n785), .A2(n784), .ZN(n788) );
  NAND2_X1 U877 ( .A1(n519), .A2(G105), .ZN(n786) );
  XOR2_X1 U878 ( .A(KEYINPUT38), .B(n786), .Z(n787) );
  NOR2_X1 U879 ( .A1(n788), .A2(n787), .ZN(n790) );
  NAND2_X1 U880 ( .A1(G117), .A2(n1012), .ZN(n789) );
  NAND2_X1 U881 ( .A1(n790), .A2(n789), .ZN(n1000) );
  AND2_X1 U882 ( .A1(n1000), .A2(G1996), .ZN(n791) );
  NOR2_X1 U883 ( .A1(n792), .A2(n791), .ZN(n854) );
  INV_X1 U884 ( .A(n854), .ZN(n793) );
  NAND2_X1 U885 ( .A1(n793), .A2(n825), .ZN(n813) );
  NAND2_X1 U886 ( .A1(n819), .A2(n813), .ZN(n808) );
  INV_X1 U887 ( .A(n808), .ZN(n794) );
  NAND2_X1 U888 ( .A1(n908), .A2(KEYINPUT33), .ZN(n795) );
  NOR2_X1 U889 ( .A1(n804), .A2(n795), .ZN(n796) );
  NAND2_X1 U890 ( .A1(n524), .A2(n797), .ZN(n810) );
  NOR2_X1 U891 ( .A1(G2090), .A2(G303), .ZN(n798) );
  NAND2_X1 U892 ( .A1(G8), .A2(n798), .ZN(n799) );
  NAND2_X1 U893 ( .A1(n800), .A2(n799), .ZN(n801) );
  AND2_X1 U894 ( .A1(n804), .A2(n801), .ZN(n806) );
  NOR2_X1 U895 ( .A1(G1981), .A2(G305), .ZN(n802) );
  XOR2_X1 U896 ( .A(n802), .B(KEYINPUT24), .Z(n803) );
  NOR2_X1 U897 ( .A1(n804), .A2(n803), .ZN(n805) );
  NOR2_X1 U898 ( .A1(n806), .A2(n805), .ZN(n807) );
  OR2_X1 U899 ( .A1(n808), .A2(n807), .ZN(n809) );
  NAND2_X1 U900 ( .A1(n810), .A2(n809), .ZN(n812) );
  XNOR2_X1 U901 ( .A(G1986), .B(G290), .ZN(n901) );
  NAND2_X1 U902 ( .A1(n901), .A2(n825), .ZN(n811) );
  NAND2_X1 U903 ( .A1(n812), .A2(n811), .ZN(n828) );
  NOR2_X1 U904 ( .A1(G1996), .A2(n1000), .ZN(n860) );
  INV_X1 U905 ( .A(n813), .ZN(n816) );
  NOR2_X1 U906 ( .A1(G1991), .A2(n1022), .ZN(n852) );
  NOR2_X1 U907 ( .A1(G1986), .A2(G290), .ZN(n814) );
  NOR2_X1 U908 ( .A1(n852), .A2(n814), .ZN(n815) );
  NOR2_X1 U909 ( .A1(n816), .A2(n815), .ZN(n817) );
  NOR2_X1 U910 ( .A1(n860), .A2(n817), .ZN(n818) );
  XNOR2_X1 U911 ( .A(n818), .B(KEYINPUT39), .ZN(n820) );
  NAND2_X1 U912 ( .A1(n820), .A2(n819), .ZN(n823) );
  NOR2_X1 U913 ( .A1(n1001), .A2(n821), .ZN(n822) );
  XNOR2_X1 U914 ( .A(KEYINPUT101), .B(n822), .ZN(n863) );
  NAND2_X1 U915 ( .A1(n823), .A2(n863), .ZN(n824) );
  XNOR2_X1 U916 ( .A(KEYINPUT102), .B(n824), .ZN(n826) );
  NAND2_X1 U917 ( .A1(n826), .A2(n825), .ZN(n827) );
  NAND2_X1 U918 ( .A1(n828), .A2(n827), .ZN(n829) );
  XNOR2_X1 U919 ( .A(n829), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U920 ( .A1(G2106), .A2(n830), .ZN(G217) );
  AND2_X1 U921 ( .A1(G15), .A2(G2), .ZN(n831) );
  NAND2_X1 U922 ( .A1(G661), .A2(n831), .ZN(G259) );
  NAND2_X1 U923 ( .A1(G3), .A2(G1), .ZN(n832) );
  NAND2_X1 U924 ( .A1(n833), .A2(n832), .ZN(G188) );
  XOR2_X1 U925 ( .A(G69), .B(KEYINPUT104), .Z(G235) );
  NAND2_X1 U927 ( .A1(n1012), .A2(G112), .ZN(n840) );
  NAND2_X1 U928 ( .A1(G136), .A2(n1015), .ZN(n835) );
  NAND2_X1 U929 ( .A1(G100), .A2(n519), .ZN(n834) );
  NAND2_X1 U930 ( .A1(n835), .A2(n834), .ZN(n838) );
  NAND2_X1 U931 ( .A1(n1011), .A2(G124), .ZN(n836) );
  XOR2_X1 U932 ( .A(KEYINPUT44), .B(n836), .Z(n837) );
  NOR2_X1 U933 ( .A1(n838), .A2(n837), .ZN(n839) );
  NAND2_X1 U934 ( .A1(n840), .A2(n839), .ZN(n841) );
  XNOR2_X1 U935 ( .A(n841), .B(KEYINPUT109), .ZN(G162) );
  NAND2_X1 U936 ( .A1(G139), .A2(n1015), .ZN(n843) );
  NAND2_X1 U937 ( .A1(G103), .A2(n519), .ZN(n842) );
  NAND2_X1 U938 ( .A1(n843), .A2(n842), .ZN(n848) );
  NAND2_X1 U939 ( .A1(n1011), .A2(G127), .ZN(n845) );
  NAND2_X1 U940 ( .A1(G115), .A2(n1012), .ZN(n844) );
  NAND2_X1 U941 ( .A1(n845), .A2(n844), .ZN(n846) );
  XOR2_X1 U942 ( .A(KEYINPUT47), .B(n846), .Z(n847) );
  NOR2_X1 U943 ( .A1(n848), .A2(n847), .ZN(n1008) );
  XOR2_X1 U944 ( .A(G2072), .B(n1008), .Z(n850) );
  XOR2_X1 U945 ( .A(G164), .B(G2078), .Z(n849) );
  NOR2_X1 U946 ( .A1(n850), .A2(n849), .ZN(n851) );
  XOR2_X1 U947 ( .A(KEYINPUT50), .B(n851), .Z(n869) );
  XNOR2_X1 U948 ( .A(G2084), .B(G160), .ZN(n858) );
  NOR2_X1 U949 ( .A1(n852), .A2(n1025), .ZN(n853) );
  NAND2_X1 U950 ( .A1(n854), .A2(n853), .ZN(n855) );
  NOR2_X1 U951 ( .A1(n856), .A2(n855), .ZN(n857) );
  NAND2_X1 U952 ( .A1(n858), .A2(n857), .ZN(n866) );
  XOR2_X1 U953 ( .A(G2090), .B(G162), .Z(n859) );
  NOR2_X1 U954 ( .A1(n860), .A2(n859), .ZN(n861) );
  XNOR2_X1 U955 ( .A(KEYINPUT51), .B(n861), .ZN(n862) );
  XNOR2_X1 U956 ( .A(n862), .B(KEYINPUT113), .ZN(n864) );
  NAND2_X1 U957 ( .A1(n864), .A2(n863), .ZN(n865) );
  NOR2_X1 U958 ( .A1(n866), .A2(n865), .ZN(n867) );
  XOR2_X1 U959 ( .A(KEYINPUT114), .B(n867), .Z(n868) );
  NOR2_X1 U960 ( .A1(n869), .A2(n868), .ZN(n870) );
  XNOR2_X1 U961 ( .A(n870), .B(KEYINPUT52), .ZN(n871) );
  XNOR2_X1 U962 ( .A(KEYINPUT55), .B(KEYINPUT115), .ZN(n890) );
  NAND2_X1 U963 ( .A1(n871), .A2(n890), .ZN(n872) );
  XNOR2_X1 U964 ( .A(KEYINPUT116), .B(n872), .ZN(n873) );
  NAND2_X1 U965 ( .A1(n873), .A2(G29), .ZN(n953) );
  XOR2_X1 U966 ( .A(G1991), .B(G25), .Z(n874) );
  NAND2_X1 U967 ( .A1(n874), .A2(G28), .ZN(n883) );
  XNOR2_X1 U968 ( .A(G2067), .B(G26), .ZN(n876) );
  XNOR2_X1 U969 ( .A(G33), .B(G2072), .ZN(n875) );
  NOR2_X1 U970 ( .A1(n876), .A2(n875), .ZN(n881) );
  XNOR2_X1 U971 ( .A(G1996), .B(G32), .ZN(n879) );
  XNOR2_X1 U972 ( .A(G27), .B(n877), .ZN(n878) );
  NOR2_X1 U973 ( .A1(n879), .A2(n878), .ZN(n880) );
  NAND2_X1 U974 ( .A1(n881), .A2(n880), .ZN(n882) );
  NOR2_X1 U975 ( .A1(n883), .A2(n882), .ZN(n884) );
  XOR2_X1 U976 ( .A(KEYINPUT53), .B(n884), .Z(n887) );
  XOR2_X1 U977 ( .A(KEYINPUT54), .B(G34), .Z(n885) );
  XNOR2_X1 U978 ( .A(G2084), .B(n885), .ZN(n886) );
  NAND2_X1 U979 ( .A1(n887), .A2(n886), .ZN(n889) );
  XNOR2_X1 U980 ( .A(G35), .B(G2090), .ZN(n888) );
  NOR2_X1 U981 ( .A1(n889), .A2(n888), .ZN(n891) );
  XNOR2_X1 U982 ( .A(n891), .B(n890), .ZN(n892) );
  NOR2_X1 U983 ( .A1(G29), .A2(n892), .ZN(n893) );
  XNOR2_X1 U984 ( .A(KEYINPUT117), .B(n893), .ZN(n894) );
  NAND2_X1 U985 ( .A1(n894), .A2(G11), .ZN(n951) );
  INV_X1 U986 ( .A(G16), .ZN(n946) );
  XOR2_X1 U987 ( .A(n946), .B(KEYINPUT56), .Z(n919) );
  XNOR2_X1 U988 ( .A(G1966), .B(G168), .ZN(n896) );
  NAND2_X1 U989 ( .A1(n896), .A2(n895), .ZN(n897) );
  XNOR2_X1 U990 ( .A(n897), .B(KEYINPUT57), .ZN(n917) );
  XOR2_X1 U991 ( .A(G299), .B(G1956), .Z(n899) );
  XOR2_X1 U992 ( .A(G301), .B(G1961), .Z(n898) );
  NAND2_X1 U993 ( .A1(n899), .A2(n898), .ZN(n900) );
  NOR2_X1 U994 ( .A1(n901), .A2(n900), .ZN(n903) );
  NAND2_X1 U995 ( .A1(n903), .A2(n902), .ZN(n907) );
  XOR2_X1 U996 ( .A(n904), .B(G1348), .Z(n905) );
  XNOR2_X1 U997 ( .A(KEYINPUT118), .B(n905), .ZN(n906) );
  NOR2_X1 U998 ( .A1(n907), .A2(n906), .ZN(n912) );
  XOR2_X1 U999 ( .A(n908), .B(KEYINPUT119), .Z(n910) );
  XNOR2_X1 U1000 ( .A(G303), .B(G1971), .ZN(n909) );
  NOR2_X1 U1001 ( .A1(n910), .A2(n909), .ZN(n911) );
  NAND2_X1 U1002 ( .A1(n912), .A2(n911), .ZN(n913) );
  XNOR2_X1 U1003 ( .A(KEYINPUT120), .B(n913), .ZN(n915) );
  XNOR2_X1 U1004 ( .A(G1341), .B(n994), .ZN(n914) );
  NOR2_X1 U1005 ( .A1(n915), .A2(n914), .ZN(n916) );
  NAND2_X1 U1006 ( .A1(n917), .A2(n916), .ZN(n918) );
  NAND2_X1 U1007 ( .A1(n919), .A2(n918), .ZN(n948) );
  XNOR2_X1 U1008 ( .A(G1966), .B(G21), .ZN(n931) );
  XNOR2_X1 U1009 ( .A(KEYINPUT121), .B(KEYINPUT122), .ZN(n920) );
  XNOR2_X1 U1010 ( .A(n920), .B(KEYINPUT60), .ZN(n929) );
  XOR2_X1 U1011 ( .A(G20), .B(G1956), .Z(n924) );
  XNOR2_X1 U1012 ( .A(G1341), .B(G19), .ZN(n922) );
  XNOR2_X1 U1013 ( .A(G1981), .B(G6), .ZN(n921) );
  NOR2_X1 U1014 ( .A1(n922), .A2(n921), .ZN(n923) );
  NAND2_X1 U1015 ( .A1(n924), .A2(n923), .ZN(n927) );
  XOR2_X1 U1016 ( .A(KEYINPUT59), .B(G1348), .Z(n925) );
  XNOR2_X1 U1017 ( .A(G4), .B(n925), .ZN(n926) );
  NOR2_X1 U1018 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1019 ( .A(n929), .B(n928), .ZN(n930) );
  NOR2_X1 U1020 ( .A1(n931), .A2(n930), .ZN(n932) );
  XOR2_X1 U1021 ( .A(KEYINPUT123), .B(n932), .Z(n941) );
  XOR2_X1 U1022 ( .A(G1976), .B(KEYINPUT124), .Z(n933) );
  XNOR2_X1 U1023 ( .A(G23), .B(n933), .ZN(n937) );
  XNOR2_X1 U1024 ( .A(G1986), .B(G24), .ZN(n935) );
  XNOR2_X1 U1025 ( .A(G1971), .B(G22), .ZN(n934) );
  NOR2_X1 U1026 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1027 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1028 ( .A(n938), .B(KEYINPUT125), .ZN(n939) );
  XNOR2_X1 U1029 ( .A(KEYINPUT58), .B(n939), .ZN(n940) );
  NAND2_X1 U1030 ( .A1(n941), .A2(n940), .ZN(n943) );
  XNOR2_X1 U1031 ( .A(G5), .B(G1961), .ZN(n942) );
  NOR2_X1 U1032 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1033 ( .A(KEYINPUT61), .B(n944), .ZN(n945) );
  NAND2_X1 U1034 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1035 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1036 ( .A(n949), .B(KEYINPUT126), .ZN(n950) );
  NOR2_X1 U1037 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1038 ( .A1(n953), .A2(n952), .ZN(n954) );
  XOR2_X1 U1039 ( .A(KEYINPUT62), .B(n954), .Z(G311) );
  XNOR2_X1 U1040 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1041 ( .A(G120), .ZN(G236) );
  INV_X1 U1042 ( .A(G96), .ZN(G221) );
  NOR2_X1 U1043 ( .A1(n956), .A2(n955), .ZN(G325) );
  INV_X1 U1044 ( .A(G325), .ZN(G261) );
  NOR2_X1 U1045 ( .A1(n957), .A2(G860), .ZN(n959) );
  XNOR2_X1 U1046 ( .A(n959), .B(n958), .ZN(G145) );
  XNOR2_X1 U1047 ( .A(G1341), .B(G2454), .ZN(n960) );
  XNOR2_X1 U1048 ( .A(n960), .B(G2430), .ZN(n961) );
  XNOR2_X1 U1049 ( .A(n961), .B(G1348), .ZN(n967) );
  XOR2_X1 U1050 ( .A(G2443), .B(G2427), .Z(n963) );
  XNOR2_X1 U1051 ( .A(G2438), .B(G2446), .ZN(n962) );
  XNOR2_X1 U1052 ( .A(n963), .B(n962), .ZN(n965) );
  XOR2_X1 U1053 ( .A(G2451), .B(G2435), .Z(n964) );
  XNOR2_X1 U1054 ( .A(n965), .B(n964), .ZN(n966) );
  XNOR2_X1 U1055 ( .A(n967), .B(n966), .ZN(n968) );
  NAND2_X1 U1056 ( .A1(n968), .A2(G14), .ZN(n969) );
  XNOR2_X1 U1057 ( .A(KEYINPUT103), .B(n969), .ZN(G401) );
  XOR2_X1 U1058 ( .A(KEYINPUT108), .B(G2474), .Z(n971) );
  XNOR2_X1 U1059 ( .A(G1991), .B(G1986), .ZN(n970) );
  XNOR2_X1 U1060 ( .A(n971), .B(n970), .ZN(n972) );
  XOR2_X1 U1061 ( .A(n972), .B(G1976), .Z(n974) );
  XNOR2_X1 U1062 ( .A(G1996), .B(G1961), .ZN(n973) );
  XNOR2_X1 U1063 ( .A(n974), .B(n973), .ZN(n979) );
  XOR2_X1 U1064 ( .A(KEYINPUT107), .B(KEYINPUT41), .Z(n977) );
  XOR2_X1 U1065 ( .A(n975), .B(G1971), .Z(n976) );
  XNOR2_X1 U1066 ( .A(n977), .B(n976), .ZN(n978) );
  XOR2_X1 U1067 ( .A(n979), .B(n978), .Z(n981) );
  XNOR2_X1 U1068 ( .A(G1966), .B(G1981), .ZN(n980) );
  XNOR2_X1 U1069 ( .A(n981), .B(n980), .ZN(G229) );
  XOR2_X1 U1070 ( .A(KEYINPUT106), .B(G2678), .Z(n983) );
  XNOR2_X1 U1071 ( .A(G2072), .B(G2090), .ZN(n982) );
  XNOR2_X1 U1072 ( .A(n983), .B(n982), .ZN(n987) );
  XOR2_X1 U1073 ( .A(KEYINPUT43), .B(KEYINPUT105), .Z(n985) );
  XNOR2_X1 U1074 ( .A(G2067), .B(KEYINPUT42), .ZN(n984) );
  XNOR2_X1 U1075 ( .A(n985), .B(n984), .ZN(n986) );
  XOR2_X1 U1076 ( .A(n987), .B(n986), .Z(n990) );
  XOR2_X1 U1077 ( .A(G2096), .B(n988), .Z(n989) );
  XNOR2_X1 U1078 ( .A(n990), .B(n989), .ZN(n992) );
  XOR2_X1 U1079 ( .A(G2078), .B(G2084), .Z(n991) );
  XNOR2_X1 U1080 ( .A(n992), .B(n991), .ZN(G227) );
  XNOR2_X1 U1081 ( .A(n994), .B(n993), .ZN(n997) );
  XOR2_X1 U1082 ( .A(G301), .B(n995), .Z(n996) );
  XNOR2_X1 U1083 ( .A(n997), .B(n996), .ZN(n998) );
  XOR2_X1 U1084 ( .A(G286), .B(n998), .Z(n999) );
  NOR2_X1 U1085 ( .A1(G37), .A2(n999), .ZN(G397) );
  XOR2_X1 U1086 ( .A(n1000), .B(G162), .Z(n1003) );
  XNOR2_X1 U1087 ( .A(G160), .B(n1001), .ZN(n1002) );
  XNOR2_X1 U1088 ( .A(n1003), .B(n1002), .ZN(n1007) );
  XOR2_X1 U1089 ( .A(KEYINPUT46), .B(KEYINPUT111), .Z(n1005) );
  XNOR2_X1 U1090 ( .A(KEYINPUT110), .B(KEYINPUT48), .ZN(n1004) );
  XNOR2_X1 U1091 ( .A(n1005), .B(n1004), .ZN(n1006) );
  XOR2_X1 U1092 ( .A(n1007), .B(n1006), .Z(n1010) );
  XNOR2_X1 U1093 ( .A(G164), .B(n1008), .ZN(n1009) );
  XNOR2_X1 U1094 ( .A(n1010), .B(n1009), .ZN(n1027) );
  NAND2_X1 U1095 ( .A1(n1011), .A2(G130), .ZN(n1014) );
  NAND2_X1 U1096 ( .A1(G118), .A2(n1012), .ZN(n1013) );
  NAND2_X1 U1097 ( .A1(n1014), .A2(n1013), .ZN(n1021) );
  NAND2_X1 U1098 ( .A1(G142), .A2(n1015), .ZN(n1018) );
  NAND2_X1 U1099 ( .A1(G106), .A2(n519), .ZN(n1017) );
  NAND2_X1 U1100 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XOR2_X1 U1101 ( .A(n1019), .B(KEYINPUT45), .Z(n1020) );
  NOR2_X1 U1102 ( .A1(n1021), .A2(n1020), .ZN(n1023) );
  XNOR2_X1 U1103 ( .A(n1023), .B(n1022), .ZN(n1024) );
  XOR2_X1 U1104 ( .A(n1025), .B(n1024), .Z(n1026) );
  XNOR2_X1 U1105 ( .A(n1027), .B(n1026), .ZN(n1028) );
  NOR2_X1 U1106 ( .A1(G37), .A2(n1028), .ZN(n1029) );
  XNOR2_X1 U1107 ( .A(KEYINPUT112), .B(n1029), .ZN(G395) );
  OR2_X1 U1108 ( .A1(n1035), .A2(G401), .ZN(n1032) );
  NOR2_X1 U1109 ( .A1(G229), .A2(G227), .ZN(n1030) );
  XNOR2_X1 U1110 ( .A(KEYINPUT49), .B(n1030), .ZN(n1031) );
  NOR2_X1 U1111 ( .A1(n1032), .A2(n1031), .ZN(n1034) );
  NOR2_X1 U1112 ( .A1(G397), .A2(G395), .ZN(n1033) );
  NAND2_X1 U1113 ( .A1(n1034), .A2(n1033), .ZN(G225) );
  INV_X1 U1114 ( .A(G225), .ZN(G308) );
  INV_X1 U1115 ( .A(n1035), .ZN(G319) );
  INV_X1 U1116 ( .A(G108), .ZN(G238) );
endmodule

