//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 1 1 0 0 1 1 1 0 1 1 0 0 1 1 1 1 1 1 0 1 0 0 1 0 1 0 0 0 1 0 1 1 0 1 1 1 0 1 1 0 0 1 1 1 1 0 0 0 1 1 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n728, new_n729,
    new_n730, new_n732, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n821, new_n822, new_n824, new_n825, new_n826, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n887, new_n888, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n904, new_n905,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n948, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958;
  XNOR2_X1  g000(.A(G197gat), .B(G204gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(G211gat), .A2(G218gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n202), .B1(KEYINPUT22), .B2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G211gat), .ZN(new_n206));
  INV_X1    g005(.A(G218gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(new_n203), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n205), .A2(new_n210), .ZN(new_n211));
  OAI211_X1 g010(.A(new_n209), .B(new_n202), .C1(KEYINPUT22), .C2(new_n204), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT72), .ZN(new_n215));
  NAND2_X1  g014(.A1(G226gat), .A2(G233gat), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(G183gat), .A2(G190gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(G169gat), .A2(G176gat), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT26), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n219), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  NOR3_X1   g021(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n218), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT27), .ZN(new_n225));
  OAI21_X1  g024(.A(KEYINPUT66), .B1(new_n225), .B2(G183gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT66), .ZN(new_n227));
  INV_X1    g026(.A(G183gat), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n227), .A2(new_n228), .A3(KEYINPUT27), .ZN(new_n229));
  AND2_X1   g028(.A1(new_n226), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n228), .A2(KEYINPUT27), .ZN(new_n231));
  AND2_X1   g030(.A1(KEYINPUT65), .A2(G190gat), .ZN(new_n232));
  NOR2_X1   g031(.A1(KEYINPUT65), .A2(G190gat), .ZN(new_n233));
  NOR3_X1   g032(.A1(new_n231), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n230), .A2(new_n234), .A3(KEYINPUT67), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT67), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n226), .A2(new_n229), .ZN(new_n237));
  OR2_X1    g036(.A1(KEYINPUT65), .A2(G190gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n225), .A2(G183gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(KEYINPUT65), .A2(G190gat), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n238), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n236), .B1(new_n237), .B2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT28), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n235), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n232), .A2(new_n233), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n228), .A2(KEYINPUT27), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n239), .A2(new_n247), .ZN(new_n248));
  NOR3_X1   g047(.A1(new_n246), .A2(new_n248), .A3(new_n243), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n224), .B1(new_n244), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n218), .A2(KEYINPUT24), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT24), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n253), .A2(G183gat), .A3(G190gat), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n255), .B1(G183gat), .B2(G190gat), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT23), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n220), .B(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n256), .A2(new_n258), .A3(new_n219), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT25), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n220), .B(KEYINPUT23), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT64), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n219), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g062(.A1(KEYINPUT64), .A2(G169gat), .A3(G176gat), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n263), .A2(KEYINPUT25), .A3(new_n264), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n261), .A2(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n255), .B1(new_n246), .B2(G183gat), .ZN(new_n267));
  AOI22_X1  g066(.A1(new_n259), .A2(new_n260), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n217), .B1(new_n251), .B2(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(KEYINPUT71), .B(KEYINPUT29), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n271), .B1(new_n251), .B2(new_n268), .ZN(new_n272));
  AOI22_X1  g071(.A1(new_n215), .A2(new_n269), .B1(new_n272), .B2(new_n216), .ZN(new_n273));
  AND3_X1   g072(.A1(new_n272), .A2(new_n215), .A3(new_n216), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n214), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT29), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n276), .B1(new_n251), .B2(new_n268), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(new_n216), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n278), .A2(new_n213), .A3(new_n269), .ZN(new_n279));
  XNOR2_X1  g078(.A(G8gat), .B(G36gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(G64gat), .B(G92gat), .ZN(new_n281));
  XOR2_X1   g080(.A(new_n280), .B(new_n281), .Z(new_n282));
  NAND4_X1  g081(.A1(new_n275), .A2(KEYINPUT30), .A3(new_n279), .A4(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(KEYINPUT73), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n282), .B1(new_n275), .B2(new_n279), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n275), .A2(new_n279), .A3(new_n282), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT30), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AND3_X1   g088(.A1(new_n284), .A2(new_n286), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(G225gat), .A2(G233gat), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(G155gat), .A2(G162gat), .ZN(new_n293));
  INV_X1    g092(.A(G155gat), .ZN(new_n294));
  INV_X1    g093(.A(G162gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(G141gat), .B(G148gat), .ZN(new_n297));
  OAI211_X1 g096(.A(new_n293), .B(new_n296), .C1(new_n297), .C2(KEYINPUT2), .ZN(new_n298));
  INV_X1    g097(.A(G141gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(G148gat), .ZN(new_n300));
  INV_X1    g099(.A(G148gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(G141gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n296), .A2(new_n293), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n293), .A2(KEYINPUT2), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n298), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(G134gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(G127gat), .ZN(new_n309));
  INV_X1    g108(.A(G127gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(G134gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(G113gat), .B(G120gat), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n312), .B1(new_n313), .B2(KEYINPUT1), .ZN(new_n314));
  INV_X1    g113(.A(G120gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(G113gat), .ZN(new_n316));
  INV_X1    g115(.A(G113gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(G120gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  XNOR2_X1  g118(.A(G127gat), .B(G134gat), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT1), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n314), .A2(new_n322), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n307), .A2(new_n323), .ZN(new_n324));
  AOI22_X1  g123(.A1(new_n298), .A2(new_n306), .B1(new_n314), .B2(new_n322), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n292), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT76), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n326), .A2(new_n327), .A3(KEYINPUT5), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n307), .A2(new_n323), .ZN(new_n329));
  NAND4_X1  g128(.A1(new_n298), .A2(new_n314), .A3(new_n306), .A4(new_n322), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n291), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT5), .ZN(new_n332));
  OAI21_X1  g131(.A(KEYINPUT76), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n314), .A2(new_n322), .A3(KEYINPUT68), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT68), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n323), .A2(new_n335), .ZN(new_n336));
  AND3_X1   g135(.A1(new_n298), .A2(KEYINPUT75), .A3(new_n306), .ZN(new_n337));
  AOI21_X1  g136(.A(KEYINPUT75), .B1(new_n298), .B2(new_n306), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n334), .B(new_n336), .C1(new_n337), .C2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT4), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n307), .A2(KEYINPUT3), .ZN(new_n342));
  XOR2_X1   g141(.A(KEYINPUT74), .B(KEYINPUT3), .Z(new_n343));
  NAND3_X1  g142(.A1(new_n298), .A2(new_n306), .A3(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n342), .A2(new_n323), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n330), .A2(new_n340), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n345), .A2(new_n291), .A3(new_n346), .ZN(new_n347));
  OAI211_X1 g146(.A(new_n328), .B(new_n333), .C1(new_n341), .C2(new_n347), .ZN(new_n348));
  XOR2_X1   g147(.A(G1gat), .B(G29gat), .Z(new_n349));
  XNOR2_X1  g148(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n349), .B(new_n350), .ZN(new_n351));
  XNOR2_X1  g150(.A(G57gat), .B(G85gat), .ZN(new_n352));
  XOR2_X1   g151(.A(new_n351), .B(new_n352), .Z(new_n353));
  INV_X1    g152(.A(KEYINPUT78), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n354), .B1(new_n330), .B2(KEYINPUT4), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n355), .B1(new_n339), .B2(KEYINPUT4), .ZN(new_n356));
  AOI22_X1  g155(.A1(new_n307), .A2(KEYINPUT3), .B1(new_n322), .B2(new_n314), .ZN(new_n357));
  AOI211_X1 g156(.A(KEYINPUT5), .B(new_n292), .C1(new_n357), .C2(new_n344), .ZN(new_n358));
  AND2_X1   g157(.A1(new_n336), .A2(new_n334), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT75), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n307), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n298), .A2(KEYINPUT75), .A3(new_n306), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND4_X1  g162(.A1(new_n359), .A2(new_n354), .A3(new_n340), .A4(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n356), .A2(new_n358), .A3(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n348), .A2(new_n353), .A3(new_n365), .ZN(new_n366));
  XOR2_X1   g165(.A(KEYINPUT79), .B(KEYINPUT6), .Z(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n353), .B1(new_n348), .B2(new_n365), .ZN(new_n369));
  OAI21_X1  g168(.A(KEYINPUT80), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n348), .A2(new_n365), .ZN(new_n371));
  INV_X1    g170(.A(new_n353), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT80), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n373), .A2(new_n374), .A3(new_n367), .A4(new_n366), .ZN(new_n375));
  INV_X1    g174(.A(new_n367), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n369), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n370), .A2(new_n375), .A3(new_n377), .ZN(new_n378));
  AND3_X1   g177(.A1(new_n278), .A2(new_n213), .A3(new_n269), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n272), .A2(new_n216), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n269), .A2(new_n215), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n272), .A2(new_n215), .A3(new_n216), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n379), .B1(new_n384), .B2(new_n214), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT73), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n385), .A2(new_n386), .A3(KEYINPUT30), .A4(new_n282), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n290), .A2(KEYINPUT81), .A3(new_n378), .A4(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT81), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n387), .A2(new_n284), .A3(new_n286), .A4(new_n289), .ZN(new_n390));
  AND3_X1   g189(.A1(new_n370), .A2(new_n375), .A3(new_n377), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n389), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  XNOR2_X1  g191(.A(KEYINPUT31), .B(G50gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n393), .B(KEYINPUT84), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n394), .B(G106gat), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(KEYINPUT29), .B1(new_n211), .B2(new_n212), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n307), .B1(new_n397), .B2(KEYINPUT3), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT83), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  OAI211_X1 g199(.A(KEYINPUT83), .B(new_n307), .C1(new_n397), .C2(KEYINPUT3), .ZN(new_n401));
  NAND2_X1  g200(.A1(G228gat), .A2(G233gat), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n344), .A2(new_n271), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n402), .B1(new_n214), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n400), .A2(new_n401), .A3(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n270), .B1(new_n211), .B2(new_n212), .ZN(new_n406));
  INV_X1    g205(.A(new_n343), .ZN(new_n407));
  OAI211_X1 g206(.A(new_n362), .B(new_n361), .C1(new_n406), .C2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n214), .A2(new_n403), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n402), .B(KEYINPUT82), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(G22gat), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n405), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n413), .B1(new_n405), .B2(new_n412), .ZN(new_n416));
  NOR3_X1   g215(.A1(new_n415), .A2(new_n416), .A3(G78gat), .ZN(new_n417));
  INV_X1    g216(.A(G78gat), .ZN(new_n418));
  AND3_X1   g217(.A1(new_n400), .A2(new_n401), .A3(new_n404), .ZN(new_n419));
  INV_X1    g218(.A(new_n411), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n420), .B1(new_n408), .B2(new_n409), .ZN(new_n421));
  OAI21_X1  g220(.A(G22gat), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n418), .B1(new_n422), .B2(new_n414), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n396), .B1(new_n417), .B2(new_n423), .ZN(new_n424));
  OAI21_X1  g223(.A(G78gat), .B1(new_n415), .B2(new_n416), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n422), .A2(new_n418), .A3(new_n414), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n425), .A2(new_n426), .A3(new_n395), .ZN(new_n427));
  AND2_X1   g226(.A1(new_n424), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n259), .A2(new_n260), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n266), .A2(new_n267), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n336), .A2(new_n334), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n237), .A2(new_n241), .ZN(new_n433));
  AOI21_X1  g232(.A(KEYINPUT28), .B1(new_n433), .B2(KEYINPUT67), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n249), .B1(new_n434), .B2(new_n242), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n431), .B(new_n432), .C1(new_n435), .C2(new_n224), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n359), .B1(new_n251), .B2(new_n268), .ZN(new_n437));
  INV_X1    g236(.A(G227gat), .ZN(new_n438));
  INV_X1    g237(.A(G233gat), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n436), .A2(new_n437), .A3(new_n440), .ZN(new_n441));
  XOR2_X1   g240(.A(G71gat), .B(G99gat), .Z(new_n442));
  XNOR2_X1  g241(.A(G15gat), .B(G43gat), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n442), .B(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(KEYINPUT33), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n441), .A2(KEYINPUT32), .A3(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT69), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n441), .A2(KEYINPUT69), .A3(KEYINPUT32), .A4(new_n445), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n441), .A2(KEYINPUT32), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT33), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n441), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n451), .A2(new_n453), .A3(new_n444), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n450), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n436), .A2(new_n437), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n456), .B1(new_n438), .B2(new_n439), .ZN(new_n457));
  OR2_X1    g256(.A1(new_n457), .A2(KEYINPUT34), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(KEYINPUT34), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n455), .A2(new_n460), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n450), .A2(new_n459), .A3(new_n458), .A4(new_n454), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n428), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n388), .A2(new_n392), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(KEYINPUT35), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT85), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n390), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n285), .B1(new_n288), .B2(new_n287), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n469), .A2(KEYINPUT85), .A3(new_n387), .A4(new_n284), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n461), .A2(KEYINPUT70), .A3(new_n462), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT70), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n455), .A2(new_n460), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n424), .A2(new_n427), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT35), .ZN(new_n477));
  XNOR2_X1  g276(.A(new_n353), .B(KEYINPUT86), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n478), .B1(new_n365), .B2(new_n348), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n377), .B1(new_n368), .B2(new_n479), .ZN(new_n480));
  AND3_X1   g279(.A1(new_n476), .A2(new_n477), .A3(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n471), .A2(new_n475), .A3(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n356), .A2(new_n364), .A3(new_n345), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(new_n292), .ZN(new_n484));
  OR2_X1    g283(.A1(new_n484), .A2(KEYINPUT39), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n329), .A2(new_n330), .A3(new_n291), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(KEYINPUT39), .ZN(new_n487));
  XOR2_X1   g286(.A(new_n487), .B(KEYINPUT87), .Z(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(new_n484), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n485), .A2(new_n489), .A3(new_n478), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT40), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n485), .A2(KEYINPUT40), .A3(new_n489), .A4(new_n478), .ZN(new_n493));
  INV_X1    g292(.A(new_n479), .ZN(new_n494));
  AND3_X1   g293(.A1(new_n492), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n468), .A2(new_n470), .A3(new_n495), .ZN(new_n496));
  OAI211_X1 g295(.A(new_n287), .B(new_n377), .C1(new_n368), .C2(new_n479), .ZN(new_n497));
  XNOR2_X1  g296(.A(KEYINPUT88), .B(KEYINPUT37), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n282), .B1(new_n385), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n384), .A2(new_n213), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT37), .ZN(new_n501));
  AND2_X1   g300(.A1(new_n278), .A2(new_n269), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n501), .B1(new_n502), .B2(new_n214), .ZN(new_n503));
  AOI21_X1  g302(.A(KEYINPUT38), .B1(new_n500), .B2(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n497), .B1(new_n499), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n385), .A2(new_n498), .ZN(new_n506));
  INV_X1    g305(.A(new_n282), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n385), .A2(new_n501), .ZN(new_n509));
  OAI21_X1  g308(.A(KEYINPUT38), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n428), .B1(new_n505), .B2(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n461), .A2(KEYINPUT36), .A3(new_n462), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT36), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n472), .A2(new_n513), .A3(new_n474), .ZN(new_n514));
  AOI22_X1  g313(.A1(new_n496), .A2(new_n511), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  AND4_X1   g314(.A1(new_n387), .A2(new_n284), .A3(new_n286), .A4(new_n289), .ZN(new_n516));
  AOI21_X1  g315(.A(KEYINPUT81), .B1(new_n516), .B2(new_n378), .ZN(new_n517));
  NOR3_X1   g316(.A1(new_n390), .A2(new_n391), .A3(new_n389), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n428), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  AOI22_X1  g318(.A1(new_n466), .A2(new_n482), .B1(new_n515), .B2(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(KEYINPUT89), .B(G50gat), .ZN(new_n521));
  INV_X1    g320(.A(G43gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  OR2_X1    g322(.A1(new_n523), .A2(KEYINPUT90), .ZN(new_n524));
  INV_X1    g323(.A(G50gat), .ZN(new_n525));
  AOI22_X1  g324(.A1(new_n523), .A2(KEYINPUT90), .B1(G43gat), .B2(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(KEYINPUT15), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g326(.A1(G29gat), .A2(G36gat), .ZN(new_n528));
  XOR2_X1   g327(.A(new_n528), .B(KEYINPUT14), .Z(new_n529));
  NAND2_X1  g328(.A1(G29gat), .A2(G36gat), .ZN(new_n530));
  XOR2_X1   g329(.A(new_n530), .B(KEYINPUT91), .Z(new_n531));
  NAND2_X1  g330(.A1(new_n522), .A2(G50gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n525), .A2(G43gat), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n532), .A2(new_n533), .A3(KEYINPUT15), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n529), .A2(new_n531), .A3(new_n534), .ZN(new_n535));
  OR3_X1    g334(.A1(new_n527), .A2(KEYINPUT92), .A3(new_n535), .ZN(new_n536));
  OAI21_X1  g335(.A(KEYINPUT92), .B1(new_n527), .B2(new_n535), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n529), .A2(new_n530), .ZN(new_n538));
  INV_X1    g337(.A(new_n534), .ZN(new_n539));
  AOI22_X1  g338(.A1(new_n536), .A2(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(G15gat), .B(G22gat), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT16), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n541), .B1(new_n542), .B2(G1gat), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n543), .B1(G1gat), .B2(new_n541), .ZN(new_n544));
  INV_X1    g343(.A(G8gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n540), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n546), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n548), .B1(new_n540), .B2(KEYINPUT17), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n536), .A2(new_n537), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n538), .A2(new_n539), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT17), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n547), .B1(new_n549), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(G229gat), .A2(G233gat), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT18), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n555), .A2(KEYINPUT18), .A3(new_n556), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n540), .B(new_n546), .ZN(new_n561));
  XOR2_X1   g360(.A(new_n556), .B(KEYINPUT13), .Z(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n559), .A2(new_n560), .A3(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(G113gat), .B(G141gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(G197gat), .ZN(new_n566));
  XOR2_X1   g365(.A(KEYINPUT11), .B(G169gat), .Z(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  XOR2_X1   g367(.A(new_n568), .B(KEYINPUT12), .Z(new_n569));
  NAND2_X1  g368(.A1(new_n564), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n569), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n559), .A2(new_n571), .A3(new_n560), .A4(new_n563), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n520), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(G99gat), .A2(G106gat), .ZN(new_n576));
  INV_X1    g375(.A(G85gat), .ZN(new_n577));
  INV_X1    g376(.A(G92gat), .ZN(new_n578));
  AOI22_X1  g377(.A1(KEYINPUT8), .A2(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT97), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(G85gat), .A2(G92gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(KEYINPUT7), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  XOR2_X1   g383(.A(G99gat), .B(G106gat), .Z(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n584), .B(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(G57gat), .ZN(new_n588));
  AND2_X1   g387(.A1(new_n588), .A2(G64gat), .ZN(new_n589));
  OR2_X1    g388(.A1(new_n589), .A2(KEYINPUT94), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(KEYINPUT94), .ZN(new_n591));
  OAI211_X1 g390(.A(new_n590), .B(new_n591), .C1(new_n588), .C2(G64gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(G71gat), .B(G78gat), .ZN(new_n593));
  AOI21_X1  g392(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n594), .B(KEYINPUT93), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n592), .A2(new_n593), .A3(new_n595), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n588), .A2(G64gat), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n595), .B1(new_n589), .B2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n593), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n587), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n584), .B(new_n585), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(new_n601), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g405(.A(KEYINPUT99), .B1(new_n606), .B2(KEYINPUT10), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n587), .A2(KEYINPUT10), .A3(new_n602), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT99), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT10), .ZN(new_n610));
  NAND4_X1  g409(.A1(new_n603), .A2(new_n605), .A3(new_n609), .A4(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n607), .A2(new_n608), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(G230gat), .A2(G233gat), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n613), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n606), .A2(new_n615), .ZN(new_n616));
  AND2_X1   g415(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(G120gat), .B(G148gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(G176gat), .B(G204gat), .ZN(new_n619));
  XOR2_X1   g418(.A(new_n618), .B(new_n619), .Z(new_n620));
  OR2_X1    g419(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n614), .A2(new_n616), .A3(new_n620), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  AND2_X1   g423(.A1(G232gat), .A2(G233gat), .ZN(new_n625));
  AOI22_X1  g424(.A1(new_n552), .A2(new_n587), .B1(KEYINPUT41), .B2(new_n625), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n604), .B1(new_n552), .B2(new_n553), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n540), .A2(KEYINPUT17), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n626), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(G190gat), .B(G218gat), .ZN(new_n630));
  OR2_X1    g429(.A1(new_n630), .A2(KEYINPUT98), .ZN(new_n631));
  XNOR2_X1  g430(.A(G134gat), .B(G162gat), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  AND3_X1   g432(.A1(new_n629), .A2(new_n631), .A3(new_n633), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n633), .B1(new_n629), .B2(new_n631), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n630), .A2(KEYINPUT98), .ZN(new_n636));
  OR2_X1    g435(.A1(new_n625), .A2(KEYINPUT41), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  OR3_X1    g438(.A1(new_n634), .A2(new_n635), .A3(new_n639), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n639), .B1(new_n634), .B2(new_n635), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n548), .B1(KEYINPUT21), .B2(new_n602), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(KEYINPUT96), .ZN(new_n645));
  NAND2_X1  g444(.A1(G231gat), .A2(G233gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(KEYINPUT95), .ZN(new_n647));
  XOR2_X1   g446(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n645), .B(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n602), .A2(KEYINPUT21), .ZN(new_n651));
  XNOR2_X1  g450(.A(G127gat), .B(G155gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(G183gat), .B(G211gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(new_n655));
  OR2_X1    g454(.A1(new_n650), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n650), .A2(new_n655), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n643), .A2(new_n659), .ZN(new_n660));
  AND3_X1   g459(.A1(new_n575), .A2(new_n624), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n391), .B(KEYINPUT100), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(G1gat), .ZN(G1324gat));
  INV_X1    g463(.A(new_n471), .ZN(new_n665));
  XOR2_X1   g464(.A(KEYINPUT16), .B(G8gat), .Z(new_n666));
  NAND4_X1  g465(.A1(new_n661), .A2(KEYINPUT42), .A3(new_n665), .A4(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n661), .A2(new_n665), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(KEYINPUT102), .ZN(new_n669));
  AND2_X1   g468(.A1(new_n669), .A2(new_n666), .ZN(new_n670));
  XNOR2_X1  g469(.A(KEYINPUT101), .B(KEYINPUT42), .ZN(new_n671));
  OAI221_X1 g470(.A(new_n667), .B1(new_n545), .B2(new_n669), .C1(new_n670), .C2(new_n671), .ZN(G1325gat));
  INV_X1    g471(.A(G15gat), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n661), .A2(new_n673), .A3(new_n475), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n514), .A2(new_n512), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  AND2_X1   g475(.A1(new_n661), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n674), .B1(new_n677), .B2(new_n673), .ZN(G1326gat));
  NAND2_X1  g477(.A1(new_n661), .A2(new_n428), .ZN(new_n679));
  XNOR2_X1  g478(.A(KEYINPUT43), .B(G22gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(G1327gat));
  NAND2_X1  g480(.A1(new_n466), .A2(new_n482), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n496), .A2(new_n511), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n519), .A2(new_n683), .A3(new_n675), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n642), .B1(new_n682), .B2(new_n684), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n623), .A2(new_n658), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n687), .A2(new_n574), .ZN(new_n688));
  AND2_X1   g487(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(G29gat), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n689), .A2(new_n690), .A3(new_n662), .ZN(new_n691));
  XOR2_X1   g490(.A(new_n691), .B(KEYINPUT45), .Z(new_n692));
  NAND2_X1  g491(.A1(new_n685), .A2(KEYINPUT44), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT44), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n694), .B1(new_n520), .B2(new_n642), .ZN(new_n695));
  AND2_X1   g494(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  AND2_X1   g495(.A1(new_n696), .A2(new_n688), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n690), .B1(new_n697), .B2(new_n662), .ZN(new_n698));
  OR2_X1    g497(.A1(new_n692), .A2(new_n698), .ZN(G1328gat));
  INV_X1    g498(.A(new_n697), .ZN(new_n700));
  OAI21_X1  g499(.A(G36gat), .B1(new_n700), .B2(new_n471), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n687), .A2(new_n642), .A3(G36gat), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n575), .A2(new_n665), .A3(new_n702), .ZN(new_n703));
  XOR2_X1   g502(.A(new_n703), .B(KEYINPUT46), .Z(new_n704));
  NAND2_X1  g503(.A1(new_n701), .A2(new_n704), .ZN(G1329gat));
  OAI21_X1  g504(.A(G43gat), .B1(new_n700), .B2(new_n675), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n689), .A2(new_n522), .A3(new_n475), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT103), .ZN(new_n709));
  AOI21_X1  g508(.A(KEYINPUT47), .B1(new_n707), .B2(new_n709), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n708), .B(new_n710), .ZN(G1330gat));
  NAND3_X1  g510(.A1(new_n697), .A2(new_n428), .A3(new_n521), .ZN(new_n712));
  AND2_X1   g511(.A1(new_n689), .A2(new_n428), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n712), .B1(new_n521), .B2(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT48), .ZN(G1331gat));
  NAND3_X1  g514(.A1(new_n660), .A2(new_n574), .A3(new_n623), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT104), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n717), .A2(new_n520), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(new_n662), .ZN(new_n719));
  XNOR2_X1  g518(.A(KEYINPUT105), .B(G57gat), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n719), .B(new_n720), .ZN(G1332gat));
  NOR3_X1   g520(.A1(new_n717), .A2(new_n471), .A3(new_n520), .ZN(new_n722));
  NOR2_X1   g521(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n723));
  AND2_X1   g522(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n722), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n725), .B1(new_n722), .B2(new_n723), .ZN(G1333gat));
  INV_X1    g525(.A(G71gat), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n718), .A2(new_n727), .A3(new_n475), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n717), .A2(new_n675), .A3(new_n520), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n728), .B1(new_n729), .B2(new_n727), .ZN(new_n730));
  XOR2_X1   g529(.A(new_n730), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g530(.A1(new_n718), .A2(new_n428), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g532(.A1(new_n573), .A2(new_n658), .ZN(new_n734));
  INV_X1    g533(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n735), .A2(new_n624), .ZN(new_n736));
  AND2_X1   g535(.A1(new_n696), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(new_n662), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n577), .B1(new_n738), .B2(KEYINPUT106), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n739), .B1(KEYINPUT106), .B2(new_n738), .ZN(new_n740));
  OAI21_X1  g539(.A(KEYINPUT107), .B1(new_n520), .B2(new_n642), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n682), .A2(new_n684), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT107), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n742), .A2(new_n743), .A3(new_n643), .ZN(new_n744));
  AND4_X1   g543(.A1(KEYINPUT51), .A2(new_n741), .A3(new_n734), .A4(new_n744), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n735), .B1(new_n685), .B2(new_n743), .ZN(new_n746));
  AOI21_X1  g545(.A(KEYINPUT51), .B1(new_n746), .B2(new_n741), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(KEYINPUT108), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT108), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n662), .A2(new_n623), .A3(new_n577), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n740), .B1(new_n752), .B2(new_n753), .ZN(G1336gat));
  AOI21_X1  g553(.A(new_n578), .B1(new_n737), .B2(new_n665), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n755), .A2(KEYINPUT52), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n665), .A2(new_n578), .A3(new_n623), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n756), .B1(new_n752), .B2(new_n757), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n748), .A2(new_n757), .ZN(new_n759));
  OAI21_X1  g558(.A(KEYINPUT52), .B1(new_n755), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n758), .A2(new_n760), .ZN(G1337gat));
  INV_X1    g560(.A(new_n475), .ZN(new_n762));
  NOR3_X1   g561(.A1(new_n624), .A2(G99gat), .A3(new_n762), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n749), .A2(new_n751), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n737), .A2(new_n676), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(G99gat), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT109), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n764), .A2(new_n766), .A3(KEYINPUT109), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(G1338gat));
  NOR3_X1   g570(.A1(new_n624), .A2(G106gat), .A3(new_n476), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n749), .A2(new_n751), .A3(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT53), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n693), .A2(new_n695), .A3(new_n428), .A4(new_n736), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(G106gat), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n773), .A2(new_n774), .A3(new_n776), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n772), .B1(new_n745), .B2(new_n747), .ZN(new_n778));
  AOI22_X1  g577(.A1(new_n778), .A2(KEYINPUT110), .B1(G106gat), .B2(new_n775), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT110), .ZN(new_n780));
  OAI211_X1 g579(.A(new_n780), .B(new_n772), .C1(new_n745), .C2(new_n747), .ZN(new_n781));
  AOI211_X1 g580(.A(KEYINPUT111), .B(new_n774), .C1(new_n779), .C2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT111), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n778), .A2(KEYINPUT110), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n784), .A2(new_n781), .A3(new_n776), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n783), .B1(new_n785), .B2(KEYINPUT53), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n777), .B1(new_n782), .B2(new_n786), .ZN(G1339gat));
  NAND2_X1  g586(.A1(new_n662), .A2(new_n471), .ZN(new_n788));
  AND2_X1   g587(.A1(new_n611), .A2(new_n608), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n615), .B1(new_n789), .B2(new_n607), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT54), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n620), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n789), .A2(new_n615), .A3(new_n607), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n614), .A2(KEYINPUT54), .A3(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n792), .A2(new_n794), .A3(KEYINPUT55), .ZN(new_n795));
  AND2_X1   g594(.A1(new_n795), .A2(new_n622), .ZN(new_n796));
  AOI21_X1  g595(.A(KEYINPUT55), .B1(new_n792), .B2(new_n794), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT112), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  AOI211_X1 g598(.A(KEYINPUT112), .B(KEYINPUT55), .C1(new_n792), .C2(new_n794), .ZN(new_n800));
  OAI211_X1 g599(.A(new_n796), .B(new_n573), .C1(new_n799), .C2(new_n800), .ZN(new_n801));
  OAI22_X1  g600(.A1(new_n555), .A2(new_n556), .B1(new_n561), .B2(new_n562), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(new_n568), .ZN(new_n803));
  AND2_X1   g602(.A1(new_n572), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n623), .A2(new_n804), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n643), .B1(new_n801), .B2(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n796), .B1(new_n799), .B2(new_n800), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n804), .A2(new_n640), .A3(new_n641), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n659), .B1(new_n806), .B2(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n660), .A2(new_n574), .A3(new_n624), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n788), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n812), .A2(new_n464), .ZN(new_n813));
  AOI21_X1  g612(.A(G113gat), .B1(new_n813), .B2(new_n573), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n810), .A2(new_n811), .ZN(new_n815));
  INV_X1    g614(.A(new_n788), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n762), .A2(new_n428), .ZN(new_n817));
  AND3_X1   g616(.A1(new_n815), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n574), .A2(new_n317), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n814), .B1(new_n818), .B2(new_n819), .ZN(G1340gat));
  AOI21_X1  g619(.A(G120gat), .B1(new_n813), .B2(new_n623), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n624), .A2(new_n315), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n821), .B1(new_n818), .B2(new_n822), .ZN(G1341gat));
  INV_X1    g622(.A(new_n818), .ZN(new_n824));
  OAI21_X1  g623(.A(G127gat), .B1(new_n824), .B2(new_n659), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n813), .A2(new_n310), .A3(new_n658), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(G1342gat));
  NOR2_X1   g626(.A1(new_n642), .A2(G134gat), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n815), .A2(new_n464), .A3(new_n816), .A4(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(KEYINPUT113), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT56), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT113), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n812), .A2(new_n832), .A3(new_n464), .A4(new_n828), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n830), .A2(new_n831), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(KEYINPUT114), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT114), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n830), .A2(new_n836), .A3(new_n831), .A4(new_n833), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n308), .B1(new_n818), .B2(new_n643), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n830), .A2(new_n833), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n839), .B1(new_n840), .B2(KEYINPUT56), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n838), .A2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT115), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n838), .A2(new_n841), .A3(KEYINPUT115), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(G1343gat));
  INV_X1    g645(.A(KEYINPUT57), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n815), .A2(new_n847), .A3(new_n428), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n788), .A2(new_n676), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT116), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n795), .A2(new_n622), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n850), .B1(new_n851), .B2(new_n797), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n792), .A2(new_n794), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT55), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n855), .A2(KEYINPUT116), .A3(new_n622), .A4(new_n795), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n852), .A2(new_n573), .A3(new_n856), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n643), .B1(new_n857), .B2(new_n805), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n659), .B1(new_n858), .B2(new_n809), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n476), .B1(new_n859), .B2(new_n811), .ZN(new_n860));
  OAI211_X1 g659(.A(new_n848), .B(new_n849), .C1(new_n860), .C2(new_n847), .ZN(new_n861));
  OAI21_X1  g660(.A(G141gat), .B1(new_n861), .B2(new_n574), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n676), .A2(new_n476), .ZN(new_n863));
  AND2_X1   g662(.A1(new_n812), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n573), .A2(new_n299), .ZN(new_n865));
  XNOR2_X1  g664(.A(new_n865), .B(KEYINPUT117), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n862), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g667(.A(KEYINPUT118), .B(KEYINPUT58), .ZN(new_n869));
  XNOR2_X1  g668(.A(new_n868), .B(new_n869), .ZN(G1344gat));
  NAND3_X1  g669(.A1(new_n864), .A2(new_n301), .A3(new_n623), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT59), .ZN(new_n872));
  AOI211_X1 g671(.A(new_n847), .B(new_n476), .C1(new_n810), .C2(new_n811), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(KEYINPUT119), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n815), .A2(KEYINPUT57), .A3(new_n428), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT119), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  OAI211_X1 g676(.A(new_n874), .B(new_n877), .C1(KEYINPUT57), .C2(new_n860), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n878), .A2(new_n623), .A3(new_n849), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n872), .B1(new_n879), .B2(G148gat), .ZN(new_n880));
  INV_X1    g679(.A(new_n861), .ZN(new_n881));
  AOI211_X1 g680(.A(KEYINPUT59), .B(new_n301), .C1(new_n881), .C2(new_n623), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n871), .B1(new_n880), .B2(new_n882), .ZN(G1345gat));
  OAI21_X1  g682(.A(G155gat), .B1(new_n861), .B2(new_n659), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n864), .A2(new_n294), .A3(new_n658), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(G1346gat));
  AOI21_X1  g685(.A(G162gat), .B1(new_n864), .B2(new_n643), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n642), .A2(new_n295), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n887), .B1(new_n881), .B2(new_n888), .ZN(G1347gat));
  INV_X1    g688(.A(KEYINPUT121), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n815), .A2(new_n817), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n662), .A2(new_n471), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n890), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(new_n893), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n891), .A2(new_n890), .A3(new_n892), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g695(.A(G169gat), .B1(new_n896), .B2(new_n574), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n662), .B1(new_n810), .B2(new_n811), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n471), .A2(new_n428), .A3(new_n463), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n900), .A2(G169gat), .A3(new_n574), .ZN(new_n901));
  XNOR2_X1  g700(.A(new_n901), .B(KEYINPUT120), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n897), .A2(new_n902), .ZN(G1348gat));
  OAI21_X1  g702(.A(G176gat), .B1(new_n896), .B2(new_n624), .ZN(new_n904));
  OR2_X1    g703(.A1(new_n624), .A2(G176gat), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n904), .B1(new_n900), .B2(new_n905), .ZN(G1349gat));
  AND3_X1   g705(.A1(new_n891), .A2(new_n890), .A3(new_n892), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n907), .A2(new_n893), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n228), .B1(new_n908), .B2(new_n658), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n900), .A2(new_n248), .A3(new_n659), .ZN(new_n910));
  OAI21_X1  g709(.A(KEYINPUT60), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g710(.A(G183gat), .B1(new_n896), .B2(new_n659), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT60), .ZN(new_n913));
  INV_X1    g712(.A(new_n910), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n911), .A2(new_n915), .ZN(G1350gat));
  NAND3_X1  g715(.A1(new_n894), .A2(new_n643), .A3(new_n895), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT61), .ZN(new_n918));
  AND3_X1   g717(.A1(new_n917), .A2(new_n918), .A3(G190gat), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n918), .B1(new_n917), .B2(G190gat), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n643), .A2(new_n245), .ZN(new_n921));
  OAI22_X1  g720(.A1(new_n919), .A2(new_n920), .B1(new_n900), .B2(new_n921), .ZN(G1351gat));
  NAND2_X1  g721(.A1(new_n863), .A2(new_n665), .ZN(new_n923));
  XOR2_X1   g722(.A(new_n923), .B(KEYINPUT122), .Z(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(new_n898), .ZN(new_n925));
  INV_X1    g724(.A(new_n925), .ZN(new_n926));
  XNOR2_X1  g725(.A(KEYINPUT123), .B(G197gat), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n926), .A2(new_n573), .A3(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT124), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n892), .A2(new_n675), .ZN(new_n930));
  INV_X1    g729(.A(new_n930), .ZN(new_n931));
  AND2_X1   g730(.A1(new_n878), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n929), .B1(new_n932), .B2(new_n573), .ZN(new_n933));
  NAND4_X1  g732(.A1(new_n878), .A2(new_n929), .A3(new_n573), .A4(new_n931), .ZN(new_n934));
  INV_X1    g733(.A(new_n927), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n928), .B1(new_n933), .B2(new_n936), .ZN(G1352gat));
  NOR3_X1   g736(.A1(new_n925), .A2(G204gat), .A3(new_n624), .ZN(new_n938));
  XNOR2_X1  g737(.A(new_n938), .B(KEYINPUT62), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n878), .A2(new_n623), .A3(new_n931), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(KEYINPUT125), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(G204gat), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n940), .A2(KEYINPUT125), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n939), .B1(new_n942), .B2(new_n943), .ZN(G1353gat));
  NAND3_X1  g743(.A1(new_n926), .A2(new_n206), .A3(new_n658), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n878), .A2(new_n658), .A3(new_n931), .ZN(new_n946));
  AND3_X1   g745(.A1(new_n946), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n947));
  AOI21_X1  g746(.A(KEYINPUT63), .B1(new_n946), .B2(G211gat), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n945), .B1(new_n947), .B2(new_n948), .ZN(G1354gat));
  OAI22_X1  g748(.A1(new_n873), .A2(KEYINPUT119), .B1(new_n860), .B2(KEYINPUT57), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n875), .A2(new_n876), .ZN(new_n951));
  OAI211_X1 g750(.A(new_n643), .B(new_n931), .C1(new_n950), .C2(new_n951), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n952), .A2(G218gat), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n926), .A2(new_n207), .A3(new_n643), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT126), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n953), .A2(KEYINPUT126), .A3(new_n954), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(G1355gat));
endmodule


