//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 1 1 0 0 0 0 1 1 1 0 1 1 1 0 1 0 0 1 0 1 0 1 0 1 1 1 1 0 1 1 0 1 1 1 0 0 1 0 1 1 0 1 0 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:01 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n728, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n910, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978;
  INV_X1    g000(.A(G140), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G125), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT16), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G125), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G140), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT74), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n188), .A2(new_n192), .A3(new_n193), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n187), .A2(KEYINPUT74), .A3(G125), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n190), .B1(new_n196), .B2(new_n189), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G146), .ZN(new_n198));
  INV_X1    g012(.A(G146), .ZN(new_n199));
  OAI211_X1 g013(.A(new_n199), .B(new_n190), .C1(new_n196), .C2(new_n189), .ZN(new_n200));
  AND2_X1   g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G110), .ZN(new_n202));
  XNOR2_X1  g016(.A(KEYINPUT67), .B(G119), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G128), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(KEYINPUT23), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT73), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n206), .B1(new_n203), .B2(G128), .ZN(new_n207));
  INV_X1    g021(.A(G119), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(KEYINPUT67), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT67), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G119), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G128), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n212), .A2(KEYINPUT73), .A3(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n205), .A2(new_n207), .A3(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n213), .A2(KEYINPUT23), .A3(G119), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n202), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n204), .B1(new_n208), .B2(G128), .ZN(new_n218));
  XNOR2_X1  g032(.A(KEYINPUT24), .B(G110), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OR3_X1    g034(.A1(new_n201), .A2(new_n217), .A3(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n215), .A2(new_n202), .A3(new_n216), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n218), .A2(new_n219), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AND2_X1   g038(.A1(new_n188), .A2(new_n192), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(new_n199), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n224), .A2(new_n198), .A3(new_n226), .ZN(new_n227));
  XNOR2_X1  g041(.A(KEYINPUT22), .B(G137), .ZN(new_n228));
  INV_X1    g042(.A(G953), .ZN(new_n229));
  AND3_X1   g043(.A1(new_n229), .A2(G221), .A3(G234), .ZN(new_n230));
  XOR2_X1   g044(.A(new_n228), .B(new_n230), .Z(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n221), .A2(new_n227), .A3(new_n232), .ZN(new_n233));
  AND3_X1   g047(.A1(new_n224), .A2(new_n198), .A3(new_n226), .ZN(new_n234));
  NOR3_X1   g048(.A1(new_n201), .A2(new_n217), .A3(new_n220), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n231), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n233), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT25), .ZN(new_n238));
  INV_X1    g052(.A(G902), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n237), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G217), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n241), .B1(G234), .B2(new_n239), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n238), .B1(new_n237), .B2(new_n239), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n242), .A2(G902), .ZN(new_n246));
  AND2_X1   g060(.A1(new_n237), .A2(new_n246), .ZN(new_n247));
  OR2_X1    g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  NOR2_X1   g062(.A1(G472), .A2(G902), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT68), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n213), .A2(KEYINPUT1), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n199), .A2(G143), .ZN(new_n252));
  INV_X1    g066(.A(G143), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G146), .ZN(new_n254));
  AND3_X1   g068(.A1(new_n251), .A2(new_n252), .A3(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT66), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n256), .B(KEYINPUT1), .C1(new_n253), .C2(G146), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n256), .B1(new_n252), .B2(KEYINPUT1), .ZN(new_n259));
  OAI21_X1  g073(.A(G128), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n252), .A2(new_n254), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n255), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(G134), .ZN(new_n263));
  OAI21_X1  g077(.A(KEYINPUT65), .B1(new_n263), .B2(G137), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT65), .ZN(new_n265));
  INV_X1    g079(.A(G137), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n265), .A2(new_n266), .A3(G134), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n263), .A2(G137), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n264), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(G131), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT11), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n271), .B1(new_n263), .B2(G137), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n266), .A2(KEYINPUT11), .A3(G134), .ZN(new_n273));
  INV_X1    g087(.A(G131), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n272), .A2(new_n273), .A3(new_n274), .A4(new_n268), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n270), .A2(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n250), .B1(new_n262), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n255), .ZN(new_n278));
  OAI21_X1  g092(.A(KEYINPUT1), .B1(new_n253), .B2(G146), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(KEYINPUT66), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n213), .B1(new_n280), .B2(new_n257), .ZN(new_n281));
  XNOR2_X1  g095(.A(G143), .B(G146), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n278), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  AND2_X1   g097(.A1(new_n270), .A2(new_n275), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n283), .A2(new_n284), .A3(KEYINPUT68), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n272), .A2(new_n273), .A3(new_n268), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(G131), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(new_n275), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT0), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(new_n213), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(KEYINPUT0), .A2(G128), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n261), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n282), .A2(new_n292), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n288), .A2(new_n296), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n277), .A2(KEYINPUT30), .A3(new_n285), .A4(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n209), .A2(new_n211), .A3(G116), .ZN(new_n299));
  INV_X1    g113(.A(G116), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(G119), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  XNOR2_X1  g116(.A(KEYINPUT2), .B(G113), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(new_n303), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n305), .A2(new_n299), .A3(new_n301), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT30), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n262), .A2(new_n276), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n261), .A2(new_n293), .ZN(new_n310));
  AOI22_X1  g124(.A1(new_n252), .A2(new_n254), .B1(new_n290), .B2(new_n292), .ZN(new_n311));
  OAI21_X1  g125(.A(KEYINPUT64), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT64), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n294), .A2(new_n313), .A3(new_n295), .ZN(new_n314));
  AOI22_X1  g128(.A1(new_n312), .A2(new_n314), .B1(new_n275), .B2(new_n287), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n308), .B1(new_n309), .B2(new_n315), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n298), .A2(new_n307), .A3(new_n316), .ZN(new_n317));
  NOR2_X1   g131(.A1(G237), .A2(G953), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G210), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT27), .ZN(new_n320));
  XNOR2_X1  g134(.A(new_n319), .B(new_n320), .ZN(new_n321));
  XNOR2_X1  g135(.A(new_n321), .B(KEYINPUT69), .ZN(new_n322));
  XNOR2_X1  g136(.A(KEYINPUT26), .B(G101), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n322), .B(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n307), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n277), .A2(new_n325), .A3(new_n285), .A4(new_n297), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n317), .A2(new_n324), .A3(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT70), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n317), .A2(KEYINPUT70), .A3(new_n324), .A4(new_n326), .ZN(new_n330));
  AND3_X1   g144(.A1(new_n329), .A2(KEYINPUT31), .A3(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n324), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n283), .A2(new_n284), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n333), .A2(new_n325), .A3(new_n297), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT28), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT71), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n334), .A2(KEYINPUT71), .A3(new_n335), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n307), .B1(new_n309), .B2(new_n315), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n335), .B1(new_n326), .B2(new_n341), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n332), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT31), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n317), .A2(new_n344), .A3(new_n324), .A4(new_n326), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n249), .B1(new_n331), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(KEYINPUT32), .ZN(new_n348));
  INV_X1    g162(.A(new_n249), .ZN(new_n349));
  AND2_X1   g163(.A1(new_n343), .A2(new_n345), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n329), .A2(KEYINPUT31), .A3(new_n330), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n349), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT32), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n348), .A2(new_n354), .ZN(new_n355));
  NOR3_X1   g169(.A1(new_n340), .A2(new_n342), .A3(new_n332), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n324), .B1(new_n317), .B2(new_n326), .ZN(new_n357));
  NOR3_X1   g171(.A1(new_n356), .A2(KEYINPUT29), .A3(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT72), .ZN(new_n359));
  INV_X1    g173(.A(new_n339), .ZN(new_n360));
  AOI21_X1  g174(.A(KEYINPUT71), .B1(new_n334), .B2(new_n335), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n359), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  AOI22_X1  g176(.A1(new_n333), .A2(new_n250), .B1(new_n288), .B2(new_n296), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n325), .B1(new_n363), .B2(new_n285), .ZN(new_n364));
  INV_X1    g178(.A(new_n326), .ZN(new_n365));
  OAI21_X1  g179(.A(KEYINPUT28), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n338), .A2(KEYINPUT72), .A3(new_n339), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n362), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n324), .A2(KEYINPUT29), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n239), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(G472), .B1(new_n358), .B2(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n248), .B1(new_n355), .B2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(G469), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT75), .ZN(new_n374));
  XNOR2_X1  g188(.A(new_n288), .B(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(G104), .ZN(new_n376));
  OAI21_X1  g190(.A(KEYINPUT3), .B1(new_n376), .B2(G107), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT3), .ZN(new_n378));
  INV_X1    g192(.A(G107), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n378), .A2(new_n379), .A3(G104), .ZN(new_n380));
  INV_X1    g194(.A(G101), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n376), .A2(G107), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n377), .A2(new_n380), .A3(new_n381), .A4(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n376), .A2(G107), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n379), .A2(G104), .ZN(new_n385));
  OAI21_X1  g199(.A(G101), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n383), .A2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT10), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  AOI22_X1  g203(.A1(new_n279), .A2(G128), .B1(new_n252), .B2(new_n254), .ZN(new_n390));
  OAI211_X1 g204(.A(new_n383), .B(new_n386), .C1(new_n390), .C2(new_n255), .ZN(new_n391));
  AOI22_X1  g205(.A1(new_n283), .A2(new_n389), .B1(new_n391), .B2(new_n388), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n377), .A2(new_n380), .A3(new_n382), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(G101), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n394), .A2(KEYINPUT4), .A3(new_n383), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT4), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n393), .A2(new_n396), .A3(G101), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n395), .A2(new_n296), .A3(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n375), .A2(new_n392), .A3(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n387), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n391), .B1(new_n283), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(new_n288), .ZN(new_n402));
  AOI21_X1  g216(.A(KEYINPUT12), .B1(new_n288), .B2(KEYINPUT76), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n403), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n405), .B1(new_n401), .B2(new_n288), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n399), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  XNOR2_X1  g221(.A(G110), .B(G140), .ZN(new_n408));
  INV_X1    g222(.A(G227), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n409), .A2(G953), .ZN(new_n410));
  XOR2_X1   g224(.A(new_n408), .B(new_n410), .Z(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n407), .A2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT77), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n283), .A2(new_n389), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n391), .A2(new_n388), .ZN(new_n416));
  AND4_X1   g230(.A1(new_n414), .A2(new_n415), .A3(new_n398), .A4(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n414), .B1(new_n392), .B2(new_n398), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n288), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n419), .A2(new_n399), .A3(new_n411), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n413), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n373), .B1(new_n421), .B2(new_n239), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n288), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n415), .A2(new_n398), .A3(new_n416), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(KEYINPUT77), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n392), .A2(new_n414), .A3(new_n398), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n424), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n399), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n412), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  OAI211_X1 g244(.A(new_n399), .B(new_n411), .C1(new_n404), .C2(new_n406), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT78), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n432), .A2(new_n433), .A3(new_n373), .A4(new_n239), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(G902), .B1(new_n430), .B2(new_n431), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n433), .B1(new_n436), .B2(new_n373), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n423), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(G221), .ZN(new_n439));
  XNOR2_X1  g253(.A(KEYINPUT9), .B(G234), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n439), .B1(new_n441), .B2(new_n239), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n438), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT85), .ZN(new_n445));
  XNOR2_X1  g259(.A(G113), .B(G122), .ZN(new_n446));
  XNOR2_X1  g260(.A(new_n446), .B(new_n376), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT19), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT83), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n196), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n194), .A2(KEYINPUT83), .A3(new_n195), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n448), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n225), .A2(KEYINPUT19), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n199), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n318), .A2(G214), .ZN(new_n455));
  NOR2_X1   g269(.A1(KEYINPUT82), .A2(G143), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n318), .B(G214), .C1(KEYINPUT82), .C2(G143), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(G131), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n457), .A2(new_n458), .A3(new_n274), .ZN(new_n461));
  AOI22_X1  g275(.A1(new_n197), .A2(G146), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n454), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n450), .A2(G146), .A3(new_n451), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n226), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n457), .A2(new_n458), .A3(KEYINPUT84), .ZN(new_n466));
  NAND2_X1  g280(.A1(KEYINPUT18), .A2(G131), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n466), .B(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n447), .B1(new_n463), .B2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT17), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n460), .A2(new_n471), .A3(new_n461), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n459), .A2(KEYINPUT17), .A3(G131), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n472), .A2(new_n198), .A3(new_n200), .A4(new_n473), .ZN(new_n474));
  AND3_X1   g288(.A1(new_n469), .A2(new_n474), .A3(new_n447), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n445), .B1(new_n470), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g290(.A1(G475), .A2(G902), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n469), .A2(new_n474), .A3(new_n447), .ZN(new_n478));
  AOI22_X1  g292(.A1(new_n454), .A2(new_n462), .B1(new_n465), .B2(new_n468), .ZN(new_n479));
  OAI211_X1 g293(.A(KEYINPUT85), .B(new_n478), .C1(new_n479), .C2(new_n447), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n476), .A2(new_n477), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(KEYINPUT20), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT86), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n481), .A2(KEYINPUT86), .A3(KEYINPUT20), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT20), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n486), .B(new_n477), .C1(new_n470), .C2(new_n475), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n484), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(G214), .B1(G237), .B2(G902), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n296), .A2(G125), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n491), .B1(new_n262), .B2(G125), .ZN(new_n492));
  XNOR2_X1  g306(.A(KEYINPUT80), .B(G224), .ZN(new_n493));
  OR2_X1    g307(.A1(new_n493), .A2(G953), .ZN(new_n494));
  AND2_X1   g308(.A1(new_n494), .A2(KEYINPUT7), .ZN(new_n495));
  OR2_X1    g309(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n299), .A2(KEYINPUT5), .A3(new_n301), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n497), .B(G113), .C1(KEYINPUT5), .C2(new_n299), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n498), .A2(new_n306), .A3(new_n400), .ZN(new_n499));
  XNOR2_X1  g313(.A(G110), .B(G122), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n307), .A2(new_n397), .ZN(new_n501));
  INV_X1    g315(.A(new_n395), .ZN(new_n502));
  OAI211_X1 g316(.A(new_n499), .B(new_n500), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n500), .B(KEYINPUT8), .ZN(new_n504));
  AND3_X1   g318(.A1(new_n498), .A2(new_n306), .A3(new_n400), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n400), .B1(new_n498), .B2(new_n306), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n492), .A2(KEYINPUT7), .A3(new_n494), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n496), .A2(new_n503), .A3(new_n507), .A4(new_n508), .ZN(new_n509));
  AND2_X1   g323(.A1(new_n509), .A2(new_n239), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n499), .B1(new_n501), .B2(new_n502), .ZN(new_n511));
  INV_X1    g325(.A(new_n500), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n511), .A2(KEYINPUT79), .A3(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n513), .A2(KEYINPUT6), .A3(new_n503), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n492), .B(new_n494), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT6), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n511), .A2(KEYINPUT79), .A3(new_n516), .A4(new_n512), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n514), .A2(new_n515), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n510), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g333(.A(G210), .B1(G237), .B2(G902), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n520), .B(KEYINPUT81), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n510), .A2(new_n518), .A3(new_n520), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n490), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  AND2_X1   g338(.A1(new_n469), .A2(new_n474), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n525), .A2(new_n447), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(KEYINPUT87), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(new_n239), .ZN(new_n528));
  NOR3_X1   g342(.A1(new_n526), .A2(KEYINPUT87), .A3(new_n475), .ZN(new_n529));
  OAI21_X1  g343(.A(G475), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT92), .ZN(new_n531));
  OAI21_X1  g345(.A(KEYINPUT89), .B1(new_n213), .B2(G143), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT89), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n533), .A2(new_n253), .A3(G128), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT13), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n213), .A2(G143), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n535), .A2(new_n536), .ZN(new_n540));
  OAI21_X1  g354(.A(G134), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  AND3_X1   g355(.A1(new_n535), .A2(new_n263), .A3(new_n538), .ZN(new_n542));
  OAI21_X1  g356(.A(KEYINPUT88), .B1(new_n300), .B2(G122), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT88), .ZN(new_n544));
  INV_X1    g358(.A(G122), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n544), .A2(new_n545), .A3(G116), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n300), .A2(G122), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(G107), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n547), .A2(new_n379), .A3(new_n548), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n542), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  AND3_X1   g366(.A1(new_n547), .A2(new_n379), .A3(new_n548), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT90), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n554), .B1(new_n548), .B2(KEYINPUT14), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n548), .A2(KEYINPUT14), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT14), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n557), .A2(new_n300), .A3(KEYINPUT90), .A4(G122), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n547), .A2(new_n555), .A3(new_n556), .A4(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n553), .B1(G107), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n535), .A2(new_n538), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(G134), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n535), .A2(new_n263), .A3(new_n538), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AOI22_X1  g378(.A1(new_n541), .A2(new_n552), .B1(new_n560), .B2(new_n564), .ZN(new_n565));
  NOR3_X1   g379(.A1(new_n440), .A2(new_n241), .A3(G953), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n531), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n552), .A2(new_n541), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n559), .A2(G107), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n564), .A2(new_n551), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n566), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n571), .A2(KEYINPUT92), .A3(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n568), .A2(new_n570), .A3(new_n566), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(KEYINPUT91), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT91), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n568), .A2(new_n570), .A3(new_n576), .A4(new_n566), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n567), .A2(new_n573), .A3(new_n575), .A4(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(new_n239), .ZN(new_n579));
  INV_X1    g393(.A(G478), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n580), .A2(KEYINPUT15), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n581), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n578), .A2(new_n239), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(G952), .ZN(new_n586));
  AOI211_X1 g400(.A(G953), .B(new_n586), .C1(G234), .C2(G237), .ZN(new_n587));
  XNOR2_X1  g401(.A(KEYINPUT21), .B(G898), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n588), .B(KEYINPUT93), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  AOI211_X1 g404(.A(new_n239), .B(new_n229), .C1(G234), .C2(G237), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n587), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n585), .A2(new_n592), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n488), .A2(new_n524), .A3(new_n530), .A4(new_n593), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n444), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n372), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n596), .B(G101), .ZN(G3));
  OAI21_X1  g411(.A(new_n239), .B1(new_n331), .B2(new_n346), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n352), .B1(new_n598), .B2(G472), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n411), .B1(new_n419), .B2(new_n399), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n399), .A2(new_n411), .ZN(new_n601));
  INV_X1    g415(.A(new_n404), .ZN(new_n602));
  INV_X1    g416(.A(new_n406), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  OAI211_X1 g418(.A(new_n373), .B(new_n239), .C1(new_n600), .C2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(KEYINPUT78), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(new_n434), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n442), .B1(new_n607), .B2(new_n423), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n245), .A2(new_n247), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n599), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  XOR2_X1   g424(.A(new_n610), .B(KEYINPUT94), .Z(new_n611));
  NAND2_X1  g425(.A1(new_n488), .A2(new_n530), .ZN(new_n612));
  INV_X1    g426(.A(new_n523), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n520), .B1(new_n510), .B2(new_n518), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n489), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n615), .A2(new_n592), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n579), .A2(G478), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT33), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n618), .B1(new_n571), .B2(new_n572), .ZN(new_n619));
  AOI22_X1  g433(.A1(new_n578), .A2(new_n618), .B1(new_n574), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n239), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n617), .B1(new_n621), .B2(G478), .ZN(new_n622));
  AND3_X1   g436(.A1(new_n612), .A2(new_n616), .A3(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n611), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(KEYINPUT95), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(KEYINPUT34), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(G104), .ZN(G6));
  INV_X1    g442(.A(KEYINPUT96), .ZN(new_n629));
  AND3_X1   g443(.A1(new_n481), .A2(KEYINPUT86), .A3(KEYINPUT20), .ZN(new_n630));
  AOI21_X1  g444(.A(KEYINPUT86), .B1(new_n481), .B2(KEYINPUT20), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n629), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n484), .A2(KEYINPUT96), .A3(new_n485), .ZN(new_n633));
  OR2_X1    g447(.A1(new_n481), .A2(KEYINPUT20), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n632), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  AND2_X1   g449(.A1(new_n585), .A2(new_n530), .ZN(new_n636));
  AND3_X1   g450(.A1(new_n635), .A2(new_n616), .A3(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n611), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(KEYINPUT35), .B(G107), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G9));
  NAND2_X1  g455(.A1(new_n221), .A2(new_n227), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n232), .A2(KEYINPUT36), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(new_n246), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n645), .B1(new_n243), .B2(new_n244), .ZN(new_n646));
  AND2_X1   g460(.A1(new_n599), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n595), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT37), .B(G110), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G12));
  NOR2_X1   g464(.A1(new_n352), .A2(new_n353), .ZN(new_n651));
  AOI211_X1 g465(.A(KEYINPUT32), .B(new_n349), .C1(new_n350), .C2(new_n351), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n371), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n646), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n654), .A2(new_n615), .ZN(new_n655));
  AND3_X1   g469(.A1(new_n653), .A2(new_n608), .A3(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(G900), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n587), .B1(new_n591), .B2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n635), .A2(new_n636), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(KEYINPUT97), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT97), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n635), .A2(new_n662), .A3(new_n636), .A4(new_n659), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n656), .A2(new_n661), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G128), .ZN(G30));
  NAND2_X1  g479(.A1(new_n522), .A2(new_n523), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT38), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(new_n668));
  NOR3_X1   g482(.A1(new_n668), .A2(new_n490), .A3(new_n646), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n669), .A2(new_n612), .A3(new_n585), .ZN(new_n670));
  XOR2_X1   g484(.A(new_n658), .B(KEYINPUT39), .Z(new_n671));
  NAND2_X1  g485(.A1(new_n608), .A2(new_n671), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n670), .B1(KEYINPUT40), .B2(new_n672), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n332), .B1(new_n365), .B2(new_n364), .ZN(new_n674));
  AND3_X1   g488(.A1(new_n329), .A2(new_n330), .A3(new_n674), .ZN(new_n675));
  OAI21_X1  g489(.A(G472), .B1(new_n675), .B2(G902), .ZN(new_n676));
  AOI21_X1  g490(.A(KEYINPUT98), .B1(new_n355), .B2(new_n676), .ZN(new_n677));
  OAI211_X1 g491(.A(KEYINPUT98), .B(new_n676), .C1(new_n651), .C2(new_n652), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  OAI221_X1 g493(.A(new_n673), .B1(KEYINPUT40), .B2(new_n672), .C1(new_n677), .C2(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G143), .ZN(G45));
  NAND2_X1  g495(.A1(new_n612), .A2(new_n622), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n682), .A2(new_n658), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n656), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G146), .ZN(G48));
  OAI21_X1  g499(.A(new_n239), .B1(new_n600), .B2(new_n604), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n686), .A2(KEYINPUT99), .A3(G469), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT99), .ZN(new_n688));
  OAI21_X1  g502(.A(new_n688), .B1(new_n436), .B2(new_n373), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n607), .A2(new_n687), .A3(new_n443), .A4(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n372), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n692), .A2(new_n624), .ZN(new_n693));
  XOR2_X1   g507(.A(KEYINPUT41), .B(G113), .Z(new_n694));
  XNOR2_X1  g508(.A(new_n693), .B(new_n694), .ZN(G15));
  NOR2_X1   g509(.A1(new_n692), .A2(new_n638), .ZN(new_n696));
  XNOR2_X1  g510(.A(KEYINPUT100), .B(G116), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(G18));
  NOR2_X1   g512(.A1(new_n690), .A2(new_n615), .ZN(new_n699));
  AND4_X1   g513(.A1(new_n488), .A2(new_n646), .A3(new_n530), .A4(new_n593), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n699), .A2(new_n653), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(KEYINPUT101), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n488), .A2(new_n646), .A3(new_n530), .A4(new_n593), .ZN(new_n703));
  NOR3_X1   g517(.A1(new_n703), .A2(new_n690), .A3(new_n615), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT101), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n704), .A2(new_n705), .A3(new_n653), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n702), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(KEYINPUT102), .B(G119), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n707), .B(new_n708), .ZN(G21));
  NAND2_X1  g523(.A1(new_n368), .A2(new_n332), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT103), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n710), .A2(new_n351), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(new_n345), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n711), .B1(new_n710), .B2(new_n351), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n249), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n598), .A2(G472), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n715), .A2(new_n609), .A3(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(new_n614), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n490), .B1(new_n718), .B2(new_n523), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n612), .A2(new_n585), .A3(new_n719), .ZN(new_n720));
  AND2_X1   g534(.A1(new_n689), .A2(new_n687), .ZN(new_n721));
  INV_X1    g535(.A(new_n592), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n721), .A2(new_n443), .A3(new_n607), .A4(new_n722), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n717), .A2(new_n720), .A3(new_n723), .ZN(new_n724));
  XOR2_X1   g538(.A(KEYINPUT104), .B(G122), .Z(new_n725));
  XNOR2_X1  g539(.A(new_n724), .B(new_n725), .ZN(G24));
  AND3_X1   g540(.A1(new_n715), .A2(new_n716), .A3(new_n646), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n727), .A2(new_n683), .A3(new_n699), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G125), .ZN(G27));
  NAND3_X1  g543(.A1(new_n522), .A2(new_n489), .A3(new_n523), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT105), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n438), .A2(new_n731), .A3(new_n443), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n422), .B1(new_n606), .B2(new_n434), .ZN(new_n733));
  OAI21_X1  g547(.A(KEYINPUT105), .B1(new_n733), .B2(new_n442), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n730), .B1(new_n732), .B2(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n735), .A2(new_n683), .A3(new_n372), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT42), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n735), .A2(new_n683), .A3(new_n372), .A4(KEYINPUT42), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G131), .ZN(G33));
  NAND4_X1  g555(.A1(new_n661), .A2(new_n372), .A3(new_n735), .A4(new_n663), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G134), .ZN(G36));
  NAND3_X1  g557(.A1(new_n488), .A2(new_n530), .A3(new_n622), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(KEYINPUT43), .ZN(new_n745));
  NOR3_X1   g559(.A1(new_n745), .A2(new_n599), .A3(new_n654), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(KEYINPUT44), .ZN(new_n747));
  INV_X1    g561(.A(new_n607), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n421), .B(KEYINPUT45), .ZN(new_n749));
  OAI21_X1  g563(.A(G469), .B1(new_n749), .B2(G902), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n748), .B1(new_n750), .B2(KEYINPUT46), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n751), .B1(KEYINPUT46), .B2(new_n750), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n752), .A2(new_n443), .A3(new_n671), .ZN(new_n753));
  OR2_X1    g567(.A1(new_n753), .A2(KEYINPUT106), .ZN(new_n754));
  INV_X1    g568(.A(new_n730), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n753), .A2(KEYINPUT106), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n754), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n747), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(new_n266), .ZN(G39));
  AND3_X1   g573(.A1(new_n752), .A2(KEYINPUT47), .A3(new_n443), .ZN(new_n760));
  AOI21_X1  g574(.A(KEYINPUT47), .B1(new_n752), .B2(new_n443), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n683), .A2(new_n248), .A3(new_n755), .ZN(new_n763));
  OR3_X1    g577(.A1(new_n762), .A2(new_n653), .A3(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G140), .ZN(G42));
  INV_X1    g579(.A(new_n720), .ZN(new_n766));
  NOR3_X1   g580(.A1(new_n444), .A2(new_n646), .A3(new_n658), .ZN(new_n767));
  OAI211_X1 g581(.A(new_n766), .B(new_n767), .C1(new_n679), .C2(new_n677), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n664), .A2(new_n768), .A3(new_n684), .A4(new_n728), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(KEYINPUT52), .ZN(new_n770));
  INV_X1    g584(.A(new_n770), .ZN(new_n771));
  OAI211_X1 g585(.A(new_n372), .B(new_n691), .C1(new_n637), .C2(new_n623), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n724), .B1(new_n702), .B2(new_n706), .ZN(new_n773));
  AND3_X1   g587(.A1(new_n578), .A2(new_n239), .A3(new_n583), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n583), .B1(new_n578), .B2(new_n239), .ZN(new_n775));
  OAI21_X1  g589(.A(KEYINPUT108), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT108), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n582), .A2(new_n777), .A3(new_n584), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n779), .A2(new_n488), .A3(new_n530), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT109), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n779), .A2(new_n488), .A3(KEYINPUT109), .A4(new_n530), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n782), .A2(new_n682), .A3(new_n783), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n524), .A2(new_n722), .ZN(new_n785));
  AND4_X1   g599(.A1(new_n609), .A2(new_n599), .A3(new_n785), .A4(new_n608), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n595), .B1(new_n372), .B2(new_n647), .ZN(new_n788));
  AND3_X1   g602(.A1(new_n787), .A2(new_n788), .A3(KEYINPUT110), .ZN(new_n789));
  AOI21_X1  g603(.A(KEYINPUT110), .B1(new_n787), .B2(new_n788), .ZN(new_n790));
  OAI211_X1 g604(.A(new_n772), .B(new_n773), .C1(new_n789), .C2(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n646), .A2(new_n530), .A3(new_n659), .ZN(new_n792));
  NOR3_X1   g606(.A1(new_n792), .A2(new_n730), .A3(new_n779), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n793), .A2(new_n653), .A3(new_n608), .A4(new_n635), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n742), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n735), .A2(new_n727), .A3(new_n683), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n795), .A2(new_n740), .A3(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT111), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n791), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  OR3_X1    g613(.A1(new_n717), .A2(new_n720), .A3(new_n723), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n701), .A2(KEYINPUT101), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n705), .B1(new_n704), .B2(new_n653), .ZN(new_n802));
  OAI211_X1 g616(.A(new_n800), .B(new_n772), .C1(new_n801), .C2(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n787), .A2(new_n788), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT110), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n787), .A2(new_n788), .A3(KEYINPUT110), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n803), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n742), .A2(new_n796), .A3(new_n794), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n809), .B1(new_n738), .B2(new_n739), .ZN(new_n810));
  AOI21_X1  g624(.A(KEYINPUT111), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n771), .B1(new_n799), .B2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT114), .ZN(new_n813));
  XNOR2_X1  g627(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n812), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n798), .B1(new_n791), .B2(new_n797), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n806), .A2(new_n807), .ZN(new_n817));
  INV_X1    g631(.A(new_n803), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n810), .A2(KEYINPUT111), .A3(new_n817), .A4(new_n818), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n770), .B1(new_n816), .B2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(new_n814), .ZN(new_n821));
  OAI21_X1  g635(.A(KEYINPUT114), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n815), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n771), .A2(KEYINPUT53), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n808), .A2(new_n810), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n823), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n828), .A2(KEYINPUT54), .ZN(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n816), .A2(new_n819), .ZN(new_n831));
  XOR2_X1   g645(.A(new_n831), .B(KEYINPUT112), .Z(new_n832));
  AOI21_X1  g646(.A(KEYINPUT53), .B1(new_n832), .B2(new_n771), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n833), .B1(new_n820), .B2(new_n821), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT54), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n830), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(new_n587), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n745), .A2(new_n837), .A3(new_n717), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n838), .A2(new_n490), .A3(new_n668), .A4(new_n691), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT115), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(KEYINPUT50), .ZN(new_n841));
  XOR2_X1   g655(.A(new_n839), .B(new_n841), .Z(new_n842));
  OAI21_X1  g656(.A(new_n842), .B1(new_n840), .B2(KEYINPUT50), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n679), .A2(new_n677), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n690), .A2(new_n730), .ZN(new_n845));
  AND4_X1   g659(.A1(new_n609), .A2(new_n844), .A3(new_n587), .A4(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n612), .A2(new_n622), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  XNOR2_X1  g662(.A(new_n848), .B(KEYINPUT117), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n745), .A2(new_n837), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n850), .A2(new_n727), .A3(new_n845), .ZN(new_n851));
  XOR2_X1   g665(.A(new_n851), .B(KEYINPUT116), .Z(new_n852));
  INV_X1    g666(.A(new_n721), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n853), .A2(new_n748), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(new_n442), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n730), .B1(new_n762), .B2(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n852), .B1(new_n838), .B2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n843), .A2(new_n849), .A3(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT51), .ZN(new_n859));
  OR2_X1    g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n858), .A2(new_n859), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n838), .A2(new_n699), .ZN(new_n862));
  XOR2_X1   g676(.A(new_n862), .B(KEYINPUT118), .Z(new_n863));
  NAND3_X1  g677(.A1(new_n850), .A2(new_n372), .A3(new_n845), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n864), .B(KEYINPUT48), .ZN(new_n865));
  INV_X1    g679(.A(new_n682), .ZN(new_n866));
  AOI211_X1 g680(.A(new_n586), .B(G953), .C1(new_n846), .C2(new_n866), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n863), .A2(new_n865), .A3(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n860), .A2(new_n861), .A3(new_n868), .ZN(new_n869));
  OAI22_X1  g683(.A1(new_n836), .A2(new_n869), .B1(G952), .B2(G953), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n854), .B(KEYINPUT49), .ZN(new_n871));
  INV_X1    g685(.A(new_n668), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n609), .A2(new_n443), .A3(new_n489), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n872), .A2(new_n873), .A3(new_n744), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n871), .A2(new_n844), .A3(new_n874), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n875), .B(KEYINPUT107), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n870), .A2(new_n876), .ZN(G75));
  NOR2_X1   g691(.A1(new_n229), .A2(G952), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n878), .B(KEYINPUT121), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n239), .B1(new_n823), .B2(new_n827), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n880), .A2(new_n521), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n514), .A2(new_n517), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(new_n515), .ZN(new_n883));
  XOR2_X1   g697(.A(new_n883), .B(KEYINPUT55), .Z(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT56), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n879), .B1(new_n881), .B2(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT120), .ZN(new_n889));
  INV_X1    g703(.A(new_n520), .ZN(new_n890));
  AOI21_X1  g704(.A(KEYINPUT119), .B1(new_n880), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n826), .B1(new_n815), .B2(new_n822), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT119), .ZN(new_n893));
  NOR4_X1   g707(.A1(new_n892), .A2(new_n893), .A3(new_n239), .A4(new_n520), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n891), .A2(new_n894), .A3(KEYINPUT56), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n889), .B1(new_n895), .B2(new_n885), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n892), .A2(new_n239), .A3(new_n520), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n886), .B1(new_n897), .B2(KEYINPUT119), .ZN(new_n898));
  OAI211_X1 g712(.A(KEYINPUT120), .B(new_n884), .C1(new_n898), .C2(new_n894), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n888), .B1(new_n896), .B2(new_n899), .ZN(G51));
  NAND2_X1  g714(.A1(G469), .A2(G902), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n901), .B(KEYINPUT57), .Z(new_n902));
  NOR2_X1   g716(.A1(new_n892), .A2(new_n835), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n902), .B1(new_n829), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(new_n432), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n880), .A2(G469), .A3(new_n749), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n878), .B1(new_n905), .B2(new_n906), .ZN(G54));
  NAND3_X1  g721(.A1(new_n880), .A2(KEYINPUT58), .A3(G475), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n476), .A2(new_n480), .ZN(new_n909));
  OAI22_X1  g723(.A1(new_n908), .A2(new_n909), .B1(G952), .B2(new_n229), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n910), .B1(new_n908), .B2(new_n909), .ZN(G60));
  NAND2_X1  g725(.A1(G478), .A2(G902), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT59), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n620), .B1(new_n836), .B2(new_n913), .ZN(new_n914));
  OAI211_X1 g728(.A(new_n620), .B(new_n913), .C1(new_n829), .C2(new_n903), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(new_n879), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n914), .A2(new_n916), .ZN(G63));
  NAND2_X1  g731(.A1(G217), .A2(G902), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(KEYINPUT122), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(KEYINPUT60), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n828), .A2(new_n644), .A3(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(new_n920), .ZN(new_n922));
  OAI211_X1 g736(.A(new_n233), .B(new_n236), .C1(new_n892), .C2(new_n922), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n921), .A2(new_n923), .A3(new_n879), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g739(.A(G953), .B1(new_n590), .B2(new_n493), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n926), .B1(new_n808), .B2(G953), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n882), .B1(G898), .B2(new_n229), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n927), .B(new_n928), .ZN(G69));
  NAND2_X1  g743(.A1(new_n298), .A2(new_n316), .ZN(new_n930));
  OR2_X1    g744(.A1(new_n452), .A2(new_n453), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n930), .B(new_n931), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n932), .B1(G900), .B2(G953), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n754), .A2(new_n372), .A3(new_n766), .A4(new_n756), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n764), .A2(new_n742), .A3(new_n935), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n936), .A2(new_n758), .ZN(new_n937));
  AND3_X1   g751(.A1(new_n664), .A2(new_n684), .A3(new_n728), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n937), .A2(new_n740), .A3(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT125), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n939), .B(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n934), .B1(new_n941), .B2(new_n229), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT124), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n680), .A2(new_n938), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT62), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n944), .B(new_n945), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n672), .A2(new_n730), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n784), .A2(new_n372), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n764), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n949), .A2(new_n758), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n946), .A2(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT123), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n946), .A2(KEYINPUT123), .A3(new_n950), .ZN(new_n954));
  AND2_X1   g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  OAI211_X1 g769(.A(new_n943), .B(new_n932), .C1(new_n955), .C2(G953), .ZN(new_n956));
  AOI21_X1  g770(.A(G953), .B1(new_n953), .B2(new_n954), .ZN(new_n957));
  INV_X1    g771(.A(new_n932), .ZN(new_n958));
  OAI21_X1  g772(.A(KEYINPUT124), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n942), .B1(new_n956), .B2(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n229), .B1(G227), .B2(G900), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(KEYINPUT126), .ZN(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n960), .B(new_n963), .ZN(G72));
  NAND2_X1  g778(.A1(new_n941), .A2(new_n808), .ZN(new_n965));
  NAND2_X1  g779(.A1(G472), .A2(G902), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT63), .Z(new_n967));
  NAND2_X1  g781(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n317), .A2(new_n326), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n969), .A2(new_n324), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n878), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n329), .A2(new_n330), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n967), .B1(new_n972), .B2(new_n357), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n971), .B1(new_n834), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n969), .A2(new_n324), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n953), .A2(new_n808), .A3(new_n954), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n975), .B1(new_n976), .B2(new_n967), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n977), .B(KEYINPUT127), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n974), .A2(new_n978), .ZN(G57));
endmodule


