//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 1 1 0 0 1 1 1 0 0 0 1 1 0 0 1 1 0 0 0 1 1 0 0 0 1 1 0 0 1 1 1 1 0 0 0 0 0 1 0 0 1 0 0 1 0 1 1 1 0 1 1 1 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:56 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n449, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n535,
    new_n536, new_n537, new_n538, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n559, new_n560,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n621, new_n624, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n852, new_n853, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1201;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT64), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  INV_X1    g022(.A(G567), .ZN(new_n448));
  NOR2_X1   g023(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT65), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G2106), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n453), .A2(new_n457), .B1(new_n448), .B2(new_n454), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT66), .Z(G319));
  OR2_X1    g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G125), .ZN(new_n463));
  INV_X1    g038(.A(G113), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n462), .A2(G137), .A3(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n465), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G101), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(KEYINPUT67), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT67), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n469), .A2(new_n474), .A3(new_n471), .ZN(new_n475));
  AND3_X1   g050(.A1(new_n467), .A2(new_n473), .A3(new_n475), .ZN(G160));
  AOI21_X1  g051(.A(new_n468), .B1(new_n460), .B2(new_n461), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  OR2_X1    g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G112), .C2(new_n468), .ZN(new_n481));
  XOR2_X1   g056(.A(new_n481), .B(KEYINPUT69), .Z(new_n482));
  AND2_X1   g057(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n483));
  NOR2_X1   g058(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n468), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(KEYINPUT68), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT68), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(new_n468), .C1(new_n483), .C2(new_n484), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  AOI211_X1 g065(.A(new_n479), .B(new_n482), .C1(G136), .C2(new_n490), .ZN(G162));
  NAND2_X1  g066(.A1(KEYINPUT4), .A2(G138), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n492), .B1(new_n460), .B2(new_n461), .ZN(new_n493));
  AND2_X1   g068(.A1(G102), .A2(G2104), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n468), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(G126), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n496), .B1(new_n460), .B2(new_n461), .ZN(new_n497));
  AND2_X1   g072(.A1(G114), .A2(G2104), .ZN(new_n498));
  OAI21_X1  g073(.A(G2105), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  INV_X1    g075(.A(G138), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n500), .B1(new_n485), .B2(new_n501), .ZN(new_n502));
  AND3_X1   g077(.A1(new_n495), .A2(new_n499), .A3(new_n502), .ZN(G164));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(KEYINPUT6), .ZN(new_n505));
  XNOR2_X1  g080(.A(new_n505), .B(KEYINPUT70), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT71), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n507), .B1(new_n504), .B2(KEYINPUT6), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT6), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n509), .A2(KEYINPUT71), .A3(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n506), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G50), .ZN(new_n515));
  OR2_X1    g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n506), .A2(new_n511), .A3(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G88), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n518), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n522));
  OR2_X1    g097(.A1(new_n522), .A2(new_n504), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n515), .A2(new_n521), .A3(new_n523), .ZN(G303));
  INV_X1    g099(.A(G303), .ZN(G166));
  NAND2_X1  g100(.A1(new_n514), .A2(G51), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n520), .A2(G89), .ZN(new_n527));
  XNOR2_X1  g102(.A(KEYINPUT72), .B(KEYINPUT7), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n528), .B(new_n529), .ZN(new_n530));
  AND2_X1   g105(.A1(G63), .A2(G651), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n530), .B1(new_n518), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n526), .A2(new_n527), .A3(new_n532), .ZN(G286));
  INV_X1    g108(.A(G286), .ZN(G168));
  NAND2_X1  g109(.A1(new_n514), .A2(G52), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n520), .A2(G90), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n518), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n537), .A2(new_n504), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n535), .A2(new_n536), .A3(new_n538), .ZN(G301));
  INV_X1    g114(.A(G301), .ZN(G171));
  OR2_X1    g115(.A1(new_n505), .A2(KEYINPUT70), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n505), .A2(KEYINPUT70), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n541), .A2(new_n542), .B1(new_n508), .B2(new_n510), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n543), .A2(G43), .A3(G543), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n543), .A2(G81), .A3(new_n518), .ZN(new_n545));
  AND2_X1   g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(G68), .A2(G543), .ZN(new_n547));
  AND2_X1   g122(.A1(new_n516), .A2(new_n517), .ZN(new_n548));
  INV_X1    g123(.A(G56), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT73), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  OAI211_X1 g127(.A(KEYINPUT73), .B(new_n547), .C1(new_n548), .C2(new_n549), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n552), .A2(G651), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n546), .A2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  NAND4_X1  g132(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND4_X1  g135(.A1(G319), .A2(G483), .A3(G661), .A4(new_n560), .ZN(G188));
  NAND2_X1  g136(.A1(new_n519), .A2(KEYINPUT74), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT74), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n543), .A2(new_n563), .A3(new_n518), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n562), .A2(new_n564), .A3(G91), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n506), .A2(G53), .A3(G543), .A4(new_n511), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(KEYINPUT9), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT9), .ZN(new_n568));
  NAND4_X1  g143(.A1(new_n543), .A2(new_n568), .A3(G53), .A4(G543), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(G65), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT75), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n548), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n518), .A2(KEYINPUT75), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n571), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  AND2_X1   g150(.A1(G78), .A2(G543), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n565), .A2(new_n570), .A3(new_n577), .ZN(G299));
  OR2_X1    g153(.A1(new_n518), .A2(G74), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n514), .A2(G49), .B1(G651), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n562), .A2(new_n564), .A3(G87), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(G288));
  NAND2_X1  g157(.A1(G73), .A2(G543), .ZN(new_n583));
  INV_X1    g158(.A(G61), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n548), .B2(new_n584), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n514), .A2(G48), .B1(G651), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n562), .A2(new_n564), .A3(G86), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(G305));
  AOI22_X1  g163(.A1(new_n518), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n589));
  OR2_X1    g164(.A1(new_n589), .A2(new_n504), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n543), .A2(G85), .A3(new_n518), .ZN(new_n591));
  XOR2_X1   g166(.A(KEYINPUT76), .B(G47), .Z(new_n592));
  NAND3_X1  g167(.A1(new_n543), .A2(G543), .A3(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT77), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n591), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n594), .B1(new_n591), .B2(new_n593), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n590), .B1(new_n596), .B2(new_n597), .ZN(G290));
  NAND2_X1  g173(.A1(G301), .A2(G868), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n562), .A2(new_n564), .A3(G92), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT10), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g177(.A1(new_n562), .A2(new_n564), .A3(KEYINPUT10), .A4(G92), .ZN(new_n603));
  AND2_X1   g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n573), .A2(new_n574), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n605), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT78), .ZN(new_n607));
  OAI21_X1  g182(.A(G651), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(G79), .A2(G543), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n518), .B(new_n572), .ZN(new_n610));
  INV_X1    g185(.A(G66), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n609), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n612), .A2(KEYINPUT78), .ZN(new_n613));
  INV_X1    g188(.A(G54), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n543), .A2(G543), .ZN(new_n615));
  OAI22_X1  g190(.A1(new_n608), .A2(new_n613), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NOR2_X1   g191(.A1(new_n604), .A2(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n599), .B1(new_n617), .B2(G868), .ZN(G284));
  OAI21_X1  g193(.A(new_n599), .B1(new_n617), .B2(G868), .ZN(G321));
  NAND2_X1  g194(.A1(G286), .A2(G868), .ZN(new_n620));
  AND3_X1   g195(.A1(new_n565), .A2(new_n570), .A3(new_n577), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n621), .B2(G868), .ZN(G297));
  OAI21_X1  g197(.A(new_n620), .B1(new_n621), .B2(G868), .ZN(G280));
  INV_X1    g198(.A(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n617), .B1(new_n624), .B2(G860), .ZN(G148));
  NAND2_X1  g200(.A1(new_n617), .A2(new_n624), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT79), .ZN(new_n627));
  INV_X1    g202(.A(G868), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n556), .A2(new_n628), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(KEYINPUT80), .B(KEYINPUT11), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(G282));
  INV_X1    g208(.A(new_n631), .ZN(G323));
  NAND2_X1  g209(.A1(new_n462), .A2(new_n470), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT12), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT13), .ZN(new_n637));
  INV_X1    g212(.A(G2100), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n477), .A2(G123), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n468), .A2(G111), .ZN(new_n641));
  OAI21_X1  g216(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n642));
  INV_X1    g217(.A(G135), .ZN(new_n643));
  OAI221_X1 g218(.A(new_n640), .B1(new_n641), .B2(new_n642), .C1(new_n489), .C2(new_n643), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n644), .A2(G2096), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n637), .A2(new_n638), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n644), .A2(G2096), .ZN(new_n647));
  NAND4_X1  g222(.A1(new_n639), .A2(new_n645), .A3(new_n646), .A4(new_n647), .ZN(G156));
  XNOR2_X1  g223(.A(KEYINPUT15), .B(G2435), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT83), .B(G2438), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n649), .B(new_n650), .Z(new_n651));
  XNOR2_X1  g226(.A(G2427), .B(G2430), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n649), .B(new_n650), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n655), .A2(new_n652), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n654), .A2(KEYINPUT14), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT84), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(G1341), .ZN(new_n659));
  INV_X1    g234(.A(G1348), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2443), .B(G2446), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT82), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(G2451), .ZN(new_n664));
  XOR2_X1   g239(.A(KEYINPUT81), .B(KEYINPUT16), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(G2454), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n664), .B(new_n666), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n661), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n661), .A2(new_n667), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n668), .A2(G14), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT85), .ZN(G401));
  XOR2_X1   g246(.A(G2084), .B(G2090), .Z(new_n672));
  XNOR2_X1  g247(.A(G2067), .B(G2678), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(G2072), .B(G2078), .Z(new_n675));
  NOR2_X1   g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT18), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n675), .B(KEYINPUT17), .ZN(new_n678));
  INV_X1    g253(.A(new_n672), .ZN(new_n679));
  INV_X1    g254(.A(new_n673), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n678), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n679), .A2(new_n675), .A3(new_n680), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n682), .A2(new_n674), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n677), .B1(new_n681), .B2(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G2096), .B(G2100), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(G227));
  XOR2_X1   g261(.A(G1971), .B(G1976), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT19), .ZN(new_n688));
  XOR2_X1   g263(.A(G1956), .B(G2474), .Z(new_n689));
  XOR2_X1   g264(.A(G1961), .B(G1966), .Z(new_n690));
  AND2_X1   g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT20), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n689), .A2(new_n690), .ZN(new_n694));
  NOR3_X1   g269(.A1(new_n688), .A2(new_n691), .A3(new_n694), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n695), .B1(new_n688), .B2(new_n694), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(G1991), .B(G1996), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT86), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n699), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1981), .B(G1986), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(G229));
  INV_X1    g280(.A(G16), .ZN(new_n706));
  NOR2_X1   g281(.A1(G171), .A2(new_n706), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(G5), .B2(new_n706), .ZN(new_n708));
  INV_X1    g283(.A(G1961), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT97), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  NOR2_X1   g287(.A1(G29), .A2(G35), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(G162), .B2(G29), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT98), .B(KEYINPUT29), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n716), .A2(G2090), .ZN(new_n717));
  NOR2_X1   g292(.A1(G27), .A2(G29), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(G164), .B2(G29), .ZN(new_n719));
  AND2_X1   g294(.A1(new_n719), .A2(G2078), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n719), .A2(G2078), .ZN(new_n721));
  XOR2_X1   g296(.A(KEYINPUT31), .B(G11), .Z(new_n722));
  INV_X1    g297(.A(G28), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n723), .A2(KEYINPUT30), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT96), .ZN(new_n725));
  AOI21_X1  g300(.A(G29), .B1(new_n723), .B2(KEYINPUT30), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n722), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(G29), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n727), .B1(new_n644), .B2(new_n728), .ZN(new_n729));
  NOR3_X1   g304(.A1(new_n720), .A2(new_n721), .A3(new_n729), .ZN(new_n730));
  AND3_X1   g305(.A1(new_n712), .A2(new_n717), .A3(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(new_n477), .ZN(new_n732));
  INV_X1    g307(.A(G129), .ZN(new_n733));
  OAI21_X1  g308(.A(KEYINPUT94), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT94), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n477), .A2(new_n735), .A3(G129), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n486), .A2(G141), .A3(new_n488), .ZN(new_n738));
  NAND3_X1  g313(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT26), .ZN(new_n740));
  OR2_X1    g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n739), .A2(new_n740), .ZN(new_n742));
  AOI22_X1  g317(.A1(new_n741), .A2(new_n742), .B1(G105), .B2(new_n470), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n737), .A2(new_n738), .A3(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT95), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  MUX2_X1   g321(.A(G32), .B(new_n746), .S(G29), .Z(new_n747));
  XNOR2_X1  g322(.A(KEYINPUT27), .B(G1996), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n706), .A2(G20), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT23), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(new_n621), .B2(new_n706), .ZN(new_n752));
  INV_X1    g327(.A(G1956), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n716), .A2(G2090), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT99), .ZN(new_n756));
  NAND4_X1  g331(.A1(new_n731), .A2(new_n749), .A3(new_n754), .A4(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(G4), .A2(G16), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT89), .Z(new_n759));
  AOI21_X1  g334(.A(new_n504), .B1(new_n612), .B2(KEYINPUT78), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n606), .A2(new_n607), .ZN(new_n761));
  AOI22_X1  g336(.A1(new_n760), .A2(new_n761), .B1(G54), .B2(new_n514), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n602), .A2(new_n603), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n759), .B1(new_n764), .B2(new_n706), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(new_n660), .ZN(new_n766));
  NAND2_X1  g341(.A1(G168), .A2(G16), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G16), .B2(G21), .ZN(new_n768));
  INV_X1    g343(.A(G1966), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(KEYINPUT24), .ZN(new_n771));
  INV_X1    g346(.A(G34), .ZN(new_n772));
  AOI21_X1  g347(.A(G29), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(new_n771), .B2(new_n772), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G160), .B2(new_n728), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n775), .A2(G2084), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n728), .A2(G33), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT25), .Z(new_n779));
  AOI22_X1  g354(.A1(new_n462), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n780));
  INV_X1    g355(.A(G139), .ZN(new_n781));
  OAI221_X1 g356(.A(new_n779), .B1(new_n780), .B2(new_n468), .C1(new_n489), .C2(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(new_n782), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n777), .B1(new_n783), .B2(new_n728), .ZN(new_n784));
  XOR2_X1   g359(.A(KEYINPUT93), .B(G2072), .Z(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n775), .A2(G2084), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n770), .A2(new_n776), .A3(new_n786), .A4(new_n787), .ZN(new_n788));
  AOI22_X1  g363(.A1(new_n708), .A2(new_n709), .B1(new_n769), .B2(new_n768), .ZN(new_n789));
  NOR2_X1   g364(.A1(G16), .A2(G19), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(new_n556), .B2(G16), .ZN(new_n791));
  XOR2_X1   g366(.A(KEYINPUT90), .B(G1341), .Z(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT91), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n791), .B(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n789), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n728), .A2(G26), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT28), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n486), .A2(G140), .A3(new_n488), .ZN(new_n798));
  OAI21_X1  g373(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n799));
  INV_X1    g374(.A(G116), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n799), .B1(new_n800), .B2(G2105), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(G128), .B2(new_n477), .ZN(new_n802));
  AND3_X1   g377(.A1(new_n798), .A2(KEYINPUT92), .A3(new_n802), .ZN(new_n803));
  AOI21_X1  g378(.A(KEYINPUT92), .B1(new_n798), .B2(new_n802), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n797), .B1(new_n805), .B2(new_n728), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(G2067), .ZN(new_n807));
  OR4_X1    g382(.A1(new_n766), .A2(new_n788), .A3(new_n795), .A4(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n757), .A2(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  MUX2_X1   g385(.A(G24), .B(G290), .S(G16), .Z(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(G1986), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n728), .A2(G25), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n490), .A2(G131), .ZN(new_n814));
  OAI21_X1  g389(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n815));
  INV_X1    g390(.A(G107), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n815), .B1(new_n816), .B2(G2105), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(G119), .B2(new_n477), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n814), .A2(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n813), .B1(new_n820), .B2(new_n728), .ZN(new_n821));
  XOR2_X1   g396(.A(KEYINPUT35), .B(G1991), .Z(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n821), .B(new_n823), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n812), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n706), .A2(G6), .ZN(new_n826));
  AND2_X1   g401(.A1(new_n586), .A2(new_n587), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n826), .B1(new_n827), .B2(new_n706), .ZN(new_n828));
  XOR2_X1   g403(.A(KEYINPUT32), .B(G1981), .Z(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n706), .A2(G22), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n831), .B1(G166), .B2(new_n706), .ZN(new_n832));
  INV_X1    g407(.A(G1971), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  NOR2_X1   g409(.A1(G16), .A2(G23), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT87), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n836), .B1(G288), .B2(new_n706), .ZN(new_n837));
  XNOR2_X1  g412(.A(KEYINPUT33), .B(G1976), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n837), .A2(new_n838), .ZN(new_n840));
  AND4_X1   g415(.A1(new_n830), .A2(new_n834), .A3(new_n839), .A4(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n825), .B1(new_n842), .B2(KEYINPUT34), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT88), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n842), .A2(KEYINPUT34), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n847), .A2(KEYINPUT36), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT36), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n845), .A2(new_n849), .A3(new_n846), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n810), .B1(new_n848), .B2(new_n850), .ZN(G311));
  INV_X1    g426(.A(new_n850), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n849), .B1(new_n845), .B2(new_n846), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n809), .B1(new_n852), .B2(new_n853), .ZN(G150));
  NOR2_X1   g429(.A1(new_n764), .A2(new_n624), .ZN(new_n855));
  XNOR2_X1  g430(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n855), .B(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n554), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n544), .A2(new_n545), .ZN(new_n859));
  NAND2_X1  g434(.A1(G80), .A2(G543), .ZN(new_n860));
  INV_X1    g435(.A(G67), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n860), .B1(new_n548), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(G651), .ZN(new_n863));
  NAND4_X1  g438(.A1(new_n506), .A2(G55), .A3(G543), .A4(new_n511), .ZN(new_n864));
  NAND4_X1  g439(.A1(new_n506), .A2(G93), .A3(new_n511), .A4(new_n518), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  NOR3_X1   g441(.A1(new_n858), .A2(new_n859), .A3(new_n866), .ZN(new_n867));
  AND3_X1   g442(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n868), .B1(new_n546), .B2(new_n554), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n857), .B(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT39), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(KEYINPUT101), .ZN(new_n874));
  AOI21_X1  g449(.A(G860), .B1(new_n871), .B2(new_n872), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n866), .A2(G860), .ZN(new_n877));
  XOR2_X1   g452(.A(new_n877), .B(KEYINPUT37), .Z(new_n878));
  NAND2_X1  g453(.A1(new_n876), .A2(new_n878), .ZN(G145));
  XNOR2_X1  g454(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n880));
  XOR2_X1   g455(.A(G162), .B(G160), .Z(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(new_n644), .ZN(new_n882));
  NOR3_X1   g457(.A1(new_n803), .A2(new_n804), .A3(G164), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n495), .A2(new_n499), .A3(new_n502), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n798), .A2(new_n802), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT92), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n798), .A2(new_n802), .A3(KEYINPUT92), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n884), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n744), .B1(new_n883), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g465(.A(G164), .B1(new_n803), .B2(new_n804), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n887), .A2(new_n884), .A3(new_n888), .ZN(new_n892));
  AND3_X1   g467(.A1(new_n737), .A2(new_n738), .A3(new_n743), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n890), .A2(new_n782), .A3(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT103), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n895), .B(new_n896), .ZN(new_n897));
  AND3_X1   g472(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n893), .B1(new_n891), .B2(new_n892), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n745), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n890), .A2(KEYINPUT95), .A3(new_n894), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(KEYINPUT102), .B1(new_n902), .B2(new_n783), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT102), .ZN(new_n904));
  AOI211_X1 g479(.A(new_n904), .B(new_n782), .C1(new_n900), .C2(new_n901), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n897), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n490), .A2(G142), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n907), .B(KEYINPUT104), .ZN(new_n908));
  OR2_X1    g483(.A1(G106), .A2(G2105), .ZN(new_n909));
  OAI211_X1 g484(.A(new_n909), .B(G2104), .C1(G118), .C2(new_n468), .ZN(new_n910));
  INV_X1    g485(.A(G130), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n910), .B1(new_n732), .B2(new_n911), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n908), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n906), .A2(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n819), .B(new_n636), .ZN(new_n915));
  INV_X1    g490(.A(new_n913), .ZN(new_n916));
  OAI211_X1 g491(.A(new_n897), .B(new_n916), .C1(new_n903), .C2(new_n905), .ZN(new_n917));
  AND3_X1   g492(.A1(new_n914), .A2(new_n915), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n915), .B1(new_n914), .B2(new_n917), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n882), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n915), .ZN(new_n921));
  NOR3_X1   g496(.A1(new_n898), .A2(new_n899), .A3(new_n745), .ZN(new_n922));
  AOI21_X1  g497(.A(KEYINPUT95), .B1(new_n890), .B2(new_n894), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n783), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(new_n904), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n902), .A2(KEYINPUT102), .A3(new_n783), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n916), .B1(new_n927), .B2(new_n897), .ZN(new_n928));
  INV_X1    g503(.A(new_n917), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n921), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n882), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n914), .A2(new_n915), .A3(new_n917), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n920), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g509(.A(KEYINPUT105), .B(G37), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n880), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n935), .ZN(new_n937));
  INV_X1    g512(.A(new_n880), .ZN(new_n938));
  AOI211_X1 g513(.A(new_n937), .B(new_n938), .C1(new_n920), .C2(new_n933), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n936), .A2(new_n939), .ZN(G395));
  XNOR2_X1  g515(.A(new_n627), .B(new_n870), .ZN(new_n941));
  AND3_X1   g516(.A1(new_n762), .A2(new_n621), .A3(new_n763), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n621), .B1(new_n762), .B2(new_n763), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  OR2_X1    g520(.A1(new_n941), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT107), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT41), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n947), .B1(new_n944), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(KEYINPUT41), .B1(new_n942), .B2(new_n943), .ZN(new_n950));
  OAI21_X1  g525(.A(G299), .B1(new_n604), .B2(new_n616), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n762), .A2(new_n763), .A3(new_n621), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n951), .A2(new_n948), .A3(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(KEYINPUT107), .B1(new_n950), .B2(new_n953), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n941), .B1(new_n949), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(G290), .A2(new_n827), .ZN(new_n956));
  OAI211_X1 g531(.A(G305), .B(new_n590), .C1(new_n597), .C2(new_n596), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(G288), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(G303), .ZN(new_n960));
  NAND2_X1  g535(.A1(G166), .A2(G288), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n958), .A2(new_n962), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n956), .A2(new_n960), .A3(new_n957), .A4(new_n961), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n965), .A2(KEYINPUT108), .ZN(new_n966));
  XOR2_X1   g541(.A(new_n966), .B(KEYINPUT42), .Z(new_n967));
  AND3_X1   g542(.A1(new_n946), .A2(new_n955), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n967), .B1(new_n946), .B2(new_n955), .ZN(new_n969));
  OAI21_X1  g544(.A(G868), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n970), .B1(G868), .B2(new_n868), .ZN(G295));
  OAI21_X1  g546(.A(new_n970), .B1(G868), .B2(new_n868), .ZN(G331));
  INV_X1    g547(.A(KEYINPUT43), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT109), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n965), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n963), .A2(KEYINPUT109), .A3(new_n964), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n866), .B1(new_n858), .B2(new_n859), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n546), .A2(new_n554), .A3(new_n868), .ZN(new_n979));
  AND3_X1   g554(.A1(new_n978), .A2(new_n979), .A3(G301), .ZN(new_n980));
  AOI21_X1  g555(.A(G301), .B1(new_n978), .B2(new_n979), .ZN(new_n981));
  OAI21_X1  g556(.A(G286), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(G171), .B1(new_n867), .B2(new_n869), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n978), .A2(new_n979), .A3(G301), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n983), .A2(G168), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n982), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(new_n944), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n986), .B1(new_n953), .B2(new_n950), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n977), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(new_n935), .ZN(new_n991));
  INV_X1    g566(.A(new_n986), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n992), .B1(new_n954), .B2(new_n949), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n993), .A2(new_n965), .A3(new_n987), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT110), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n993), .A2(KEYINPUT110), .A3(new_n987), .A4(new_n965), .ZN(new_n997));
  AOI211_X1 g572(.A(new_n973), .B(new_n991), .C1(new_n996), .C2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n996), .A2(new_n997), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n993), .A2(new_n987), .ZN(new_n1000));
  AOI21_X1  g575(.A(G37), .B1(new_n1000), .B2(new_n977), .ZN(new_n1001));
  AOI21_X1  g576(.A(KEYINPUT43), .B1(new_n999), .B2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g577(.A(KEYINPUT44), .B1(new_n998), .B2(new_n1002), .ZN(new_n1003));
  AOI211_X1 g578(.A(KEYINPUT43), .B(new_n991), .C1(new_n996), .C2(new_n997), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n973), .B1(new_n999), .B2(new_n1001), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1003), .B1(new_n1006), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g582(.A(G1384), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n884), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT45), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n467), .A2(new_n473), .A3(G40), .A4(new_n475), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(G1996), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1015), .A2(new_n746), .ZN(new_n1016));
  XOR2_X1   g591(.A(new_n1016), .B(KEYINPUT111), .Z(new_n1017));
  XNOR2_X1  g592(.A(new_n805), .B(G2067), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1018), .B1(new_n1014), .B2(new_n893), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1017), .B1(new_n1013), .B2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n820), .A2(new_n822), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n819), .A2(new_n823), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1013), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1020), .A2(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g599(.A(G290), .B(G1986), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1024), .B1(new_n1013), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(G303), .A2(G8), .ZN(new_n1027));
  XOR2_X1   g602(.A(new_n1027), .B(KEYINPUT55), .Z(new_n1028));
  XNOR2_X1  g603(.A(new_n1028), .B(KEYINPUT114), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n884), .A2(KEYINPUT45), .A3(new_n1008), .ZN(new_n1030));
  XNOR2_X1  g605(.A(new_n1030), .B(KEYINPUT112), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1012), .B1(new_n1010), .B2(new_n1009), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(new_n833), .ZN(new_n1034));
  AND4_X1   g609(.A1(G40), .A2(new_n467), .A3(new_n473), .A4(new_n475), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1009), .A2(KEYINPUT50), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT50), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n884), .A2(new_n1037), .A3(new_n1008), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1035), .A2(new_n1036), .A3(new_n1038), .ZN(new_n1039));
  OR3_X1    g614(.A1(new_n1039), .A2(KEYINPUT113), .A3(G2090), .ZN(new_n1040));
  OAI21_X1  g615(.A(KEYINPUT113), .B1(new_n1039), .B2(G2090), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1034), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  AND2_X1   g617(.A1(new_n1042), .A2(G8), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1029), .A2(new_n1043), .ZN(new_n1044));
  OR2_X1    g619(.A1(G305), .A2(G1981), .ZN(new_n1045));
  INV_X1    g620(.A(G86), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n586), .B1(new_n1046), .B2(new_n519), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(G1981), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1045), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT49), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1045), .A2(KEYINPUT49), .A3(new_n1048), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1012), .A2(new_n1009), .ZN(new_n1053));
  INV_X1    g628(.A(G8), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1051), .A2(new_n1052), .A3(new_n1055), .ZN(new_n1056));
  AOI211_X1 g631(.A(new_n1054), .B(new_n1053), .C1(new_n959), .C2(G1976), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT52), .ZN(new_n1058));
  OR2_X1    g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1057), .B(new_n1058), .C1(G1976), .C2(new_n959), .ZN(new_n1060));
  AND3_X1   g635(.A1(new_n1056), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1034), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT115), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1063), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1038), .A2(new_n1063), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(new_n1035), .ZN(new_n1066));
  NOR3_X1   g641(.A1(new_n1064), .A2(new_n1066), .A3(G2090), .ZN(new_n1067));
  OAI21_X1  g642(.A(G8), .B1(new_n1062), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1028), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1044), .A2(new_n1061), .A3(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT120), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1035), .A2(new_n1011), .A3(new_n1030), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(new_n769), .ZN(new_n1074));
  XOR2_X1   g649(.A(KEYINPUT116), .B(G2084), .Z(new_n1075));
  NAND4_X1  g650(.A1(new_n1035), .A2(new_n1036), .A3(new_n1038), .A4(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT119), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1074), .A2(KEYINPUT119), .A3(new_n1076), .ZN(new_n1080));
  AOI21_X1  g655(.A(G286), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(KEYINPUT51), .A2(G8), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1072), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  AND3_X1   g658(.A1(new_n1074), .A2(KEYINPUT119), .A3(new_n1076), .ZN(new_n1084));
  AOI21_X1  g659(.A(KEYINPUT119), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1085));
  OAI21_X1  g660(.A(G168), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1086), .A2(KEYINPUT120), .A3(KEYINPUT51), .A4(G8), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1054), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1088));
  NOR2_X1   g663(.A1(G168), .A2(new_n1054), .ZN(new_n1089));
  OR3_X1    g664(.A1(new_n1088), .A2(KEYINPUT51), .A3(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1083), .A2(new_n1087), .A3(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1079), .A2(new_n1089), .A3(new_n1080), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(KEYINPUT62), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT118), .ZN(new_n1095));
  OR2_X1    g670(.A1(new_n1039), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1039), .A2(new_n1095), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1096), .A2(new_n709), .A3(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT53), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1099), .B1(new_n1033), .B2(G2078), .ZN(new_n1100));
  OR3_X1    g675(.A1(new_n1073), .A2(new_n1099), .A3(G2078), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1098), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(G171), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT62), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1091), .A2(new_n1105), .A3(new_n1092), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1094), .A2(new_n1104), .A3(new_n1106), .ZN(new_n1107));
  XNOR2_X1  g682(.A(new_n621), .B(KEYINPUT57), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n753), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1109));
  XNOR2_X1  g684(.A(KEYINPUT56), .B(G2072), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1031), .A2(new_n1032), .A3(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1108), .A2(new_n1109), .A3(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1096), .A2(new_n660), .A3(new_n1097), .ZN(new_n1113));
  INV_X1    g688(.A(G2067), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1053), .A2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n764), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1111), .A2(new_n1109), .ZN(new_n1117));
  XNOR2_X1  g692(.A(G299), .B(KEYINPUT57), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1119), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1112), .B1(new_n1116), .B2(new_n1120), .ZN(new_n1121));
  XNOR2_X1  g696(.A(KEYINPUT58), .B(G1341), .ZN(new_n1122));
  OAI22_X1  g697(.A1(new_n1033), .A2(G1996), .B1(new_n1053), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(new_n556), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(KEYINPUT59), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT59), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1123), .A2(new_n1126), .A3(new_n556), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1112), .A2(new_n1119), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT61), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  AND3_X1   g706(.A1(new_n1113), .A2(KEYINPUT60), .A3(new_n1115), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1132), .A2(new_n764), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1112), .A2(new_n1119), .A3(KEYINPUT61), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1128), .A2(new_n1131), .A3(new_n1133), .A4(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(KEYINPUT60), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1136));
  NOR3_X1   g711(.A1(new_n1132), .A2(new_n1136), .A3(new_n764), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1121), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT54), .ZN(new_n1139));
  XOR2_X1   g714(.A(KEYINPUT121), .B(G2078), .Z(new_n1140));
  NAND4_X1  g715(.A1(new_n1031), .A2(KEYINPUT53), .A3(new_n1032), .A4(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1098), .A2(new_n1100), .A3(new_n1141), .ZN(new_n1142));
  OAI211_X1 g717(.A(new_n1103), .B(new_n1139), .C1(G171), .C2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(KEYINPUT122), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT122), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1098), .A2(new_n1100), .A3(new_n1145), .A4(new_n1141), .ZN(new_n1146));
  AOI21_X1  g721(.A(G301), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1102), .A2(G301), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(KEYINPUT54), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1143), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1138), .A2(new_n1150), .A3(new_n1093), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1071), .B1(new_n1107), .B2(new_n1151), .ZN(new_n1152));
  NOR2_X1   g727(.A1(G288), .A2(G1976), .ZN(new_n1153));
  AND2_X1   g728(.A1(new_n1056), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1045), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1055), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1088), .A2(G168), .ZN(new_n1157));
  XNOR2_X1  g732(.A(new_n1157), .B(KEYINPUT117), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1061), .A2(new_n1158), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1043), .A2(new_n1028), .ZN(new_n1160));
  OAI21_X1  g735(.A(KEYINPUT63), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT63), .ZN(new_n1162));
  AND2_X1   g737(.A1(new_n1158), .A2(new_n1162), .ZN(new_n1163));
  AOI22_X1  g738(.A1(new_n1163), .A2(new_n1070), .B1(new_n1043), .B2(new_n1029), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1061), .ZN(new_n1165));
  OAI211_X1 g740(.A(new_n1156), .B(new_n1161), .C1(new_n1164), .C2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1026), .B1(new_n1152), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1018), .A2(new_n893), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1168), .A2(new_n1013), .ZN(new_n1169));
  XOR2_X1   g744(.A(new_n1169), .B(KEYINPUT125), .Z(new_n1170));
  NAND3_X1  g745(.A1(new_n1015), .A2(KEYINPUT124), .A3(KEYINPUT46), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT124), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT46), .ZN(new_n1173));
  OAI211_X1 g748(.A(new_n1013), .B(new_n1014), .C1(new_n1172), .C2(new_n1173), .ZN(new_n1174));
  AOI22_X1  g749(.A1(new_n1171), .A2(new_n1174), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1170), .A2(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT126), .ZN(new_n1177));
  XNOR2_X1  g752(.A(new_n1176), .B(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT47), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  XNOR2_X1  g755(.A(new_n1176), .B(KEYINPUT126), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1181), .A2(KEYINPUT47), .ZN(new_n1182));
  XOR2_X1   g757(.A(new_n1022), .B(KEYINPUT123), .Z(new_n1183));
  AOI22_X1  g758(.A1(new_n1020), .A2(new_n1183), .B1(new_n1114), .B2(new_n805), .ZN(new_n1184));
  OR3_X1    g759(.A1(new_n1184), .A2(new_n1012), .A3(new_n1011), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT127), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1024), .A2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1020), .A2(KEYINPUT127), .A3(new_n1023), .ZN(new_n1188));
  NOR4_X1   g763(.A1(G290), .A2(G1986), .A3(new_n1012), .A4(new_n1011), .ZN(new_n1189));
  XOR2_X1   g764(.A(new_n1189), .B(KEYINPUT48), .Z(new_n1190));
  NAND3_X1  g765(.A1(new_n1187), .A2(new_n1188), .A3(new_n1190), .ZN(new_n1191));
  AND4_X1   g766(.A1(new_n1180), .A2(new_n1182), .A3(new_n1185), .A4(new_n1191), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1167), .A2(new_n1192), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g768(.A(G319), .ZN(new_n1195));
  NOR2_X1   g769(.A1(new_n1195), .A2(G227), .ZN(new_n1196));
  AND3_X1   g770(.A1(new_n670), .A2(new_n704), .A3(new_n1196), .ZN(new_n1197));
  OAI21_X1  g771(.A(new_n1197), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1198));
  AOI21_X1  g772(.A(new_n937), .B1(new_n920), .B2(new_n933), .ZN(new_n1199));
  NOR2_X1   g773(.A1(new_n1198), .A2(new_n1199), .ZN(G308));
  NAND2_X1  g774(.A1(new_n934), .A2(new_n935), .ZN(new_n1201));
  OAI211_X1 g775(.A(new_n1201), .B(new_n1197), .C1(new_n1005), .C2(new_n1004), .ZN(G225));
endmodule


