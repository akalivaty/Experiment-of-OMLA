//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 1 1 0 0 1 0 0 1 1 0 0 0 0 1 1 1 1 1 0 1 0 0 0 1 0 1 1 0 1 1 0 0 1 1 1 0 1 1 0 0 1 0 1 0 1 1 1 0 1 1 1 1 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n800, new_n801, new_n802, new_n803, new_n804, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n818, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n843, new_n844, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n897,
    new_n898, new_n900, new_n901, new_n903, new_n904, new_n905, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n979, new_n980, new_n981;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT93), .ZN(new_n203));
  XNOR2_X1  g002(.A(G15gat), .B(G43gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n204), .B(KEYINPUT75), .ZN(new_n205));
  XOR2_X1   g004(.A(G71gat), .B(G99gat), .Z(new_n206));
  XNOR2_X1  g005(.A(new_n205), .B(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(G227gat), .A2(G233gat), .ZN(new_n209));
  XOR2_X1   g008(.A(new_n209), .B(KEYINPUT64), .Z(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212));
  AND2_X1   g011(.A1(KEYINPUT68), .A2(KEYINPUT24), .ZN(new_n213));
  NOR2_X1   g012(.A1(KEYINPUT68), .A2(KEYINPUT24), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT69), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OAI211_X1 g016(.A(KEYINPUT69), .B(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n218));
  INV_X1    g017(.A(G183gat), .ZN(new_n219));
  INV_X1    g018(.A(G190gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g020(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n222));
  AND2_X1   g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n217), .A2(new_n218), .A3(new_n223), .ZN(new_n224));
  NOR2_X1   g023(.A1(G169gat), .A2(G176gat), .ZN(new_n225));
  OAI21_X1  g024(.A(KEYINPUT23), .B1(new_n225), .B2(KEYINPUT67), .ZN(new_n226));
  NAND2_X1  g025(.A1(G169gat), .A2(G176gat), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT67), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT23), .ZN(new_n229));
  OAI211_X1 g028(.A(new_n228), .B(new_n229), .C1(G169gat), .C2(G176gat), .ZN(new_n230));
  AND4_X1   g029(.A1(KEYINPUT25), .A2(new_n226), .A3(new_n227), .A4(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n224), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n226), .A2(new_n227), .A3(new_n230), .ZN(new_n233));
  AOI21_X1  g032(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT66), .ZN(new_n235));
  OAI22_X1  g034(.A1(new_n234), .A2(new_n235), .B1(new_n222), .B2(KEYINPUT65), .ZN(new_n236));
  AND2_X1   g035(.A1(new_n234), .A2(new_n235), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NOR2_X1   g037(.A1(G183gat), .A2(G190gat), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n239), .B1(KEYINPUT65), .B2(new_n222), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n233), .B1(new_n238), .B2(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n232), .B1(new_n241), .B2(KEYINPUT25), .ZN(new_n242));
  INV_X1    g041(.A(new_n212), .ZN(new_n243));
  NOR3_X1   g042(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT73), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n244), .B(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n227), .ZN(new_n247));
  INV_X1    g046(.A(new_n225), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n247), .B1(new_n248), .B2(KEYINPUT26), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n243), .B1(new_n246), .B2(new_n249), .ZN(new_n250));
  XOR2_X1   g049(.A(KEYINPUT72), .B(KEYINPUT28), .Z(new_n251));
  INV_X1    g050(.A(KEYINPUT70), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n252), .B1(new_n219), .B2(KEYINPUT27), .ZN(new_n253));
  AOI21_X1  g052(.A(G190gat), .B1(new_n219), .B2(KEYINPUT27), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT27), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n255), .A2(KEYINPUT70), .A3(G183gat), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n253), .A2(new_n254), .A3(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT71), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n253), .A2(new_n254), .A3(KEYINPUT71), .A4(new_n256), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n251), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n219), .A2(KEYINPUT27), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n263), .A2(KEYINPUT28), .A3(new_n254), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n250), .B1(new_n261), .B2(new_n265), .ZN(new_n266));
  AND2_X1   g065(.A1(new_n242), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(G113gat), .B(G120gat), .ZN(new_n268));
  INV_X1    g067(.A(G127gat), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n269), .A2(G134gat), .ZN(new_n270));
  INV_X1    g069(.A(G134gat), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n271), .A2(G127gat), .ZN(new_n272));
  OAI22_X1  g071(.A1(new_n268), .A2(KEYINPUT1), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(G120gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(G113gat), .ZN(new_n275));
  INV_X1    g074(.A(G113gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(G120gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G127gat), .B(G134gat), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT1), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n278), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  AND2_X1   g080(.A1(new_n273), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n267), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n242), .A2(new_n266), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n273), .A2(new_n281), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n211), .B1(new_n283), .B2(new_n286), .ZN(new_n287));
  OAI211_X1 g086(.A(KEYINPUT74), .B(new_n208), .C1(new_n287), .C2(KEYINPUT33), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT32), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  AND2_X1   g089(.A1(new_n208), .A2(KEYINPUT33), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n288), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n283), .A2(new_n211), .A3(new_n286), .ZN(new_n293));
  XOR2_X1   g092(.A(new_n293), .B(KEYINPUT34), .Z(new_n294));
  INV_X1    g093(.A(KEYINPUT74), .ZN(new_n295));
  OAI211_X1 g094(.A(new_n295), .B(new_n208), .C1(new_n287), .C2(KEYINPUT33), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n283), .A2(new_n286), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(new_n210), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(KEYINPUT32), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  AND3_X1   g099(.A1(new_n292), .A2(new_n294), .A3(new_n300), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n294), .B1(new_n300), .B2(new_n292), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n203), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n292), .A2(new_n300), .ZN(new_n304));
  INV_X1    g103(.A(new_n294), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n292), .A2(new_n294), .A3(new_n300), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n306), .A2(KEYINPUT93), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n303), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(G225gat), .A2(G233gat), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(G148gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(G141gat), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(KEYINPUT81), .B(G141gat), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n314), .B1(new_n315), .B2(G148gat), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT2), .ZN(new_n317));
  INV_X1    g116(.A(G155gat), .ZN(new_n318));
  INV_X1    g117(.A(G162gat), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n317), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(G155gat), .A2(G162gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT80), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n324), .A2(new_n318), .A3(new_n319), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n321), .A2(KEYINPUT79), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT79), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n327), .A2(G155gat), .A3(G162gat), .ZN(new_n328));
  OAI21_X1  g127(.A(KEYINPUT80), .B1(G155gat), .B2(G162gat), .ZN(new_n329));
  NAND4_X1  g128(.A1(new_n325), .A2(new_n326), .A3(new_n328), .A4(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(G141gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(G148gat), .ZN(new_n332));
  AOI22_X1  g131(.A1(new_n313), .A2(new_n332), .B1(KEYINPUT2), .B2(new_n321), .ZN(new_n333));
  OAI22_X1  g132(.A1(new_n316), .A2(new_n323), .B1(new_n330), .B2(new_n333), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n334), .A2(new_n285), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n313), .A2(new_n332), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n321), .A2(KEYINPUT2), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  AND2_X1   g137(.A1(new_n325), .A2(new_n329), .ZN(new_n339));
  AND2_X1   g138(.A1(new_n326), .A2(new_n328), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n331), .A2(KEYINPUT81), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT81), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(G141gat), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n342), .A2(new_n344), .A3(G148gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(new_n313), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(new_n322), .ZN(new_n347));
  AOI22_X1  g146(.A1(new_n341), .A2(new_n347), .B1(new_n281), .B2(new_n273), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n311), .B1(new_n335), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(KEYINPUT5), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT3), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n341), .A2(new_n347), .A3(new_n351), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n330), .A2(new_n333), .ZN(new_n353));
  AOI22_X1  g152(.A1(new_n345), .A2(new_n313), .B1(new_n321), .B2(new_n320), .ZN(new_n354));
  OAI21_X1  g153(.A(KEYINPUT3), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n352), .A2(new_n355), .A3(new_n285), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT4), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n357), .B1(new_n334), .B2(new_n285), .ZN(new_n358));
  NAND4_X1  g157(.A1(new_n282), .A2(KEYINPUT4), .A3(new_n347), .A4(new_n341), .ZN(new_n359));
  NAND4_X1  g158(.A1(new_n356), .A2(new_n310), .A3(new_n358), .A4(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n350), .A2(new_n360), .ZN(new_n361));
  AND2_X1   g160(.A1(new_n359), .A2(new_n358), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n362), .A2(KEYINPUT5), .A3(new_n310), .A4(new_n356), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  XNOR2_X1  g163(.A(G1gat), .B(G29gat), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n365), .B(KEYINPUT0), .ZN(new_n366));
  XNOR2_X1  g165(.A(G57gat), .B(G85gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n366), .B(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  AOI21_X1  g168(.A(KEYINPUT6), .B1(new_n364), .B2(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n361), .A2(new_n363), .A3(new_n368), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT6), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n372), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(G226gat), .A2(G233gat), .ZN(new_n377));
  XOR2_X1   g176(.A(new_n377), .B(KEYINPUT76), .Z(new_n378));
  AND2_X1   g177(.A1(new_n244), .A2(new_n245), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n244), .A2(new_n245), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n249), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(new_n212), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n259), .A2(new_n260), .ZN(new_n383));
  INV_X1    g182(.A(new_n251), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n382), .B1(new_n385), .B2(new_n264), .ZN(new_n386));
  OAI21_X1  g185(.A(KEYINPUT66), .B1(new_n243), .B2(KEYINPUT24), .ZN(new_n387));
  OR2_X1    g186(.A1(new_n222), .A2(KEYINPUT65), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n234), .A2(new_n235), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n387), .A2(new_n388), .A3(new_n240), .A4(new_n389), .ZN(new_n390));
  AND2_X1   g189(.A1(new_n226), .A2(new_n227), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n390), .A2(new_n230), .A3(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT25), .ZN(new_n393));
  AOI22_X1  g192(.A1(new_n392), .A2(new_n393), .B1(new_n224), .B2(new_n231), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n378), .B1(new_n386), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(G211gat), .A2(G218gat), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT22), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NOR2_X1   g197(.A1(G197gat), .A2(G204gat), .ZN(new_n399));
  AND2_X1   g198(.A1(G197gat), .A2(G204gat), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n398), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  XOR2_X1   g200(.A(G211gat), .B(G218gat), .Z(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(G211gat), .B(G218gat), .ZN(new_n404));
  XNOR2_X1  g203(.A(G197gat), .B(G204gat), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n404), .A2(new_n405), .A3(new_n398), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n403), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n395), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT77), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT29), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n411), .B1(new_n386), .B2(new_n394), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n410), .B1(new_n412), .B2(new_n377), .ZN(new_n413));
  AOI21_X1  g212(.A(KEYINPUT29), .B1(new_n242), .B2(new_n266), .ZN(new_n414));
  INV_X1    g213(.A(new_n377), .ZN(new_n415));
  NOR3_X1   g214(.A1(new_n414), .A2(KEYINPUT77), .A3(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n409), .B1(new_n413), .B2(new_n416), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n415), .B1(new_n386), .B2(new_n394), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n418), .B1(new_n414), .B2(new_n378), .ZN(new_n419));
  INV_X1    g218(.A(new_n407), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  XOR2_X1   g220(.A(G8gat), .B(G36gat), .Z(new_n422));
  XNOR2_X1  g221(.A(new_n422), .B(KEYINPUT78), .ZN(new_n423));
  XNOR2_X1  g222(.A(G64gat), .B(G92gat), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n423), .B(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n417), .A2(new_n421), .A3(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT30), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n417), .A2(KEYINPUT30), .A3(new_n421), .A4(new_n426), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n417), .A2(new_n421), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(new_n425), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n376), .A2(new_n429), .A3(new_n430), .A4(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT92), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n433), .B(new_n434), .ZN(new_n435));
  XNOR2_X1  g234(.A(G78gat), .B(G106gat), .ZN(new_n436));
  XNOR2_X1  g235(.A(KEYINPUT31), .B(G50gat), .ZN(new_n437));
  XOR2_X1   g236(.A(new_n436), .B(new_n437), .Z(new_n438));
  AOI21_X1  g237(.A(new_n407), .B1(new_n352), .B2(new_n411), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n401), .A2(new_n402), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n404), .B1(new_n398), .B2(new_n405), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n411), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  AOI22_X1  g241(.A1(new_n442), .A2(new_n351), .B1(new_n347), .B2(new_n341), .ZN(new_n443));
  OAI21_X1  g242(.A(KEYINPUT83), .B1(new_n439), .B2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT83), .ZN(new_n445));
  AOI21_X1  g244(.A(KEYINPUT29), .B1(new_n403), .B2(new_n406), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n334), .B1(new_n446), .B2(KEYINPUT3), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n353), .A2(new_n354), .ZN(new_n448));
  AOI21_X1  g247(.A(KEYINPUT29), .B1(new_n448), .B2(new_n351), .ZN(new_n449));
  OAI211_X1 g248(.A(new_n445), .B(new_n447), .C1(new_n449), .C2(new_n407), .ZN(new_n450));
  NAND2_X1  g249(.A1(G228gat), .A2(G233gat), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n444), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n451), .ZN(new_n453));
  OAI211_X1 g252(.A(KEYINPUT83), .B(new_n453), .C1(new_n439), .C2(new_n443), .ZN(new_n454));
  AND3_X1   g253(.A1(new_n452), .A2(new_n454), .A3(G22gat), .ZN(new_n455));
  AOI21_X1  g254(.A(G22gat), .B1(new_n452), .B2(new_n454), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n438), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT84), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n452), .A2(new_n454), .ZN(new_n460));
  INV_X1    g259(.A(G22gat), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT85), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n452), .A2(new_n454), .A3(G22gat), .ZN(new_n465));
  INV_X1    g264(.A(new_n438), .ZN(new_n466));
  AND2_X1   g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n456), .A2(KEYINPUT85), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n464), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  OAI211_X1 g268(.A(KEYINPUT84), .B(new_n438), .C1(new_n455), .C2(new_n456), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n459), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(KEYINPUT86), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT86), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n459), .A2(new_n469), .A3(new_n473), .A4(new_n470), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  AND4_X1   g274(.A1(new_n202), .A2(new_n309), .A3(new_n435), .A4(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n371), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n364), .A2(new_n369), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(new_n373), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n477), .B1(new_n479), .B2(KEYINPUT82), .ZN(new_n480));
  AOI211_X1 g279(.A(KEYINPUT82), .B(KEYINPUT6), .C1(new_n364), .C2(new_n369), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n374), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n429), .A2(new_n430), .A3(new_n432), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n306), .A2(new_n307), .ZN(new_n486));
  AOI21_X1  g285(.A(KEYINPUT85), .B1(new_n460), .B2(new_n461), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n465), .A2(new_n466), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AOI22_X1  g288(.A1(new_n489), .A2(new_n468), .B1(new_n457), .B2(new_n458), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n473), .B1(new_n490), .B2(new_n470), .ZN(new_n491));
  AND4_X1   g290(.A1(new_n473), .A2(new_n459), .A3(new_n469), .A4(new_n470), .ZN(new_n492));
  OAI211_X1 g291(.A(new_n485), .B(new_n486), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(KEYINPUT35), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(KEYINPUT94), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT94), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n493), .A2(new_n496), .A3(KEYINPUT35), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n476), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT87), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT82), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n371), .B1(new_n370), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n375), .B1(new_n501), .B2(new_n481), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n426), .B1(new_n417), .B2(new_n421), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n503), .B1(new_n428), .B2(new_n427), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n502), .A2(new_n504), .A3(new_n430), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n472), .A2(new_n505), .A3(new_n474), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT36), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n508), .B1(new_n301), .B2(new_n302), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n306), .A2(KEYINPUT36), .A3(new_n307), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n499), .B1(new_n507), .B2(new_n511), .ZN(new_n512));
  AND2_X1   g311(.A1(new_n509), .A2(new_n510), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n513), .A2(KEYINPUT87), .A3(new_n506), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n372), .A2(new_n427), .A3(new_n375), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT38), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n426), .B1(new_n431), .B2(KEYINPUT37), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT89), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT37), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n377), .B1(new_n242), .B2(new_n266), .ZN(new_n520));
  INV_X1    g319(.A(new_n378), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n520), .B1(new_n412), .B2(new_n521), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n519), .B1(new_n522), .B2(new_n407), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n412), .A2(new_n410), .A3(new_n377), .ZN(new_n524));
  OAI21_X1  g323(.A(KEYINPUT77), .B1(new_n414), .B2(new_n415), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n408), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n518), .B1(new_n523), .B2(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(KEYINPUT37), .B1(new_n419), .B2(new_n420), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n417), .A2(KEYINPUT89), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n516), .B1(new_n517), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT91), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n515), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NOR3_X1   g332(.A1(new_n523), .A2(new_n526), .A3(new_n518), .ZN(new_n534));
  AOI21_X1  g333(.A(KEYINPUT89), .B1(new_n417), .B2(new_n528), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n421), .ZN(new_n537));
  OAI21_X1  g336(.A(KEYINPUT37), .B1(new_n537), .B2(new_n526), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(new_n425), .ZN(new_n539));
  OAI21_X1  g338(.A(KEYINPUT38), .B1(new_n536), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(KEYINPUT91), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n425), .A2(new_n516), .ZN(new_n542));
  OAI211_X1 g341(.A(new_n420), .B(new_n395), .C1(new_n413), .C2(new_n416), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n519), .B1(new_n419), .B2(new_n407), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n530), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT90), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  OAI211_X1 g347(.A(KEYINPUT90), .B(new_n545), .C1(new_n534), .C2(new_n535), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n533), .A2(new_n541), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n362), .A2(new_n356), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(new_n311), .ZN(new_n553));
  OR3_X1    g352(.A1(new_n335), .A2(new_n348), .A3(new_n311), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n553), .A2(KEYINPUT39), .A3(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(KEYINPUT88), .B(KEYINPUT39), .ZN(new_n556));
  OAI211_X1 g355(.A(new_n555), .B(new_n369), .C1(new_n553), .C2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT40), .ZN(new_n558));
  AND2_X1   g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n557), .A2(new_n558), .ZN(new_n560));
  NOR3_X1   g359(.A1(new_n559), .A2(new_n560), .A3(new_n477), .ZN(new_n561));
  AOI22_X1  g360(.A1(new_n472), .A2(new_n474), .B1(new_n561), .B2(new_n484), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n551), .A2(new_n562), .ZN(new_n563));
  AND3_X1   g362(.A1(new_n512), .A2(new_n514), .A3(new_n563), .ZN(new_n564));
  OR2_X1    g363(.A1(new_n498), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(G15gat), .B(G22gat), .ZN(new_n566));
  OR2_X1    g365(.A1(new_n566), .A2(G1gat), .ZN(new_n567));
  AOI21_X1  g366(.A(G8gat), .B1(new_n567), .B2(KEYINPUT96), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT16), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n566), .B1(new_n569), .B2(G1gat), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n568), .B(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(G29gat), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n574), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n575));
  AND2_X1   g374(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n576));
  NOR2_X1   g375(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n575), .B1(new_n578), .B2(G36gat), .ZN(new_n579));
  OR2_X1    g378(.A1(new_n579), .A2(KEYINPUT15), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(KEYINPUT15), .ZN(new_n581));
  XNOR2_X1  g380(.A(G43gat), .B(G50gat), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n583), .B1(new_n581), .B2(new_n582), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n573), .A2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(KEYINPUT98), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n584), .B(KEYINPUT17), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n572), .B(KEYINPUT97), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AND2_X1   g388(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(G229gat), .A2(G233gat), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n590), .A2(KEYINPUT18), .A3(new_n591), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n586), .B1(new_n573), .B2(new_n584), .ZN(new_n593));
  XOR2_X1   g392(.A(new_n591), .B(KEYINPUT13), .Z(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n586), .A2(new_n591), .A3(new_n589), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT18), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n592), .A2(new_n595), .A3(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(G113gat), .B(G141gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(G197gat), .ZN(new_n601));
  XOR2_X1   g400(.A(KEYINPUT11), .B(G169gat), .Z(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(KEYINPUT95), .B(KEYINPUT12), .ZN(new_n604));
  XOR2_X1   g403(.A(new_n603), .B(new_n604), .Z(new_n605));
  NAND2_X1  g404(.A1(new_n599), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n605), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n592), .A2(new_n607), .A3(new_n595), .A4(new_n598), .ZN(new_n608));
  AND2_X1   g407(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(G71gat), .B(G78gat), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT99), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(G57gat), .B(G64gat), .ZN(new_n615));
  NOR3_X1   g414(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n611), .A2(new_n612), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  OAI211_X1 g417(.A(new_n612), .B(new_n611), .C1(new_n615), .C2(new_n614), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n620), .A2(KEYINPUT21), .ZN(new_n621));
  NAND2_X1  g420(.A1(G231gat), .A2(G233gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(new_n269), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n573), .B1(KEYINPUT21), .B2(new_n620), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(G183gat), .B(G211gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(KEYINPUT100), .ZN(new_n628));
  XNOR2_X1  g427(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(new_n318), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n628), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n626), .B(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(G85gat), .A2(G92gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(KEYINPUT7), .ZN(new_n634));
  NAND2_X1  g433(.A1(G99gat), .A2(G106gat), .ZN(new_n635));
  INV_X1    g434(.A(G85gat), .ZN(new_n636));
  INV_X1    g435(.A(G92gat), .ZN(new_n637));
  AOI22_X1  g436(.A1(KEYINPUT8), .A2(new_n635), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  AND2_X1   g437(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(G99gat), .B(G106gat), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(KEYINPUT101), .ZN(new_n642));
  OR2_X1    g441(.A1(new_n639), .A2(new_n640), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n587), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(G190gat), .B(G218gat), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT41), .ZN(new_n648));
  NAND2_X1  g447(.A1(G232gat), .A2(G233gat), .ZN(new_n649));
  OAI22_X1  g448(.A1(new_n647), .A2(KEYINPUT102), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n644), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n650), .B1(new_n651), .B2(new_n584), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n645), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n647), .A2(KEYINPUT102), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT103), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n653), .B(new_n655), .ZN(new_n656));
  XOR2_X1   g455(.A(G134gat), .B(G162gat), .Z(new_n657));
  NAND2_X1  g456(.A1(new_n649), .A2(new_n648), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(new_n659));
  OR2_X1    g458(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n656), .A2(new_n659), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n632), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT108), .ZN(new_n664));
  INV_X1    g463(.A(G230gat), .ZN(new_n665));
  INV_X1    g464(.A(G233gat), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n620), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n644), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g468(.A(new_n640), .B(KEYINPUT104), .Z(new_n670));
  NOR2_X1   g469(.A1(new_n670), .A2(new_n639), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT105), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NOR3_X1   g472(.A1(new_n670), .A2(KEYINPUT105), .A3(new_n639), .ZN(new_n674));
  OAI211_X1 g473(.A(new_n642), .B(new_n620), .C1(new_n673), .C2(new_n674), .ZN(new_n675));
  XOR2_X1   g474(.A(KEYINPUT106), .B(KEYINPUT10), .Z(new_n676));
  NAND3_X1  g475(.A1(new_n669), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n651), .A2(KEYINPUT10), .A3(new_n620), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n667), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  AOI211_X1 g478(.A(new_n665), .B(new_n666), .C1(new_n669), .C2(new_n675), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n664), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  XOR2_X1   g480(.A(G120gat), .B(G148gat), .Z(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(KEYINPUT107), .ZN(new_n683));
  XNOR2_X1  g482(.A(G176gat), .B(G204gat), .ZN(new_n684));
  XOR2_X1   g483(.A(new_n683), .B(new_n684), .Z(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  OR2_X1    g485(.A1(new_n681), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n681), .A2(new_n686), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n663), .A2(new_n690), .ZN(new_n691));
  AND3_X1   g490(.A1(new_n565), .A2(new_n610), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(new_n483), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g493(.A1(new_n692), .A2(new_n484), .ZN(new_n695));
  AND2_X1   g494(.A1(new_n695), .A2(G8gat), .ZN(new_n696));
  XNOR2_X1  g495(.A(KEYINPUT16), .B(G8gat), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(KEYINPUT42), .B1(new_n696), .B2(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n699), .B1(KEYINPUT42), .B2(new_n698), .ZN(G1325gat));
  INV_X1    g499(.A(G15gat), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n692), .A2(new_n701), .A3(new_n309), .ZN(new_n702));
  AND2_X1   g501(.A1(new_n692), .A2(new_n511), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n702), .B1(new_n703), .B2(new_n701), .ZN(G1326gat));
  INV_X1    g503(.A(new_n475), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n692), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g505(.A(KEYINPUT43), .B(G22gat), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n706), .B(new_n707), .ZN(G1327gat));
  NOR3_X1   g507(.A1(new_n609), .A2(new_n632), .A3(new_n690), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n662), .A2(KEYINPUT44), .ZN(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT110), .ZN(new_n713));
  INV_X1    g512(.A(new_n549), .ZN(new_n714));
  AOI21_X1  g513(.A(KEYINPUT90), .B1(new_n530), .B2(new_n545), .ZN(new_n715));
  OAI22_X1  g514(.A1(new_n714), .A2(new_n715), .B1(new_n531), .B2(new_n532), .ZN(new_n716));
  OAI211_X1 g515(.A(new_n532), .B(KEYINPUT38), .C1(new_n536), .C2(new_n539), .ZN(new_n717));
  INV_X1    g516(.A(new_n515), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n716), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n561), .A2(new_n484), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n475), .A2(new_n721), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n513), .B1(new_n720), .B2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT109), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n506), .A2(new_n724), .ZN(new_n725));
  NAND4_X1  g524(.A1(new_n472), .A2(new_n505), .A3(KEYINPUT109), .A4(new_n474), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n713), .B1(new_n723), .B2(new_n727), .ZN(new_n728));
  AND2_X1   g527(.A1(new_n725), .A2(new_n726), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n511), .B1(new_n551), .B2(new_n562), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n729), .A2(KEYINPUT110), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n728), .A2(new_n731), .ZN(new_n732));
  NAND4_X1  g531(.A1(new_n309), .A2(new_n435), .A3(new_n202), .A4(new_n475), .ZN(new_n733));
  INV_X1    g532(.A(new_n497), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n496), .B1(new_n493), .B2(KEYINPUT35), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n733), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n712), .B1(new_n732), .B2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(new_n662), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n738), .B1(new_n498), .B2(new_n564), .ZN(new_n739));
  AOI22_X1  g538(.A1(new_n737), .A2(KEYINPUT111), .B1(KEYINPUT44), .B2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT111), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n495), .A2(new_n497), .ZN(new_n742));
  AOI22_X1  g541(.A1(new_n728), .A2(new_n731), .B1(new_n742), .B2(new_n733), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n741), .B1(new_n743), .B2(new_n712), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n710), .B1(new_n740), .B2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  OAI21_X1  g545(.A(G29gat), .B1(new_n746), .B2(new_n502), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n739), .A2(new_n710), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n748), .A2(new_n574), .A3(new_n483), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(KEYINPUT45), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n747), .A2(new_n750), .ZN(G1328gat));
  INV_X1    g550(.A(KEYINPUT112), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n565), .A2(new_n738), .A3(new_n709), .ZN(new_n753));
  INV_X1    g552(.A(new_n484), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n754), .A2(G36gat), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n752), .B1(new_n753), .B2(new_n756), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n748), .A2(KEYINPUT112), .A3(new_n755), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT113), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n760), .A2(KEYINPUT46), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n759), .B(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n760), .A2(KEYINPUT46), .ZN(new_n763));
  OAI21_X1  g562(.A(G36gat), .B1(new_n746), .B2(new_n754), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n762), .A2(new_n763), .A3(new_n764), .ZN(G1329gat));
  NOR3_X1   g564(.A1(new_n723), .A2(new_n713), .A3(new_n727), .ZN(new_n766));
  AOI21_X1  g565(.A(KEYINPUT110), .B1(new_n729), .B2(new_n730), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n736), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n768), .A2(KEYINPUT111), .A3(new_n711), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n739), .A2(KEYINPUT44), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n744), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n771), .A2(new_n511), .A3(new_n709), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT114), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n771), .A2(KEYINPUT114), .A3(new_n511), .A4(new_n709), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n774), .A2(G43gat), .A3(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(new_n309), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n753), .A2(G43gat), .A3(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT47), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n776), .A2(new_n780), .ZN(new_n781));
  AND2_X1   g580(.A1(new_n772), .A2(G43gat), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n779), .B1(new_n782), .B2(new_n778), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n781), .A2(new_n783), .ZN(G1330gat));
  XNOR2_X1  g583(.A(KEYINPUT116), .B(KEYINPUT48), .ZN(new_n785));
  INV_X1    g584(.A(G50gat), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n786), .B1(new_n745), .B2(new_n705), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n753), .A2(G50gat), .A3(new_n475), .ZN(new_n788));
  OAI211_X1 g587(.A(KEYINPUT115), .B(new_n785), .C1(new_n787), .C2(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(new_n785), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n771), .A2(new_n705), .A3(new_n709), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n788), .B1(new_n791), .B2(G50gat), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT115), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n790), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n789), .A2(new_n794), .ZN(G1331gat));
  NOR3_X1   g594(.A1(new_n610), .A2(new_n663), .A3(new_n689), .ZN(new_n796));
  AND2_X1   g595(.A1(new_n768), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(new_n483), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n798), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g598(.A1(new_n768), .A2(new_n796), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n800), .A2(new_n754), .ZN(new_n801));
  NOR2_X1   g600(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n802));
  AND2_X1   g601(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n801), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n804), .B1(new_n801), .B2(new_n802), .ZN(G1333gat));
  NAND3_X1  g604(.A1(new_n797), .A2(KEYINPUT118), .A3(new_n309), .ZN(new_n806));
  INV_X1    g605(.A(G71gat), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT118), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n808), .B1(new_n800), .B2(new_n777), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n806), .A2(new_n807), .A3(new_n809), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n513), .A2(new_n807), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n797), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n812), .A2(KEYINPUT117), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT117), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n814), .B1(new_n797), .B2(new_n811), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n810), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  XNOR2_X1  g615(.A(new_n816), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g616(.A1(new_n797), .A2(new_n705), .ZN(new_n818));
  XNOR2_X1  g617(.A(new_n818), .B(G78gat), .ZN(G1335gat));
  INV_X1    g618(.A(new_n632), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(new_n609), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n821), .A2(new_n689), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n771), .A2(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(G85gat), .B1(new_n823), .B2(new_n502), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n821), .A2(new_n662), .ZN(new_n825));
  AND3_X1   g624(.A1(new_n768), .A2(KEYINPUT51), .A3(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(KEYINPUT51), .B1(new_n768), .B2(new_n825), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  XNOR2_X1  g627(.A(new_n828), .B(KEYINPUT119), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n690), .A2(new_n636), .A3(new_n483), .ZN(new_n830));
  XNOR2_X1  g629(.A(new_n830), .B(KEYINPUT120), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n824), .B1(new_n829), .B2(new_n831), .ZN(G1336gat));
  XNOR2_X1  g631(.A(KEYINPUT121), .B(KEYINPUT52), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n771), .A2(new_n484), .A3(new_n822), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(G92gat), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n690), .A2(new_n637), .A3(new_n484), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n828), .A2(new_n838), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n834), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  OAI211_X1 g639(.A(new_n836), .B(new_n833), .C1(new_n828), .C2(new_n838), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(G1337gat));
  OAI21_X1  g641(.A(G99gat), .B1(new_n823), .B2(new_n513), .ZN(new_n843));
  OR3_X1    g642(.A1(new_n777), .A2(G99gat), .A3(new_n689), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n843), .B1(new_n829), .B2(new_n844), .ZN(G1338gat));
  INV_X1    g644(.A(KEYINPUT122), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n846), .A2(KEYINPUT53), .ZN(new_n847));
  OAI211_X1 g646(.A(new_n705), .B(new_n690), .C1(new_n826), .C2(new_n827), .ZN(new_n848));
  INV_X1    g647(.A(G106gat), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n847), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n846), .A2(KEYINPUT53), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n771), .A2(G106gat), .A3(new_n705), .A4(new_n822), .ZN(new_n852));
  AND3_X1   g651(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n851), .B1(new_n850), .B2(new_n852), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n853), .A2(new_n854), .ZN(G1339gat));
  NOR2_X1   g654(.A1(new_n590), .A2(new_n591), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n593), .A2(new_n594), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n603), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n608), .A2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT54), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n679), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n677), .A2(new_n667), .A3(new_n678), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n685), .B1(new_n679), .B2(new_n860), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT55), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  OR3_X1    g666(.A1(new_n679), .A2(new_n680), .A3(new_n686), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n863), .A2(KEYINPUT55), .A3(new_n864), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  OAI221_X1 g669(.A(new_n662), .B1(new_n689), .B2(new_n859), .C1(new_n609), .C2(new_n870), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n869), .A2(new_n868), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n872), .A2(new_n608), .A3(new_n867), .A4(new_n858), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n632), .B1(new_n873), .B2(new_n738), .ZN(new_n874));
  AOI22_X1  g673(.A1(new_n871), .A2(new_n874), .B1(new_n691), .B2(new_n609), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n475), .A2(new_n486), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  NOR4_X1   g676(.A1(new_n875), .A2(new_n502), .A3(new_n484), .A4(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(G113gat), .B1(new_n878), .B2(new_n610), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT123), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n880), .B1(new_n875), .B2(new_n705), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n609), .A2(new_n632), .A3(new_n662), .A4(new_n689), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n873), .A2(new_n738), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(new_n820), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n662), .B1(new_n859), .B2(new_n689), .ZN(new_n885));
  INV_X1    g684(.A(new_n870), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n885), .B1(new_n610), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n882), .B1(new_n884), .B2(new_n887), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n888), .A2(KEYINPUT123), .A3(new_n475), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n777), .B1(new_n881), .B2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n484), .A2(new_n502), .ZN(new_n892));
  INV_X1    g691(.A(new_n892), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n609), .A2(new_n276), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n879), .B1(new_n894), .B2(new_n895), .ZN(G1340gat));
  AOI21_X1  g695(.A(G120gat), .B1(new_n878), .B2(new_n690), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n689), .A2(new_n274), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n897), .B1(new_n894), .B2(new_n898), .ZN(G1341gat));
  NAND3_X1  g698(.A1(new_n878), .A2(new_n269), .A3(new_n632), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n891), .A2(new_n820), .A3(new_n893), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n900), .B1(new_n901), .B2(new_n269), .ZN(G1342gat));
  NAND3_X1  g701(.A1(new_n878), .A2(new_n271), .A3(new_n738), .ZN(new_n903));
  XOR2_X1   g702(.A(new_n903), .B(KEYINPUT56), .Z(new_n904));
  NOR3_X1   g703(.A1(new_n891), .A2(new_n662), .A3(new_n893), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n904), .B1(new_n271), .B2(new_n905), .ZN(G1343gat));
  INV_X1    g705(.A(new_n315), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n888), .A2(new_n705), .ZN(new_n908));
  OR2_X1    g707(.A1(new_n908), .A2(KEYINPUT57), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n511), .B1(new_n908), .B2(KEYINPUT57), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n909), .A2(new_n892), .A3(new_n910), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n907), .B1(new_n911), .B2(new_n609), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n513), .A2(new_n705), .ZN(new_n913));
  NOR4_X1   g712(.A1(new_n875), .A2(new_n502), .A3(new_n484), .A4(new_n913), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n914), .A2(new_n331), .A3(new_n610), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n912), .A2(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT58), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n917), .B1(new_n915), .B2(KEYINPUT124), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n916), .B(new_n918), .ZN(G1344gat));
  OAI21_X1  g718(.A(G148gat), .B1(new_n911), .B2(new_n689), .ZN(new_n920));
  XNOR2_X1  g719(.A(new_n920), .B(KEYINPUT59), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n914), .A2(new_n312), .A3(new_n690), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(G1345gat));
  NAND2_X1  g722(.A1(new_n632), .A2(G155gat), .ZN(new_n924));
  XNOR2_X1  g723(.A(new_n924), .B(KEYINPUT125), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n914), .A2(new_n632), .ZN(new_n926));
  OAI22_X1  g725(.A1(new_n911), .A2(new_n925), .B1(new_n926), .B2(G155gat), .ZN(new_n927));
  INV_X1    g726(.A(new_n927), .ZN(G1346gat));
  OAI21_X1  g727(.A(G162gat), .B1(new_n911), .B2(new_n662), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n914), .A2(new_n319), .A3(new_n738), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(G1347gat));
  NOR4_X1   g730(.A1(new_n875), .A2(new_n483), .A3(new_n754), .A4(new_n877), .ZN(new_n932));
  AOI21_X1  g731(.A(G169gat), .B1(new_n932), .B2(new_n610), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n754), .A2(new_n483), .ZN(new_n934));
  AND2_X1   g733(.A1(new_n890), .A2(new_n934), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n610), .A2(G169gat), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n933), .B1(new_n935), .B2(new_n936), .ZN(G1348gat));
  AOI21_X1  g736(.A(G176gat), .B1(new_n932), .B2(new_n690), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n881), .A2(new_n889), .ZN(new_n939));
  AND4_X1   g738(.A1(G176gat), .A2(new_n309), .A3(new_n690), .A4(new_n934), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n938), .B1(new_n939), .B2(new_n940), .ZN(G1349gat));
  NAND4_X1  g740(.A1(new_n939), .A2(new_n309), .A3(new_n632), .A4(new_n934), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT126), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND4_X1  g743(.A1(new_n890), .A2(KEYINPUT126), .A3(new_n632), .A4(new_n934), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n944), .A2(G183gat), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n219), .A2(KEYINPUT27), .ZN(new_n947));
  NAND4_X1  g746(.A1(new_n932), .A2(new_n263), .A3(new_n947), .A4(new_n632), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(KEYINPUT60), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT60), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n946), .A2(new_n951), .A3(new_n948), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n950), .A2(new_n952), .ZN(G1350gat));
  NAND3_X1  g752(.A1(new_n932), .A2(new_n220), .A3(new_n738), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT61), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n935), .A2(new_n738), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n955), .B1(new_n956), .B2(G190gat), .ZN(new_n957));
  AOI211_X1 g756(.A(KEYINPUT61), .B(new_n220), .C1(new_n935), .C2(new_n738), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n954), .B1(new_n957), .B2(new_n958), .ZN(G1351gat));
  NAND3_X1  g758(.A1(new_n909), .A2(new_n910), .A3(new_n934), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n610), .A2(G197gat), .ZN(new_n961));
  NOR4_X1   g760(.A1(new_n875), .A2(new_n483), .A3(new_n754), .A4(new_n913), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n962), .A2(new_n610), .ZN(new_n963));
  OAI22_X1  g762(.A1(new_n960), .A2(new_n961), .B1(new_n963), .B2(G197gat), .ZN(new_n964));
  INV_X1    g763(.A(new_n964), .ZN(G1352gat));
  INV_X1    g764(.A(G204gat), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n962), .A2(new_n966), .A3(new_n690), .ZN(new_n967));
  XOR2_X1   g766(.A(new_n967), .B(KEYINPUT62), .Z(new_n968));
  NOR2_X1   g767(.A1(new_n960), .A2(new_n689), .ZN(new_n969));
  AND2_X1   g768(.A1(new_n969), .A2(KEYINPUT127), .ZN(new_n970));
  OAI21_X1  g769(.A(G204gat), .B1(new_n969), .B2(KEYINPUT127), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n968), .B1(new_n970), .B2(new_n971), .ZN(G1353gat));
  OAI21_X1  g771(.A(G211gat), .B1(new_n960), .B2(new_n820), .ZN(new_n973));
  INV_X1    g772(.A(KEYINPUT63), .ZN(new_n974));
  XNOR2_X1  g773(.A(new_n973), .B(new_n974), .ZN(new_n975));
  INV_X1    g774(.A(G211gat), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n962), .A2(new_n976), .A3(new_n632), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n975), .A2(new_n977), .ZN(G1354gat));
  OAI21_X1  g777(.A(G218gat), .B1(new_n960), .B2(new_n662), .ZN(new_n979));
  INV_X1    g778(.A(G218gat), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n962), .A2(new_n980), .A3(new_n738), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n979), .A2(new_n981), .ZN(G1355gat));
endmodule


