

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n588, n589, n590, n591,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760;

  INV_X1 U381 ( .A(KEYINPUT108), .ZN(n361) );
  NAND2_X2 U382 ( .A1(n682), .A2(n683), .ZN(n362) );
  BUF_X1 U383 ( .A(G143), .Z(n759) );
  INV_X1 U384 ( .A(G128), .ZN(n467) );
  XNOR2_X2 U385 ( .A(n545), .B(n396), .ZN(n554) );
  XNOR2_X2 U386 ( .A(n377), .B(KEYINPUT88), .ZN(n545) );
  XNOR2_X2 U387 ( .A(KEYINPUT73), .B(KEYINPUT22), .ZN(n439) );
  XNOR2_X2 U388 ( .A(KEYINPUT15), .B(G902), .ZN(n608) );
  XNOR2_X1 U389 ( .A(n360), .B(KEYINPUT46), .ZN(n593) );
  NAND2_X1 U390 ( .A1(n760), .A2(n757), .ZN(n360) );
  NOR2_X2 U391 ( .A1(n738), .A2(n749), .ZN(n665) );
  XNOR2_X2 U392 ( .A(n588), .B(KEYINPUT41), .ZN(n702) );
  XNOR2_X2 U393 ( .A(n362), .B(n361), .ZN(n687) );
  AND2_X2 U394 ( .A1(n635), .A2(n634), .ZN(n626) );
  XNOR2_X1 U395 ( .A(KEYINPUT77), .B(KEYINPUT98), .ZN(n441) );
  XNOR2_X1 U396 ( .A(G122), .B(G104), .ZN(n406) );
  XNOR2_X1 U397 ( .A(G146), .B(G101), .ZN(n458) );
  INV_X1 U398 ( .A(G104), .ZN(n381) );
  INV_X1 U399 ( .A(G953), .ZN(n703) );
  INV_X1 U400 ( .A(n558), .ZN(n559) );
  XNOR2_X1 U401 ( .A(n479), .B(n478), .ZN(n669) );
  NOR2_X1 U402 ( .A1(n594), .A2(n593), .ZN(n595) );
  NOR2_X1 U403 ( .A1(n572), .A2(n571), .ZN(n577) );
  NOR2_X1 U404 ( .A1(n504), .A2(n543), .ZN(n492) );
  NOR2_X1 U405 ( .A1(n667), .A2(n666), .ZN(n490) );
  XNOR2_X1 U406 ( .A(n673), .B(KEYINPUT6), .ZN(n543) );
  BUF_X1 U407 ( .A(n485), .Z(n673) );
  XNOR2_X1 U408 ( .A(n422), .B(n421), .ZN(n513) );
  OR2_X1 U409 ( .A1(n669), .A2(n670), .ZN(n666) );
  AND2_X1 U410 ( .A1(n369), .A2(n372), .ZN(n368) );
  XNOR2_X1 U411 ( .A(n403), .B(KEYINPUT94), .ZN(n404) );
  XNOR2_X1 U412 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X2 U413 ( .A(n616), .B(KEYINPUT90), .ZN(n662) );
  XNOR2_X1 U414 ( .A(n431), .B(KEYINPUT4), .ZN(n453) );
  XNOR2_X2 U415 ( .A(G146), .B(G125), .ZN(n410) );
  XOR2_X2 U416 ( .A(KEYINPUT5), .B(KEYINPUT99), .Z(n442) );
  XNOR2_X2 U417 ( .A(KEYINPUT67), .B(KEYINPUT10), .ZN(n409) );
  XNOR2_X2 U418 ( .A(G116), .B(G113), .ZN(n375) );
  XNOR2_X1 U419 ( .A(G110), .B(G107), .ZN(n382) );
  NAND2_X1 U420 ( .A1(n635), .A2(n634), .ZN(n655) );
  NAND2_X1 U421 ( .A1(n611), .A2(n610), .ZN(n635) );
  BUF_X1 U422 ( .A(n565), .Z(n580) );
  XNOR2_X1 U423 ( .A(n376), .B(n375), .ZN(n446) );
  XNOR2_X1 U424 ( .A(n379), .B(G119), .ZN(n376) );
  NAND2_X2 U425 ( .A1(n368), .A2(n367), .ZN(n507) );
  NAND2_X1 U426 ( .A1(n371), .A2(n475), .ZN(n370) );
  XNOR2_X1 U427 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n386) );
  INV_X1 U428 ( .A(KEYINPUT33), .ZN(n491) );
  XNOR2_X1 U429 ( .A(n446), .B(n380), .ZN(n732) );
  INV_X1 U430 ( .A(KEYINPUT85), .ZN(n534) );
  XNOR2_X1 U431 ( .A(n453), .B(n388), .ZN(n366) );
  XNOR2_X1 U432 ( .A(n498), .B(KEYINPUT35), .ZN(n527) );
  INV_X1 U433 ( .A(KEYINPUT34), .ZN(n494) );
  INV_X1 U434 ( .A(n613), .ZN(n614) );
  XNOR2_X1 U435 ( .A(n419), .B(n418), .ZN(n642) );
  XOR2_X1 U436 ( .A(n734), .B(n383), .Z(n363) );
  INV_X1 U437 ( .A(n608), .ZN(n374) );
  BUF_X1 U438 ( .A(n446), .Z(n364) );
  BUF_X1 U439 ( .A(n612), .Z(n738) );
  BUF_X1 U440 ( .A(n484), .Z(n519) );
  XNOR2_X1 U441 ( .A(n732), .B(n363), .ZN(n365) );
  OR2_X2 U442 ( .A1(n656), .A2(n374), .ZN(n373) );
  XNOR2_X1 U443 ( .A(n365), .B(n366), .ZN(n656) );
  OR2_X1 U444 ( .A1(n648), .A2(n370), .ZN(n367) );
  NAND2_X1 U445 ( .A1(n648), .A2(n462), .ZN(n369) );
  INV_X1 U446 ( .A(n462), .ZN(n371) );
  NAND2_X1 U447 ( .A1(n462), .A2(G902), .ZN(n372) );
  XNOR2_X2 U448 ( .A(n507), .B(n463), .ZN(n667) );
  XNOR2_X2 U449 ( .A(n456), .B(n469), .ZN(n748) );
  XNOR2_X2 U450 ( .A(n453), .B(n452), .ZN(n456) );
  XNOR2_X2 U451 ( .A(n384), .B(n467), .ZN(n431) );
  XNOR2_X2 U452 ( .A(n373), .B(n392), .ZN(n565) );
  NOR2_X2 U453 ( .A1(n565), .A2(n395), .ZN(n377) );
  XNOR2_X1 U454 ( .A(n615), .B(n614), .ZN(n617) );
  NAND2_X2 U455 ( .A1(n484), .A2(n482), .ZN(n483) );
  XNOR2_X2 U456 ( .A(n483), .B(KEYINPUT32), .ZN(n624) );
  AND2_X1 U457 ( .A1(n476), .A2(G217), .ZN(n378) );
  INV_X1 U458 ( .A(G137), .ZN(n443) );
  XNOR2_X1 U459 ( .A(n444), .B(n443), .ZN(n445) );
  NOR2_X1 U460 ( .A1(G953), .A2(G237), .ZN(n415) );
  INV_X1 U461 ( .A(KEYINPUT78), .ZN(n605) );
  XNOR2_X1 U462 ( .A(n364), .B(n445), .ZN(n450) );
  XNOR2_X1 U463 ( .A(n749), .B(n605), .ZN(n606) );
  XNOR2_X1 U464 ( .A(n492), .B(n491), .ZN(n692) );
  XNOR2_X1 U465 ( .A(n417), .B(n416), .ZN(n418) );
  BUF_X1 U466 ( .A(n692), .Z(n701) );
  XNOR2_X1 U467 ( .A(n455), .B(G472), .ZN(n485) );
  BUF_X1 U468 ( .A(n627), .Z(n628) );
  XNOR2_X1 U469 ( .A(n420), .B(n639), .ZN(n421) );
  XNOR2_X1 U470 ( .A(n472), .B(n471), .ZN(n473) );
  BUF_X1 U471 ( .A(n648), .Z(n650) );
  INV_X1 U472 ( .A(KEYINPUT39), .ZN(n582) );
  XNOR2_X1 U473 ( .A(n474), .B(n473), .ZN(n637) );
  INV_X1 U474 ( .A(KEYINPUT123), .ZN(n618) );
  XNOR2_X2 U475 ( .A(G101), .B(KEYINPUT3), .ZN(n379) );
  XNOR2_X1 U476 ( .A(KEYINPUT16), .B(G122), .ZN(n380) );
  XNOR2_X1 U477 ( .A(n382), .B(n381), .ZN(n734) );
  XNOR2_X1 U478 ( .A(KEYINPUT71), .B(KEYINPUT72), .ZN(n383) );
  XNOR2_X2 U479 ( .A(KEYINPUT82), .B(G143), .ZN(n384) );
  NAND2_X1 U480 ( .A1(n703), .A2(G224), .ZN(n385) );
  XNOR2_X1 U481 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U482 ( .A(n387), .B(n410), .ZN(n388) );
  NOR2_X1 U483 ( .A1(G902), .A2(G237), .ZN(n389) );
  XNOR2_X1 U484 ( .A(n389), .B(KEYINPUT76), .ZN(n394) );
  INV_X1 U485 ( .A(G210), .ZN(n654) );
  OR2_X1 U486 ( .A1(n394), .A2(n654), .ZN(n391) );
  INV_X1 U487 ( .A(KEYINPUT91), .ZN(n390) );
  INV_X1 U488 ( .A(G214), .ZN(n393) );
  OR2_X1 U489 ( .A1(n394), .A2(n393), .ZN(n683) );
  INV_X1 U490 ( .A(n683), .ZN(n395) );
  XNOR2_X1 U491 ( .A(KEYINPUT66), .B(KEYINPUT19), .ZN(n396) );
  NAND2_X1 U492 ( .A1(G237), .A2(G234), .ZN(n397) );
  XNOR2_X1 U493 ( .A(n397), .B(KEYINPUT92), .ZN(n398) );
  XNOR2_X1 U494 ( .A(KEYINPUT14), .B(n398), .ZN(n401) );
  NAND2_X1 U495 ( .A1(n401), .A2(G902), .ZN(n399) );
  XNOR2_X1 U496 ( .A(n399), .B(KEYINPUT93), .ZN(n536) );
  INV_X1 U497 ( .A(G898), .ZN(n400) );
  AND2_X1 U498 ( .A1(n400), .A2(G953), .ZN(n736) );
  AND2_X1 U499 ( .A1(n536), .A2(n736), .ZN(n402) );
  NAND2_X1 U500 ( .A1(G952), .A2(n401), .ZN(n699) );
  NOR2_X1 U501 ( .A1(G953), .A2(n699), .ZN(n538) );
  NOR2_X1 U502 ( .A1(n402), .A2(n538), .ZN(n403) );
  NOR2_X2 U503 ( .A1(n554), .A2(n404), .ZN(n405) );
  XNOR2_X2 U504 ( .A(n405), .B(KEYINPUT0), .ZN(n493) );
  XOR2_X1 U505 ( .A(KEYINPUT11), .B(KEYINPUT100), .Z(n407) );
  XNOR2_X1 U506 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U507 ( .A(KEYINPUT12), .B(n408), .Z(n413) );
  INV_X1 U508 ( .A(n409), .ZN(n411) );
  XNOR2_X1 U509 ( .A(n411), .B(n410), .ZN(n747) );
  XNOR2_X1 U510 ( .A(G131), .B(n747), .ZN(n412) );
  XNOR2_X1 U511 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U512 ( .A(n414), .B(G140), .Z(n419) );
  XOR2_X1 U513 ( .A(KEYINPUT79), .B(n415), .Z(n447) );
  NAND2_X1 U514 ( .A1(n447), .A2(G214), .ZN(n417) );
  XNOR2_X1 U515 ( .A(n759), .B(G113), .ZN(n416) );
  NOR2_X1 U516 ( .A1(G902), .A2(n642), .ZN(n422) );
  XNOR2_X1 U517 ( .A(KEYINPUT101), .B(KEYINPUT13), .ZN(n420) );
  INV_X1 U518 ( .A(G475), .ZN(n639) );
  XOR2_X1 U519 ( .A(KEYINPUT102), .B(KEYINPUT7), .Z(n424) );
  XNOR2_X1 U520 ( .A(G107), .B(KEYINPUT9), .ZN(n423) );
  XNOR2_X1 U521 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U522 ( .A(n425), .B(G134), .Z(n427) );
  XNOR2_X1 U523 ( .A(G116), .B(G122), .ZN(n426) );
  XNOR2_X1 U524 ( .A(n427), .B(n426), .ZN(n433) );
  NAND2_X1 U525 ( .A1(n703), .A2(G234), .ZN(n429) );
  INV_X1 U526 ( .A(KEYINPUT8), .ZN(n428) );
  XNOR2_X1 U527 ( .A(n429), .B(n428), .ZN(n470) );
  NAND2_X1 U528 ( .A1(n470), .A2(G217), .ZN(n430) );
  XNOR2_X1 U529 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U530 ( .A(n433), .B(n432), .ZN(n613) );
  INV_X1 U531 ( .A(G902), .ZN(n475) );
  NAND2_X1 U532 ( .A1(n613), .A2(n475), .ZN(n435) );
  XNOR2_X1 U533 ( .A(G478), .B(KEYINPUT103), .ZN(n434) );
  XNOR2_X1 U534 ( .A(n435), .B(n434), .ZN(n512) );
  INV_X1 U535 ( .A(n512), .ZN(n496) );
  NOR2_X1 U536 ( .A1(n513), .A2(n496), .ZN(n685) );
  NAND2_X1 U537 ( .A1(n608), .A2(G234), .ZN(n436) );
  XNOR2_X1 U538 ( .A(n436), .B(KEYINPUT20), .ZN(n476) );
  AND2_X1 U539 ( .A1(n476), .A2(G221), .ZN(n437) );
  XNOR2_X1 U540 ( .A(n437), .B(KEYINPUT21), .ZN(n540) );
  AND2_X1 U541 ( .A1(n685), .A2(n540), .ZN(n438) );
  NAND2_X1 U542 ( .A1(n493), .A2(n438), .ZN(n440) );
  XNOR2_X2 U543 ( .A(n440), .B(n439), .ZN(n484) );
  XNOR2_X1 U544 ( .A(n442), .B(n441), .ZN(n444) );
  NAND2_X1 U545 ( .A1(n447), .A2(G210), .ZN(n448) );
  XNOR2_X1 U546 ( .A(n448), .B(G146), .ZN(n449) );
  XNOR2_X1 U547 ( .A(n450), .B(n449), .ZN(n454) );
  XNOR2_X1 U548 ( .A(G134), .B(G131), .ZN(n451) );
  XNOR2_X1 U549 ( .A(n451), .B(KEYINPUT68), .ZN(n452) );
  XNOR2_X1 U550 ( .A(n454), .B(n456), .ZN(n627) );
  NAND2_X1 U551 ( .A1(n627), .A2(n475), .ZN(n455) );
  XNOR2_X1 U552 ( .A(n543), .B(KEYINPUT81), .ZN(n481) );
  XNOR2_X1 U553 ( .A(G140), .B(G137), .ZN(n469) );
  NAND2_X1 U554 ( .A1(n703), .A2(G227), .ZN(n457) );
  XNOR2_X1 U555 ( .A(n457), .B(KEYINPUT95), .ZN(n459) );
  XNOR2_X1 U556 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U557 ( .A(n363), .B(n460), .ZN(n461) );
  XNOR2_X1 U558 ( .A(n748), .B(n461), .ZN(n648) );
  XNOR2_X1 U559 ( .A(KEYINPUT70), .B(G469), .ZN(n462) );
  XOR2_X1 U560 ( .A(KEYINPUT64), .B(KEYINPUT1), .Z(n463) );
  INV_X1 U561 ( .A(n667), .ZN(n598) );
  XOR2_X1 U562 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n465) );
  XNOR2_X1 U563 ( .A(G110), .B(KEYINPUT96), .ZN(n464) );
  XNOR2_X1 U564 ( .A(n465), .B(n464), .ZN(n466) );
  XOR2_X1 U565 ( .A(n747), .B(n466), .Z(n474) );
  XNOR2_X1 U566 ( .A(n467), .B(G119), .ZN(n468) );
  XNOR2_X1 U567 ( .A(n469), .B(n468), .ZN(n472) );
  NAND2_X1 U568 ( .A1(G221), .A2(n470), .ZN(n471) );
  NAND2_X1 U569 ( .A1(n637), .A2(n475), .ZN(n479) );
  XOR2_X1 U570 ( .A(KEYINPUT25), .B(KEYINPUT80), .Z(n477) );
  XNOR2_X1 U571 ( .A(n477), .B(n378), .ZN(n478) );
  NAND2_X1 U572 ( .A1(n598), .A2(n669), .ZN(n480) );
  NOR2_X1 U573 ( .A1(n481), .A2(n480), .ZN(n482) );
  XNOR2_X1 U574 ( .A(n485), .B(KEYINPUT105), .ZN(n558) );
  NAND2_X1 U575 ( .A1(n558), .A2(n669), .ZN(n486) );
  NOR2_X1 U576 ( .A1(n598), .A2(n486), .ZN(n487) );
  NAND2_X1 U577 ( .A1(n519), .A2(n487), .ZN(n621) );
  NAND2_X1 U578 ( .A1(n624), .A2(n621), .ZN(n489) );
  INV_X1 U579 ( .A(KEYINPUT87), .ZN(n488) );
  XNOR2_X1 U580 ( .A(n489), .B(n488), .ZN(n523) );
  INV_X1 U581 ( .A(n540), .ZN(n670) );
  XNOR2_X1 U582 ( .A(n490), .B(KEYINPUT75), .ZN(n504) );
  BUF_X2 U583 ( .A(n493), .Z(n508) );
  NAND2_X1 U584 ( .A1(n692), .A2(n508), .ZN(n495) );
  XNOR2_X1 U585 ( .A(n495), .B(n494), .ZN(n497) );
  AND2_X1 U586 ( .A1(n513), .A2(n496), .ZN(n566) );
  NAND2_X1 U587 ( .A1(n497), .A2(n566), .ZN(n498) );
  NAND2_X1 U588 ( .A1(n527), .A2(KEYINPUT86), .ZN(n499) );
  NAND2_X1 U589 ( .A1(n499), .A2(KEYINPUT44), .ZN(n500) );
  NOR2_X1 U590 ( .A1(n523), .A2(n500), .ZN(n503) );
  INV_X1 U591 ( .A(KEYINPUT86), .ZN(n501) );
  NOR2_X1 U592 ( .A1(n501), .A2(KEYINPUT44), .ZN(n502) );
  NOR2_X1 U593 ( .A1(n503), .A2(n502), .ZN(n522) );
  INV_X1 U594 ( .A(n508), .ZN(n505) );
  INV_X1 U595 ( .A(n673), .ZN(n510) );
  OR2_X1 U596 ( .A1(n504), .A2(n510), .ZN(n676) );
  NOR2_X2 U597 ( .A1(n505), .A2(n676), .ZN(n506) );
  XNOR2_X1 U598 ( .A(n506), .B(KEYINPUT31), .ZN(n724) );
  INV_X1 U599 ( .A(n507), .ZN(n552) );
  NOR2_X1 U600 ( .A1(n552), .A2(n666), .ZN(n563) );
  NAND2_X1 U601 ( .A1(n508), .A2(n563), .ZN(n509) );
  XNOR2_X1 U602 ( .A(n509), .B(KEYINPUT97), .ZN(n511) );
  NAND2_X1 U603 ( .A1(n511), .A2(n510), .ZN(n712) );
  NAND2_X1 U604 ( .A1(n724), .A2(n712), .ZN(n514) );
  AND2_X1 U605 ( .A1(n513), .A2(n512), .ZN(n719) );
  NOR2_X1 U606 ( .A1(n513), .A2(n512), .ZN(n716) );
  NOR2_X1 U607 ( .A1(n719), .A2(n716), .ZN(n574) );
  INV_X1 U608 ( .A(n574), .ZN(n688) );
  NAND2_X1 U609 ( .A1(n514), .A2(n688), .ZN(n515) );
  XNOR2_X1 U610 ( .A(n515), .B(KEYINPUT104), .ZN(n520) );
  INV_X1 U611 ( .A(n669), .ZN(n516) );
  NAND2_X1 U612 ( .A1(n543), .A2(n516), .ZN(n517) );
  NOR2_X1 U613 ( .A1(n598), .A2(n517), .ZN(n518) );
  NAND2_X1 U614 ( .A1(n519), .A2(n518), .ZN(n622) );
  NAND2_X1 U615 ( .A1(n520), .A2(n622), .ZN(n521) );
  NOR2_X1 U616 ( .A1(n522), .A2(n521), .ZN(n532) );
  INV_X1 U617 ( .A(n523), .ZN(n525) );
  INV_X1 U618 ( .A(KEYINPUT44), .ZN(n524) );
  NAND2_X1 U619 ( .A1(n525), .A2(n524), .ZN(n526) );
  NAND2_X1 U620 ( .A1(n526), .A2(KEYINPUT86), .ZN(n530) );
  BUF_X1 U621 ( .A(n527), .Z(n528) );
  INV_X1 U622 ( .A(n528), .ZN(n529) );
  NAND2_X1 U623 ( .A1(n530), .A2(n529), .ZN(n531) );
  AND2_X2 U624 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X2 U625 ( .A(n533), .B(KEYINPUT45), .ZN(n612) );
  NOR2_X2 U626 ( .A1(n612), .A2(n608), .ZN(n535) );
  XNOR2_X1 U627 ( .A(n535), .B(n534), .ZN(n607) );
  NAND2_X1 U628 ( .A1(G953), .A2(n536), .ZN(n537) );
  NOR2_X1 U629 ( .A1(G900), .A2(n537), .ZN(n539) );
  NOR2_X1 U630 ( .A1(n539), .A2(n538), .ZN(n562) );
  NAND2_X1 U631 ( .A1(n669), .A2(n540), .ZN(n541) );
  NOR2_X1 U632 ( .A1(n562), .A2(n541), .ZN(n542) );
  XNOR2_X1 U633 ( .A(KEYINPUT69), .B(n542), .ZN(n550) );
  INV_X1 U634 ( .A(n719), .ZN(n722) );
  OR2_X1 U635 ( .A1(n722), .A2(n543), .ZN(n544) );
  NOR2_X1 U636 ( .A1(n550), .A2(n544), .ZN(n597) );
  BUF_X1 U637 ( .A(n545), .Z(n546) );
  NAND2_X1 U638 ( .A1(n597), .A2(n546), .ZN(n548) );
  XOR2_X1 U639 ( .A(KEYINPUT36), .B(KEYINPUT110), .Z(n547) );
  XNOR2_X1 U640 ( .A(n548), .B(n547), .ZN(n549) );
  NAND2_X1 U641 ( .A1(n549), .A2(n598), .ZN(n729) );
  NOR2_X1 U642 ( .A1(n550), .A2(n558), .ZN(n551) );
  XOR2_X1 U643 ( .A(KEYINPUT28), .B(n551), .Z(n553) );
  NOR2_X1 U644 ( .A1(n553), .A2(n552), .ZN(n589) );
  BUF_X1 U645 ( .A(n554), .Z(n555) );
  INV_X1 U646 ( .A(n555), .ZN(n556) );
  NAND2_X1 U647 ( .A1(n589), .A2(n556), .ZN(n573) );
  NAND2_X1 U648 ( .A1(n573), .A2(KEYINPUT47), .ZN(n557) );
  NAND2_X1 U649 ( .A1(n729), .A2(n557), .ZN(n572) );
  NAND2_X1 U650 ( .A1(KEYINPUT47), .A2(n574), .ZN(n569) );
  NAND2_X1 U651 ( .A1(n559), .A2(n683), .ZN(n560) );
  XNOR2_X1 U652 ( .A(n560), .B(KEYINPUT30), .ZN(n561) );
  NOR2_X1 U653 ( .A1(n562), .A2(n561), .ZN(n564) );
  NAND2_X1 U654 ( .A1(n564), .A2(n563), .ZN(n581) );
  INV_X1 U655 ( .A(n580), .ZN(n601) );
  NAND2_X1 U656 ( .A1(n566), .A2(n601), .ZN(n567) );
  OR2_X1 U657 ( .A1(n581), .A2(n567), .ZN(n568) );
  XNOR2_X2 U658 ( .A(KEYINPUT106), .B(n568), .ZN(n758) );
  NAND2_X1 U659 ( .A1(n569), .A2(n758), .ZN(n570) );
  XOR2_X1 U660 ( .A(KEYINPUT83), .B(n570), .Z(n571) );
  INV_X1 U661 ( .A(n573), .ZN(n720) );
  NOR2_X1 U662 ( .A1(KEYINPUT47), .A2(n574), .ZN(n575) );
  NAND2_X1 U663 ( .A1(n720), .A2(n575), .ZN(n576) );
  NAND2_X1 U664 ( .A1(n577), .A2(n576), .ZN(n594) );
  XOR2_X1 U665 ( .A(KEYINPUT107), .B(KEYINPUT40), .Z(n585) );
  INV_X1 U666 ( .A(KEYINPUT74), .ZN(n578) );
  XNOR2_X1 U667 ( .A(n578), .B(KEYINPUT38), .ZN(n579) );
  XNOR2_X1 U668 ( .A(n580), .B(n579), .ZN(n586) );
  NOR2_X1 U669 ( .A1(n586), .A2(n581), .ZN(n583) );
  XNOR2_X1 U670 ( .A(n583), .B(n582), .ZN(n596) );
  NAND2_X1 U671 ( .A1(n596), .A2(n719), .ZN(n584) );
  XNOR2_X1 U672 ( .A(n585), .B(n584), .ZN(n757) );
  XOR2_X1 U673 ( .A(KEYINPUT109), .B(KEYINPUT42), .Z(n591) );
  INV_X1 U674 ( .A(n586), .ZN(n682) );
  NAND2_X1 U675 ( .A1(n687), .A2(n685), .ZN(n588) );
  NAND2_X1 U676 ( .A1(n702), .A2(n589), .ZN(n590) );
  XNOR2_X1 U677 ( .A(n591), .B(n590), .ZN(n760) );
  XNOR2_X1 U678 ( .A(n595), .B(KEYINPUT48), .ZN(n604) );
  AND2_X1 U679 ( .A1(n596), .A2(n716), .ZN(n731) );
  NAND2_X1 U680 ( .A1(n597), .A2(n683), .ZN(n599) );
  NOR2_X1 U681 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U682 ( .A(n600), .B(KEYINPUT43), .ZN(n602) );
  NOR2_X1 U683 ( .A1(n602), .A2(n601), .ZN(n623) );
  NOR2_X1 U684 ( .A1(n731), .A2(n623), .ZN(n603) );
  NAND2_X1 U685 ( .A1(n604), .A2(n603), .ZN(n749) );
  NAND2_X1 U686 ( .A1(n607), .A2(n606), .ZN(n611) );
  NAND2_X1 U687 ( .A1(n374), .A2(KEYINPUT2), .ZN(n609) );
  XOR2_X1 U688 ( .A(KEYINPUT65), .B(n609), .Z(n610) );
  NAND2_X1 U689 ( .A1(n665), .A2(KEYINPUT2), .ZN(n634) );
  NAND2_X1 U690 ( .A1(n626), .A2(G478), .ZN(n615) );
  NOR2_X1 U691 ( .A1(n703), .A2(G952), .ZN(n616) );
  NOR2_X2 U692 ( .A1(n617), .A2(n662), .ZN(n619) );
  XNOR2_X1 U693 ( .A(n619), .B(n618), .ZN(G63) );
  XOR2_X1 U694 ( .A(G110), .B(KEYINPUT111), .Z(n620) );
  XNOR2_X1 U695 ( .A(n621), .B(n620), .ZN(G12) );
  XNOR2_X1 U696 ( .A(n622), .B(G101), .ZN(G3) );
  XOR2_X1 U697 ( .A(G140), .B(n623), .Z(G42) );
  BUF_X1 U698 ( .A(n624), .Z(n625) );
  XNOR2_X1 U699 ( .A(n625), .B(G119), .ZN(G21) );
  XOR2_X1 U700 ( .A(n528), .B(G122), .Z(G24) );
  NAND2_X1 U701 ( .A1(n626), .A2(G472), .ZN(n630) );
  XOR2_X1 U702 ( .A(KEYINPUT62), .B(n628), .Z(n629) );
  XNOR2_X1 U703 ( .A(n630), .B(n629), .ZN(n631) );
  NOR2_X2 U704 ( .A1(n631), .A2(n662), .ZN(n633) );
  XNOR2_X1 U705 ( .A(KEYINPUT89), .B(KEYINPUT63), .ZN(n632) );
  XNOR2_X1 U706 ( .A(n633), .B(n632), .ZN(G57) );
  INV_X1 U707 ( .A(n655), .ZN(n647) );
  NAND2_X1 U708 ( .A1(n647), .A2(G217), .ZN(n636) );
  XOR2_X1 U709 ( .A(n637), .B(n636), .Z(n638) );
  NOR2_X1 U710 ( .A1(n638), .A2(n662), .ZN(G66) );
  NOR2_X1 U711 ( .A1(n655), .A2(n639), .ZN(n644) );
  XNOR2_X1 U712 ( .A(KEYINPUT121), .B(KEYINPUT122), .ZN(n640) );
  XOR2_X1 U713 ( .A(n640), .B(KEYINPUT59), .Z(n641) );
  XNOR2_X1 U714 ( .A(n642), .B(n641), .ZN(n643) );
  XNOR2_X1 U715 ( .A(n644), .B(n643), .ZN(n645) );
  NOR2_X1 U716 ( .A1(n645), .A2(n662), .ZN(n646) );
  XNOR2_X1 U717 ( .A(n646), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U718 ( .A1(n647), .A2(G469), .ZN(n652) );
  XOR2_X1 U719 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n649) );
  XNOR2_X1 U720 ( .A(n650), .B(n649), .ZN(n651) );
  XNOR2_X1 U721 ( .A(n652), .B(n651), .ZN(n653) );
  NOR2_X1 U722 ( .A1(n653), .A2(n662), .ZN(G54) );
  NOR2_X1 U723 ( .A1(n655), .A2(n654), .ZN(n661) );
  BUF_X1 U724 ( .A(n656), .Z(n657) );
  XNOR2_X1 U725 ( .A(KEYINPUT84), .B(KEYINPUT54), .ZN(n658) );
  XNOR2_X1 U726 ( .A(n658), .B(KEYINPUT55), .ZN(n659) );
  XNOR2_X1 U727 ( .A(n657), .B(n659), .ZN(n660) );
  XNOR2_X1 U728 ( .A(n661), .B(n660), .ZN(n663) );
  NOR2_X1 U729 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U730 ( .A(n664), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U731 ( .A(n665), .B(KEYINPUT2), .ZN(n708) );
  XNOR2_X1 U732 ( .A(KEYINPUT51), .B(KEYINPUT115), .ZN(n680) );
  NAND2_X1 U733 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U734 ( .A(n668), .B(KEYINPUT50), .ZN(n675) );
  AND2_X1 U735 ( .A1(n670), .A2(n669), .ZN(n671) );
  XOR2_X1 U736 ( .A(KEYINPUT49), .B(n671), .Z(n672) );
  NOR2_X1 U737 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U738 ( .A1(n675), .A2(n674), .ZN(n677) );
  NAND2_X1 U739 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U740 ( .A(n678), .B(KEYINPUT114), .ZN(n679) );
  XNOR2_X1 U741 ( .A(n680), .B(n679), .ZN(n681) );
  NAND2_X1 U742 ( .A1(n681), .A2(n702), .ZN(n695) );
  NOR2_X1 U743 ( .A1(n683), .A2(n682), .ZN(n684) );
  XOR2_X1 U744 ( .A(KEYINPUT116), .B(n684), .Z(n686) );
  NAND2_X1 U745 ( .A1(n686), .A2(n685), .ZN(n690) );
  NAND2_X1 U746 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U747 ( .A1(n690), .A2(n689), .ZN(n691) );
  XOR2_X1 U748 ( .A(KEYINPUT117), .B(n691), .Z(n693) );
  NAND2_X1 U749 ( .A1(n693), .A2(n701), .ZN(n694) );
  NAND2_X1 U750 ( .A1(n695), .A2(n694), .ZN(n697) );
  XOR2_X1 U751 ( .A(KEYINPUT52), .B(KEYINPUT118), .Z(n696) );
  XNOR2_X1 U752 ( .A(n697), .B(n696), .ZN(n698) );
  NOR2_X1 U753 ( .A1(n699), .A2(n698), .ZN(n700) );
  XOR2_X1 U754 ( .A(KEYINPUT119), .B(n700), .Z(n706) );
  NAND2_X1 U755 ( .A1(n702), .A2(n701), .ZN(n704) );
  NAND2_X1 U756 ( .A1(n704), .A2(n703), .ZN(n705) );
  NOR2_X1 U757 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U758 ( .A1(n708), .A2(n707), .ZN(n710) );
  XOR2_X1 U759 ( .A(KEYINPUT120), .B(KEYINPUT53), .Z(n709) );
  XNOR2_X1 U760 ( .A(n710), .B(n709), .ZN(G75) );
  NOR2_X1 U761 ( .A1(n722), .A2(n712), .ZN(n711) );
  XOR2_X1 U762 ( .A(G104), .B(n711), .Z(G6) );
  INV_X1 U763 ( .A(n716), .ZN(n725) );
  NOR2_X1 U764 ( .A1(n725), .A2(n712), .ZN(n714) );
  XNOR2_X1 U765 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n713) );
  XNOR2_X1 U766 ( .A(n714), .B(n713), .ZN(n715) );
  XNOR2_X1 U767 ( .A(G107), .B(n715), .ZN(G9) );
  XOR2_X1 U768 ( .A(G128), .B(KEYINPUT29), .Z(n718) );
  NAND2_X1 U769 ( .A1(n720), .A2(n716), .ZN(n717) );
  XNOR2_X1 U770 ( .A(n718), .B(n717), .ZN(G30) );
  NAND2_X1 U771 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U772 ( .A(n721), .B(G146), .ZN(G48) );
  NOR2_X1 U773 ( .A1(n722), .A2(n724), .ZN(n723) );
  XOR2_X1 U774 ( .A(G113), .B(n723), .Z(G15) );
  NOR2_X1 U775 ( .A1(n725), .A2(n724), .ZN(n726) );
  XOR2_X1 U776 ( .A(KEYINPUT112), .B(n726), .Z(n727) );
  XNOR2_X1 U777 ( .A(G116), .B(n727), .ZN(G18) );
  XNOR2_X1 U778 ( .A(KEYINPUT113), .B(KEYINPUT37), .ZN(n728) );
  XNOR2_X1 U779 ( .A(n729), .B(n728), .ZN(n730) );
  XNOR2_X1 U780 ( .A(G125), .B(n730), .ZN(G27) );
  XOR2_X1 U781 ( .A(G134), .B(n731), .Z(G36) );
  BUF_X1 U782 ( .A(n732), .Z(n733) );
  XNOR2_X1 U783 ( .A(n734), .B(KEYINPUT125), .ZN(n735) );
  XNOR2_X1 U784 ( .A(n733), .B(n735), .ZN(n737) );
  NOR2_X1 U785 ( .A1(n737), .A2(n736), .ZN(n745) );
  NOR2_X1 U786 ( .A1(n738), .A2(G953), .ZN(n739) );
  XOR2_X1 U787 ( .A(KEYINPUT124), .B(n739), .Z(n743) );
  NAND2_X1 U788 ( .A1(G953), .A2(G224), .ZN(n740) );
  XNOR2_X1 U789 ( .A(KEYINPUT61), .B(n740), .ZN(n741) );
  NAND2_X1 U790 ( .A1(n741), .A2(G898), .ZN(n742) );
  NAND2_X1 U791 ( .A1(n743), .A2(n742), .ZN(n744) );
  XNOR2_X1 U792 ( .A(n745), .B(n744), .ZN(n746) );
  XNOR2_X1 U793 ( .A(KEYINPUT126), .B(n746), .ZN(G69) );
  XOR2_X1 U794 ( .A(n748), .B(n747), .Z(n752) );
  XNOR2_X1 U795 ( .A(n749), .B(n752), .ZN(n750) );
  NOR2_X1 U796 ( .A1(G953), .A2(n750), .ZN(n751) );
  XNOR2_X1 U797 ( .A(n751), .B(KEYINPUT127), .ZN(n756) );
  XOR2_X1 U798 ( .A(G227), .B(n752), .Z(n753) );
  NAND2_X1 U799 ( .A1(n753), .A2(G900), .ZN(n754) );
  NAND2_X1 U800 ( .A1(n754), .A2(G953), .ZN(n755) );
  NAND2_X1 U801 ( .A1(n756), .A2(n755), .ZN(G72) );
  XNOR2_X1 U802 ( .A(G131), .B(n757), .ZN(G33) );
  XNOR2_X1 U803 ( .A(n759), .B(n758), .ZN(G45) );
  XNOR2_X1 U804 ( .A(G137), .B(n760), .ZN(G39) );
endmodule

