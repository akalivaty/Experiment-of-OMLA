//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 1 1 0 1 1 0 0 0 1 1 1 0 1 0 1 0 1 0 0 0 1 0 0 0 0 1 0 0 0 1 0 0 1 1 1 1 0 1 1 0 0 1 1 0 1 0 0 0 1 1 0 1 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:32 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n542, new_n543, new_n544, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n557, new_n558,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n576, new_n577, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n592, new_n595, new_n596, new_n598,
    new_n599, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n817, new_n818, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1153, new_n1154,
    new_n1155;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT64), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT65), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g024(.A1(G218), .A2(G219), .A3(G220), .A4(G221), .ZN(new_n450));
  XNOR2_X1  g025(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT67), .Z(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  NAND2_X1  g032(.A1(new_n452), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OR2_X1    g034(.A1(new_n454), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  AND2_X1   g037(.A1(KEYINPUT68), .A2(KEYINPUT3), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT68), .A2(KEYINPUT3), .ZN(new_n464));
  OAI21_X1  g039(.A(G2104), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT69), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n466), .B1(KEYINPUT3), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  OAI211_X1 g044(.A(new_n466), .B(G2104), .C1(new_n463), .C2(new_n464), .ZN(new_n470));
  AOI21_X1  g045(.A(G2105), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G137), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT3), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(G125), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n473), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n467), .A2(G2105), .ZN(new_n480));
  AOI22_X1  g055(.A1(new_n479), .A2(G2105), .B1(G101), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n472), .A2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G160));
  INV_X1    g058(.A(G2105), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n484), .B1(new_n469), .B2(new_n470), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  OR2_X1    g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G112), .C2(new_n484), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n489), .B1(G136), .B2(new_n471), .ZN(G162));
  INV_X1    g065(.A(KEYINPUT71), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n484), .A2(G138), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n492), .B1(new_n469), .B2(new_n470), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n491), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT68), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(new_n475), .ZN(new_n497));
  NAND2_X1  g072(.A1(KEYINPUT68), .A2(KEYINPUT3), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n467), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n474), .A2(KEYINPUT69), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n470), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n492), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n503), .A2(KEYINPUT71), .A3(KEYINPUT4), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n495), .A2(new_n504), .ZN(new_n505));
  NOR3_X1   g080(.A1(new_n477), .A2(KEYINPUT4), .A3(new_n492), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n501), .A2(G126), .A3(G2105), .ZN(new_n508));
  OAI21_X1  g083(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n509));
  INV_X1    g084(.A(G114), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n509), .B1(new_n510), .B2(G2105), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n508), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT70), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n508), .A2(KEYINPUT70), .A3(new_n512), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n505), .A2(new_n507), .B1(new_n515), .B2(new_n516), .ZN(G164));
  OAI21_X1  g092(.A(KEYINPUT5), .B1(KEYINPUT72), .B2(G543), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT73), .ZN(new_n519));
  INV_X1    g094(.A(G543), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND4_X1  g096(.A1(KEYINPUT72), .A2(KEYINPUT73), .A3(KEYINPUT5), .A4(G543), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  XNOR2_X1  g098(.A(KEYINPUT6), .B(G651), .ZN(new_n524));
  AND2_X1   g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(G543), .ZN(new_n526));
  INV_X1    g101(.A(new_n526), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n525), .A2(G88), .B1(G50), .B2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(G651), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n523), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n531), .A2(KEYINPUT74), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(KEYINPUT74), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(G166));
  NAND2_X1  g109(.A1(new_n525), .A2(G89), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n527), .A2(G51), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n523), .A2(G63), .A3(G651), .ZN(new_n537));
  XOR2_X1   g112(.A(KEYINPUT75), .B(KEYINPUT7), .Z(new_n538));
  NAND3_X1  g113(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n538), .B(new_n539), .ZN(new_n540));
  AND4_X1   g115(.A1(new_n535), .A2(new_n536), .A3(new_n537), .A4(new_n540), .ZN(G168));
  AOI22_X1  g116(.A1(new_n523), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n542), .A2(new_n529), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n525), .A2(G90), .B1(G52), .B2(new_n527), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(G301));
  INV_X1    g120(.A(G301), .ZN(G171));
  AND2_X1   g121(.A1(G68), .A2(G543), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n547), .B1(new_n523), .B2(G56), .ZN(new_n548));
  OR3_X1    g123(.A1(new_n548), .A2(KEYINPUT76), .A3(new_n529), .ZN(new_n549));
  OAI21_X1  g124(.A(KEYINPUT76), .B1(new_n548), .B2(new_n529), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n525), .A2(G81), .B1(G43), .B2(new_n527), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT77), .ZN(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND4_X1  g133(.A1(G319), .A2(G483), .A3(G661), .A4(new_n558), .ZN(G188));
  INV_X1    g134(.A(G53), .ZN(new_n560));
  OR3_X1    g135(.A1(new_n526), .A2(KEYINPUT9), .A3(new_n560), .ZN(new_n561));
  OAI21_X1  g136(.A(KEYINPUT9), .B1(new_n526), .B2(new_n560), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n561), .A2(new_n562), .B1(new_n525), .B2(G91), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n523), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n529), .B2(new_n564), .ZN(G299));
  INV_X1    g140(.A(G168), .ZN(G286));
  INV_X1    g141(.A(G166), .ZN(G303));
  NAND2_X1  g142(.A1(new_n525), .A2(G87), .ZN(new_n568));
  OAI21_X1  g143(.A(G651), .B1(new_n523), .B2(G74), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n527), .A2(G49), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(G288));
  AOI22_X1  g146(.A1(new_n523), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n572));
  OR2_X1    g147(.A1(new_n572), .A2(new_n529), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n525), .A2(G86), .B1(G48), .B2(new_n527), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(G305));
  AOI22_X1  g150(.A1(new_n525), .A2(G85), .B1(G47), .B2(new_n527), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n523), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n529), .B2(new_n577), .ZN(G290));
  INV_X1    g153(.A(G868), .ZN(new_n579));
  NOR2_X1   g154(.A1(G301), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n525), .A2(G92), .ZN(new_n581));
  XOR2_X1   g156(.A(new_n581), .B(KEYINPUT10), .Z(new_n582));
  NAND2_X1  g157(.A1(new_n523), .A2(G66), .ZN(new_n583));
  INV_X1    g158(.A(G79), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n584), .B2(new_n520), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n585), .A2(G651), .B1(G54), .B2(new_n527), .ZN(new_n586));
  AND3_X1   g161(.A1(new_n582), .A2(KEYINPUT78), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g162(.A(KEYINPUT78), .B1(new_n582), .B2(new_n586), .ZN(new_n588));
  OR2_X1    g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n580), .B1(new_n589), .B2(new_n579), .ZN(G284));
  XNOR2_X1  g165(.A(G284), .B(KEYINPUT79), .ZN(G321));
  NAND2_X1  g166(.A1(G299), .A2(new_n579), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n592), .B1(new_n579), .B2(G168), .ZN(G280));
  XOR2_X1   g168(.A(G280), .B(KEYINPUT80), .Z(G297));
  XOR2_X1   g169(.A(KEYINPUT81), .B(G559), .Z(new_n595));
  OAI21_X1  g170(.A(new_n589), .B1(G860), .B2(new_n595), .ZN(new_n596));
  XOR2_X1   g171(.A(new_n596), .B(KEYINPUT82), .Z(G148));
  NAND2_X1  g172(.A1(new_n589), .A2(new_n595), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(G868), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n599), .B1(G868), .B2(new_n553), .ZN(G323));
  XNOR2_X1  g175(.A(KEYINPUT83), .B(KEYINPUT11), .ZN(new_n601));
  XNOR2_X1  g176(.A(G323), .B(new_n601), .ZN(G282));
  NAND2_X1  g177(.A1(new_n471), .A2(G135), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n485), .A2(G123), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n484), .A2(G111), .ZN(new_n605));
  OAI21_X1  g180(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n606));
  OAI211_X1 g181(.A(new_n603), .B(new_n604), .C1(new_n605), .C2(new_n606), .ZN(new_n607));
  OR2_X1    g182(.A1(new_n607), .A2(G2096), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(G2096), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n484), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT12), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT13), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(G2100), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n608), .A2(new_n609), .A3(new_n613), .ZN(G156));
  XNOR2_X1  g189(.A(G2427), .B(G2438), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(G2430), .ZN(new_n616));
  XNOR2_X1  g191(.A(KEYINPUT15), .B(G2435), .ZN(new_n617));
  OR2_X1    g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n616), .A2(new_n617), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n618), .A2(KEYINPUT14), .A3(new_n619), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT85), .ZN(new_n621));
  INV_X1    g196(.A(G1341), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(G1348), .ZN(new_n624));
  XNOR2_X1  g199(.A(G2451), .B(G2454), .ZN(new_n625));
  XNOR2_X1  g200(.A(G2443), .B(G2446), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n624), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n624), .A2(new_n629), .ZN(new_n631));
  AND3_X1   g206(.A1(new_n630), .A2(G14), .A3(new_n631), .ZN(G401));
  XOR2_X1   g207(.A(G2072), .B(G2078), .Z(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(G2084), .B(G2090), .Z(new_n635));
  XNOR2_X1  g210(.A(G2067), .B(G2678), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT18), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n633), .B(KEYINPUT17), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n636), .B(KEYINPUT86), .ZN(new_n640));
  AND2_X1   g215(.A1(new_n640), .A2(new_n635), .ZN(new_n641));
  AOI21_X1  g216(.A(new_n638), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n635), .B1(new_n640), .B2(new_n633), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n643), .A2(KEYINPUT87), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n644), .B1(new_n640), .B2(new_n639), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n643), .A2(KEYINPUT87), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n642), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G2096), .B(G2100), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(G227));
  XNOR2_X1  g224(.A(G1971), .B(G1976), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT19), .ZN(new_n651));
  XNOR2_X1  g226(.A(G1956), .B(G2474), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT88), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1961), .B(G1966), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(KEYINPUT89), .B(KEYINPUT20), .Z(new_n657));
  OR2_X1    g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  OR2_X1    g233(.A1(new_n653), .A2(new_n655), .ZN(new_n659));
  AOI21_X1  g234(.A(new_n651), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n659), .A2(new_n656), .A3(new_n651), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n657), .B1(new_n656), .B2(new_n651), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT90), .ZN(new_n665));
  XOR2_X1   g240(.A(G1981), .B(G1986), .Z(new_n666));
  XNOR2_X1  g241(.A(G1991), .B(G1996), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n665), .B(new_n670), .ZN(G229));
  INV_X1    g246(.A(G29), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n672), .A2(KEYINPUT91), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(KEYINPUT91), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n675), .A2(G35), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n676), .B1(G162), .B2(new_n675), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(KEYINPUT29), .Z(new_n678));
  INV_X1    g253(.A(G2090), .ZN(new_n679));
  AND2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(G115), .A2(G2104), .ZN(new_n681));
  INV_X1    g256(.A(G127), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n681), .B1(new_n477), .B2(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(KEYINPUT98), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n484), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n685), .B1(new_n684), .B2(new_n683), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n471), .A2(G139), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n484), .A2(G103), .A3(G2104), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n688), .B(KEYINPUT25), .Z(new_n689));
  NAND3_X1  g264(.A1(new_n686), .A2(new_n687), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT99), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n691), .A2(new_n672), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n692), .B1(new_n672), .B2(G33), .ZN(new_n693));
  INV_X1    g268(.A(G2072), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n680), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT96), .B(G1348), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(G16), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G4), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(new_n589), .B2(new_n699), .ZN(new_n701));
  OAI221_X1 g276(.A(new_n696), .B1(new_n679), .B2(new_n678), .C1(new_n698), .C2(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(new_n675), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(G27), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n704), .B(KEYINPUT107), .Z(new_n705));
  INV_X1    g280(.A(G164), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n705), .B1(new_n706), .B2(new_n675), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT108), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n702), .B1(G2078), .B2(new_n708), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n708), .A2(G2078), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT24), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n711), .A2(G34), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(G34), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n703), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(new_n482), .B2(new_n672), .ZN(new_n715));
  INV_X1    g290(.A(G2084), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(KEYINPUT105), .Z(new_n718));
  NOR2_X1   g293(.A1(G171), .A2(new_n699), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(G5), .B2(new_n699), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  AND2_X1   g296(.A1(new_n672), .A2(G32), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT100), .B(KEYINPUT26), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT101), .ZN(new_n724));
  NAND3_X1  g299(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n724), .A2(new_n725), .ZN(new_n727));
  AOI22_X1  g302(.A1(new_n726), .A2(new_n727), .B1(G105), .B2(new_n480), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n471), .A2(G141), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n485), .A2(G129), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n728), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(KEYINPUT102), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT102), .ZN(new_n733));
  NAND4_X1  g308(.A1(new_n728), .A2(new_n733), .A3(new_n729), .A4(new_n730), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n722), .B1(new_n735), .B2(G29), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT27), .B(G1996), .ZN(new_n737));
  OAI221_X1 g312(.A(new_n718), .B1(new_n721), .B2(G1961), .C1(new_n736), .C2(new_n737), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT106), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n607), .A2(new_n703), .ZN(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT31), .B(G11), .ZN(new_n741));
  XOR2_X1   g316(.A(KEYINPUT104), .B(G28), .Z(new_n742));
  NOR2_X1   g317(.A1(new_n742), .A2(KEYINPUT30), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n742), .A2(KEYINPUT30), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(new_n672), .ZN(new_n745));
  NAND2_X1  g320(.A1(G168), .A2(G16), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G16), .B2(G21), .ZN(new_n747));
  XOR2_X1   g322(.A(KEYINPUT103), .B(G1966), .Z(new_n748));
  OAI221_X1 g323(.A(new_n741), .B1(new_n743), .B2(new_n745), .C1(new_n747), .C2(new_n748), .ZN(new_n749));
  AOI211_X1 g324(.A(new_n740), .B(new_n749), .C1(new_n748), .C2(new_n747), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n703), .A2(G26), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT28), .Z(new_n752));
  NAND2_X1  g327(.A1(new_n471), .A2(G140), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n485), .A2(G128), .ZN(new_n754));
  OR2_X1    g329(.A1(G104), .A2(G2105), .ZN(new_n755));
  OAI211_X1 g330(.A(new_n755), .B(G2104), .C1(G116), .C2(new_n484), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n753), .A2(new_n754), .A3(new_n756), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n752), .B1(new_n757), .B2(G29), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G2067), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n699), .A2(G20), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT23), .Z(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G299), .B2(G16), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(G1956), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n715), .A2(new_n716), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n721), .B2(G1961), .ZN(new_n765));
  NAND4_X1  g340(.A1(new_n750), .A2(new_n759), .A3(new_n763), .A4(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n701), .A2(new_n698), .ZN(new_n767));
  AOI22_X1  g342(.A1(new_n693), .A2(new_n694), .B1(new_n736), .B2(new_n737), .ZN(new_n768));
  INV_X1    g343(.A(G19), .ZN(new_n769));
  OR3_X1    g344(.A1(new_n769), .A2(KEYINPUT97), .A3(G16), .ZN(new_n770));
  OAI21_X1  g345(.A(KEYINPUT97), .B1(new_n769), .B2(G16), .ZN(new_n771));
  OAI211_X1 g346(.A(new_n770), .B(new_n771), .C1(new_n553), .C2(new_n699), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(new_n622), .ZN(new_n773));
  NAND3_X1  g348(.A1(new_n767), .A2(new_n768), .A3(new_n773), .ZN(new_n774));
  NOR3_X1   g349(.A1(new_n739), .A2(new_n766), .A3(new_n774), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n709), .A2(new_n710), .A3(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(G16), .A2(G22), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(G166), .B2(G16), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(G1971), .Z(new_n779));
  OR2_X1    g354(.A1(new_n779), .A2(KEYINPUT95), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n779), .A2(KEYINPUT95), .ZN(new_n781));
  NOR2_X1   g356(.A1(G6), .A2(G16), .ZN(new_n782));
  INV_X1    g357(.A(G305), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n782), .B1(new_n783), .B2(G16), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT32), .ZN(new_n785));
  INV_X1    g360(.A(G1981), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n699), .A2(G23), .ZN(new_n788));
  INV_X1    g363(.A(G288), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n788), .B1(new_n789), .B2(new_n699), .ZN(new_n790));
  XOR2_X1   g365(.A(KEYINPUT33), .B(G1976), .Z(new_n791));
  XOR2_X1   g366(.A(new_n790), .B(new_n791), .Z(new_n792));
  NAND4_X1  g367(.A1(new_n780), .A2(new_n781), .A3(new_n787), .A4(new_n792), .ZN(new_n793));
  OR2_X1    g368(.A1(new_n793), .A2(KEYINPUT34), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n793), .A2(KEYINPUT34), .ZN(new_n795));
  MUX2_X1   g370(.A(G24), .B(G290), .S(G16), .Z(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(G1986), .Z(new_n797));
  NAND2_X1  g372(.A1(new_n703), .A2(G25), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(KEYINPUT92), .Z(new_n799));
  OR2_X1    g374(.A1(G95), .A2(G2105), .ZN(new_n800));
  OAI211_X1 g375(.A(new_n800), .B(G2104), .C1(G107), .C2(new_n484), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(KEYINPUT93), .Z(new_n802));
  NAND2_X1  g377(.A1(new_n471), .A2(G131), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n485), .A2(G119), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n802), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(KEYINPUT94), .Z(new_n806));
  OAI21_X1  g381(.A(new_n799), .B1(new_n806), .B2(new_n703), .ZN(new_n807));
  XOR2_X1   g382(.A(KEYINPUT35), .B(G1991), .Z(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n797), .B1(new_n807), .B2(new_n809), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(new_n809), .B2(new_n807), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n794), .A2(new_n795), .A3(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n812), .A2(KEYINPUT36), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n812), .A2(KEYINPUT36), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n776), .B1(new_n814), .B2(new_n815), .ZN(G311));
  INV_X1    g391(.A(new_n776), .ZN(new_n817));
  INV_X1    g392(.A(new_n815), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n817), .B1(new_n818), .B2(new_n813), .ZN(G150));
  NAND2_X1  g394(.A1(new_n589), .A2(G559), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT38), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n525), .A2(G93), .ZN(new_n822));
  INV_X1    g397(.A(G55), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n822), .B1(new_n823), .B2(new_n526), .ZN(new_n824));
  AOI22_X1  g399(.A1(new_n523), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n825), .A2(new_n529), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n553), .A2(new_n827), .ZN(new_n828));
  OR2_X1    g403(.A1(new_n824), .A2(new_n826), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(new_n552), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n821), .B(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT39), .ZN(new_n833));
  AOI21_X1  g408(.A(G860), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(new_n833), .B2(new_n832), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n829), .A2(G860), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(KEYINPUT37), .Z(new_n837));
  NAND2_X1  g412(.A1(new_n835), .A2(new_n837), .ZN(G145));
  NAND2_X1  g413(.A1(new_n735), .A2(new_n757), .ZN(new_n839));
  INV_X1    g414(.A(new_n757), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n732), .A2(new_n734), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n471), .A2(G142), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n485), .A2(G130), .ZN(new_n844));
  OR2_X1    g419(.A1(G106), .A2(G2105), .ZN(new_n845));
  OAI211_X1 g420(.A(new_n845), .B(G2104), .C1(G118), .C2(new_n484), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n843), .A2(new_n844), .A3(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n842), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n839), .A2(new_n847), .A3(new_n841), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n805), .B(new_n611), .ZN(new_n851));
  AND3_X1   g426(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n851), .B1(new_n849), .B2(new_n850), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n691), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n849), .A2(new_n850), .ZN(new_n855));
  INV_X1    g430(.A(new_n851), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n691), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n506), .B1(new_n495), .B2(new_n504), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n861), .A2(new_n513), .ZN(new_n862));
  AND3_X1   g437(.A1(new_n854), .A2(new_n860), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n862), .B1(new_n854), .B2(new_n860), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n607), .B(new_n482), .ZN(new_n866));
  XOR2_X1   g441(.A(new_n866), .B(G162), .Z(new_n867));
  AOI21_X1  g442(.A(G37), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n854), .A2(new_n860), .ZN(new_n869));
  INV_X1    g444(.A(new_n862), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n854), .A2(new_n860), .A3(new_n862), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n867), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  AOI21_X1  g449(.A(KEYINPUT40), .B1(new_n868), .B2(new_n874), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n871), .A2(new_n867), .A3(new_n872), .ZN(new_n876));
  INV_X1    g451(.A(G37), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT40), .ZN(new_n879));
  NOR3_X1   g454(.A1(new_n878), .A2(new_n879), .A3(new_n873), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n875), .A2(new_n880), .ZN(G395));
  XNOR2_X1  g456(.A(new_n598), .B(new_n831), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n582), .A2(new_n586), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(G299), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(KEYINPUT41), .ZN(new_n885));
  OR2_X1    g460(.A1(new_n882), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n882), .ZN(new_n887));
  INV_X1    g462(.A(new_n884), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n886), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(KEYINPUT42), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT42), .ZN(new_n891));
  OAI211_X1 g466(.A(new_n886), .B(new_n891), .C1(new_n887), .C2(new_n888), .ZN(new_n892));
  XNOR2_X1  g467(.A(G166), .B(G288), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n783), .B(G290), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n893), .B(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  AND3_X1   g471(.A1(new_n890), .A2(new_n892), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n896), .B1(new_n890), .B2(new_n892), .ZN(new_n898));
  OAI21_X1  g473(.A(G868), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n899), .B1(G868), .B2(new_n827), .ZN(G295));
  OAI21_X1  g475(.A(new_n899), .B1(G868), .B2(new_n827), .ZN(G331));
  INV_X1    g476(.A(KEYINPUT44), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n543), .A2(new_n544), .A3(KEYINPUT109), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(G168), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(KEYINPUT110), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT110), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n903), .A2(G168), .A3(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n831), .A2(new_n905), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n905), .A2(new_n907), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n909), .A2(new_n830), .A3(new_n828), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g486(.A1(G171), .A2(KEYINPUT109), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n908), .A2(new_n910), .A3(new_n912), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(new_n885), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n914), .A2(new_n888), .A3(new_n915), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n917), .A2(KEYINPUT113), .A3(new_n918), .ZN(new_n919));
  OAI211_X1 g494(.A(new_n919), .B(new_n896), .C1(KEYINPUT113), .C2(new_n917), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT43), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT111), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n918), .A2(new_n922), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n914), .A2(KEYINPUT111), .A3(new_n888), .A4(new_n915), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n923), .A2(new_n917), .A3(new_n895), .A4(new_n924), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n920), .A2(new_n921), .A3(new_n877), .A4(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n923), .A2(new_n924), .A3(new_n917), .ZN(new_n927));
  AOI21_X1  g502(.A(G37), .B1(new_n927), .B2(new_n896), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n921), .B1(new_n928), .B2(new_n925), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT112), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n926), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  AOI211_X1 g506(.A(KEYINPUT112), .B(new_n921), .C1(new_n928), .C2(new_n925), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n902), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  AND4_X1   g508(.A1(KEYINPUT43), .A2(new_n920), .A3(new_n877), .A4(new_n925), .ZN(new_n934));
  AOI21_X1  g509(.A(KEYINPUT43), .B1(new_n928), .B2(new_n925), .ZN(new_n935));
  OAI21_X1  g510(.A(KEYINPUT44), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n933), .A2(new_n936), .ZN(G397));
  INV_X1    g512(.A(G1384), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n938), .B1(new_n861), .B2(new_n513), .ZN(new_n939));
  XNOR2_X1  g514(.A(KEYINPUT114), .B(KEYINPUT45), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  AND3_X1   g516(.A1(new_n472), .A2(G40), .A3(new_n481), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  NOR3_X1   g518(.A1(new_n941), .A2(G1996), .A3(new_n943), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n944), .B(KEYINPUT115), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n941), .A2(new_n943), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(G2067), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n757), .B(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n950), .B1(new_n735), .B2(G1996), .ZN(new_n951));
  OAI22_X1  g526(.A1(new_n945), .A2(new_n735), .B1(new_n947), .B2(new_n951), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n805), .B(new_n808), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n947), .A2(new_n953), .ZN(new_n954));
  OR2_X1    g529(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  XNOR2_X1  g530(.A(G290), .B(G1986), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n955), .B1(new_n946), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n942), .A2(new_n716), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT50), .ZN(new_n959));
  OAI211_X1 g534(.A(new_n959), .B(new_n938), .C1(new_n861), .C2(new_n513), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n515), .A2(new_n516), .ZN(new_n961));
  AOI21_X1  g536(.A(KEYINPUT71), .B1(new_n503), .B2(KEYINPUT4), .ZN(new_n962));
  AOI211_X1 g537(.A(new_n491), .B(new_n494), .C1(new_n501), .C2(new_n502), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n507), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(G1384), .B1(new_n961), .B2(new_n964), .ZN(new_n965));
  OAI211_X1 g540(.A(KEYINPUT117), .B(new_n960), .C1(new_n965), .C2(new_n959), .ZN(new_n966));
  INV_X1    g541(.A(new_n513), .ZN(new_n967));
  AOI21_X1  g542(.A(G1384), .B1(new_n964), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT117), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n968), .A2(new_n969), .A3(new_n959), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n958), .B1(new_n966), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(new_n748), .ZN(new_n972));
  INV_X1    g547(.A(new_n940), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n943), .B1(new_n965), .B2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT45), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n939), .A2(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n972), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(G286), .B1(new_n971), .B2(new_n977), .ZN(new_n978));
  AND3_X1   g553(.A1(new_n508), .A2(KEYINPUT70), .A3(new_n512), .ZN(new_n979));
  AOI21_X1  g554(.A(KEYINPUT70), .B1(new_n508), .B2(new_n512), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  OAI211_X1 g556(.A(new_n938), .B(new_n973), .C1(new_n981), .C2(new_n861), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n942), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n968), .A2(KEYINPUT45), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n748), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n960), .A2(KEYINPUT117), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n969), .B1(new_n968), .B2(new_n959), .ZN(new_n987));
  OAI21_X1  g562(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n986), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  OAI211_X1 g564(.A(G168), .B(new_n985), .C1(new_n989), .C2(new_n958), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n978), .A2(new_n990), .A3(G8), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(KEYINPUT51), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT51), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n990), .A2(new_n993), .A3(G8), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT53), .ZN(new_n996));
  OAI211_X1 g571(.A(KEYINPUT45), .B(new_n938), .C1(new_n861), .C2(new_n513), .ZN(new_n997));
  OAI211_X1 g572(.A(new_n942), .B(new_n997), .C1(new_n965), .C2(new_n973), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n996), .B1(new_n998), .B2(G2078), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n943), .B1(new_n966), .B2(new_n970), .ZN(new_n1000));
  XOR2_X1   g575(.A(KEYINPUT121), .B(G1961), .Z(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n999), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n996), .A2(G2078), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n997), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(KEYINPUT122), .B1(new_n941), .B2(new_n942), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT122), .ZN(new_n1008));
  AOI211_X1 g583(.A(new_n1008), .B(new_n943), .C1(new_n939), .C2(new_n940), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1005), .B1(new_n1007), .B2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g586(.A(G171), .B1(new_n1003), .B2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n974), .A2(new_n1004), .A3(new_n976), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n999), .B(new_n1013), .C1(new_n1000), .C2(new_n1002), .ZN(new_n1014));
  OAI211_X1 g589(.A(new_n1012), .B(KEYINPUT54), .C1(G171), .C2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n532), .A2(G8), .A3(new_n533), .ZN(new_n1016));
  XNOR2_X1  g591(.A(new_n1016), .B(KEYINPUT55), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  AOI211_X1 g593(.A(G2090), .B(new_n943), .C1(new_n966), .C2(new_n970), .ZN(new_n1019));
  XOR2_X1   g594(.A(KEYINPUT116), .B(G1971), .Z(new_n1020));
  AOI21_X1  g595(.A(new_n943), .B1(new_n968), .B2(KEYINPUT45), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n940), .B1(G164), .B2(G1384), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1020), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  OAI211_X1 g598(.A(new_n1018), .B(G8), .C1(new_n1019), .C2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n789), .A2(G1976), .ZN(new_n1025));
  INV_X1    g600(.A(G1976), .ZN(new_n1026));
  AOI21_X1  g601(.A(KEYINPUT52), .B1(G288), .B2(new_n1026), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n938), .B(new_n942), .C1(new_n861), .C2(new_n513), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1028), .A2(KEYINPUT118), .A3(G8), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(KEYINPUT118), .B1(new_n1028), .B2(G8), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n1025), .B(new_n1027), .C1(new_n1030), .C2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT49), .ZN(new_n1033));
  NOR2_X1   g608(.A1(G305), .A2(G1981), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n786), .B1(new_n573), .B2(new_n574), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1033), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1038));
  NOR3_X1   g613(.A1(new_n1034), .A2(KEYINPUT49), .A3(new_n1036), .ZN(new_n1039));
  OAI22_X1  g614(.A1(new_n1030), .A2(new_n1031), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1032), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT52), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1028), .A2(G8), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT118), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(new_n1029), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1042), .B1(new_n1046), .B2(new_n1025), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1041), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n965), .A2(new_n959), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n939), .A2(KEYINPUT50), .ZN(new_n1050));
  AND4_X1   g625(.A1(new_n679), .A2(new_n1049), .A3(new_n942), .A4(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(G8), .B1(new_n1051), .B2(new_n1023), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(new_n1017), .ZN(new_n1053));
  AND3_X1   g628(.A1(new_n1024), .A2(new_n1048), .A3(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n995), .A2(new_n1015), .A3(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1014), .A2(G171), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1001), .B1(new_n989), .B2(new_n943), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n997), .B(new_n1004), .C1(new_n1006), .C2(new_n1009), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1057), .A2(G301), .A3(new_n999), .A4(new_n1058), .ZN(new_n1059));
  AND3_X1   g634(.A1(new_n1056), .A2(new_n1059), .A3(KEYINPUT123), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT54), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1061), .B1(new_n1059), .B2(KEYINPUT123), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g638(.A(KEYINPUT124), .B1(new_n1055), .B2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1024), .A2(new_n1048), .A3(new_n1053), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1065), .B1(new_n992), .B2(new_n994), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT124), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1056), .A2(new_n1059), .A3(KEYINPUT123), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1003), .A2(new_n1011), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT123), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1069), .A2(new_n1070), .A3(G301), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1068), .A2(new_n1071), .A3(new_n1061), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1066), .A2(new_n1067), .A3(new_n1072), .A4(new_n1015), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1049), .A2(new_n942), .A3(new_n1050), .ZN(new_n1074));
  INV_X1    g649(.A(G1956), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  XNOR2_X1  g651(.A(KEYINPUT56), .B(G2072), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1021), .A2(new_n1022), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT119), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT57), .ZN(new_n1080));
  OAI21_X1  g655(.A(G299), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1082));
  XNOR2_X1  g657(.A(new_n1081), .B(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1076), .A2(new_n1078), .A3(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(new_n589), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n697), .B1(new_n989), .B2(new_n943), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n968), .A2(new_n948), .A3(new_n942), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1085), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1083), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1084), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1089), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(new_n1084), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT61), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  XOR2_X1   g669(.A(KEYINPUT58), .B(G1341), .Z(new_n1095));
  NAND2_X1  g670(.A1(new_n1028), .A2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1096), .B1(new_n998), .B2(G1996), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(new_n553), .ZN(new_n1098));
  NAND2_X1  g673(.A1(KEYINPUT120), .A2(KEYINPUT59), .ZN(new_n1099));
  XOR2_X1   g674(.A(new_n1098), .B(new_n1099), .Z(new_n1100));
  NAND3_X1  g675(.A1(new_n1091), .A2(KEYINPUT61), .A3(new_n1084), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1094), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT60), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1085), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1086), .A2(KEYINPUT60), .A3(new_n589), .A4(new_n1087), .ZN(new_n1107));
  AND3_X1   g682(.A1(new_n1105), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1090), .B1(new_n1102), .B2(new_n1108), .ZN(new_n1109));
  AND3_X1   g684(.A1(new_n1064), .A2(new_n1073), .A3(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1040), .A2(new_n1026), .A3(new_n789), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(new_n1035), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(new_n1046), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1048), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1113), .B1(new_n1114), .B2(new_n1024), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT63), .ZN(new_n1116));
  OAI211_X1 g691(.A(G8), .B(G168), .C1(new_n971), .C2(new_n977), .ZN(new_n1117));
  OAI21_X1  g692(.A(G8), .B1(new_n1019), .B2(new_n1023), .ZN(new_n1118));
  AOI211_X1 g693(.A(new_n1116), .B(new_n1117), .C1(new_n1118), .C2(new_n1017), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1119), .A2(new_n1024), .A3(new_n1048), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1116), .B1(new_n1065), .B2(new_n1117), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1115), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1065), .A2(new_n1056), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT62), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n992), .A2(new_n1124), .A3(new_n994), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1123), .A2(new_n1125), .A3(KEYINPUT125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n995), .A2(KEYINPUT62), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(KEYINPUT125), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1122), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n957), .B1(new_n1110), .B2(new_n1130), .ZN(new_n1131));
  XNOR2_X1  g706(.A(new_n945), .B(KEYINPUT46), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n946), .B1(new_n735), .B2(new_n950), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT126), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1132), .A2(KEYINPUT126), .A3(new_n1133), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1136), .A2(KEYINPUT47), .A3(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n955), .A2(KEYINPUT127), .ZN(new_n1139));
  OR3_X1    g714(.A1(new_n952), .A2(KEYINPUT127), .A3(new_n954), .ZN(new_n1140));
  NOR3_X1   g715(.A1(new_n947), .A2(G1986), .A3(G290), .ZN(new_n1141));
  XOR2_X1   g716(.A(new_n1141), .B(KEYINPUT48), .Z(new_n1142));
  NAND3_X1  g717(.A1(new_n1139), .A2(new_n1140), .A3(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1138), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(new_n806), .ZN(new_n1145));
  NOR3_X1   g720(.A1(new_n952), .A2(new_n809), .A3(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1146), .B1(new_n948), .B2(new_n840), .ZN(new_n1147));
  NOR3_X1   g722(.A1(new_n1147), .A2(new_n943), .A3(new_n941), .ZN(new_n1148));
  AOI21_X1  g723(.A(KEYINPUT47), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1149));
  NOR3_X1   g724(.A1(new_n1144), .A2(new_n1148), .A3(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1131), .A2(new_n1150), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g726(.A1(new_n931), .A2(new_n932), .ZN(new_n1153));
  NOR4_X1   g727(.A1(G401), .A2(new_n461), .A3(G227), .A4(G229), .ZN(new_n1154));
  OAI21_X1  g728(.A(new_n1154), .B1(new_n878), .B2(new_n873), .ZN(new_n1155));
  NOR2_X1   g729(.A1(new_n1153), .A2(new_n1155), .ZN(G308));
  OAI221_X1 g730(.A(new_n1154), .B1(new_n878), .B2(new_n873), .C1(new_n931), .C2(new_n932), .ZN(G225));
endmodule


