//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 0 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 0 1 0 0 1 0 0 1 0 1 0 0 0 1 1 0 1 1 0 1 1 0 1 1 0 0 1 1 1 1 1 0 1 1 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:00 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1250, new_n1251,
    new_n1252;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  XOR2_X1   g0005(.A(KEYINPUT65), .B(G238), .Z(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  XNOR2_X1  g0007(.A(KEYINPUT66), .B(G244), .ZN(new_n208));
  AOI22_X1  g0008(.A1(new_n207), .A2(G68), .B1(G77), .B2(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G50), .A2(G226), .B1(G107), .B2(G264), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G116), .A2(G270), .ZN(new_n212));
  AND3_X1   g0012(.A1(new_n210), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(G232), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n209), .B(new_n213), .C1(new_n201), .C2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G20), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  XOR2_X1   g0017(.A(new_n217), .B(KEYINPUT1), .Z(new_n218));
  NAND2_X1  g0018(.A1(new_n203), .A2(G50), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G13), .ZN(new_n221));
  INV_X1    g0021(.A(new_n221), .ZN(new_n222));
  NAND3_X1  g0022(.A1(new_n220), .A2(G20), .A3(new_n222), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n216), .A2(G13), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n224), .B(G250), .C1(G257), .C2(G264), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT64), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT0), .ZN(new_n227));
  NAND3_X1  g0027(.A1(new_n218), .A2(new_n223), .A3(new_n227), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(new_n214), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT2), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G264), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n235), .B(G270), .Z(new_n236));
  XOR2_X1   g0036(.A(new_n233), .B(new_n236), .Z(G358));
  XNOR2_X1  g0037(.A(G50), .B(G68), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT67), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G58), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G77), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G87), .B(G97), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G107), .ZN(new_n243));
  INV_X1    g0043(.A(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n241), .B(new_n245), .ZN(G351));
  INV_X1    g0046(.A(KEYINPUT13), .ZN(new_n247));
  OR2_X1    g0047(.A1(KEYINPUT3), .A2(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(KEYINPUT3), .A2(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G1698), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n250), .A2(G226), .A3(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(G33), .A2(G97), .ZN(new_n253));
  AND2_X1   g0053(.A1(KEYINPUT3), .A2(G33), .ZN(new_n254));
  NOR2_X1   g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  OAI211_X1 g0055(.A(G232), .B(G1698), .C1(new_n254), .C2(new_n255), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n252), .A2(new_n253), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(KEYINPUT74), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n221), .B1(G33), .B2(G41), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT74), .ZN(new_n260));
  NAND4_X1  g0060(.A1(new_n252), .A2(new_n260), .A3(new_n253), .A4(new_n256), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n258), .A2(new_n259), .A3(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G41), .ZN(new_n263));
  INV_X1    g0063(.A(G45), .ZN(new_n264));
  AOI21_X1  g0064(.A(G1), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT68), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n265), .A2(new_n266), .A3(G274), .ZN(new_n267));
  INV_X1    g0067(.A(G1), .ZN(new_n268));
  OAI211_X1 g0068(.A(new_n268), .B(G274), .C1(G41), .C2(G45), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(KEYINPUT68), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n267), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(KEYINPUT75), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT75), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n267), .A2(new_n273), .A3(new_n270), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n259), .A2(new_n265), .ZN(new_n275));
  AOI22_X1  g0075(.A1(new_n272), .A2(new_n274), .B1(G238), .B2(new_n275), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n247), .B1(new_n262), .B2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n262), .A2(new_n276), .A3(new_n247), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n278), .A2(G190), .A3(new_n279), .ZN(new_n280));
  AND3_X1   g0080(.A1(new_n262), .A2(new_n276), .A3(new_n247), .ZN(new_n281));
  OAI21_X1  g0081(.A(G200), .B1(new_n281), .B2(new_n277), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n202), .A2(G20), .ZN(new_n283));
  INV_X1    g0083(.A(G20), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G33), .ZN(new_n285));
  INV_X1    g0085(.A(G77), .ZN(new_n286));
  NOR2_X1   g0086(.A1(G20), .A2(G33), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G50), .ZN(new_n289));
  OAI221_X1 g0089(.A(new_n283), .B1(new_n285), .B2(new_n286), .C1(new_n288), .C2(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(new_n221), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n290), .A2(KEYINPUT11), .A3(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n292), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n294), .B1(G1), .B2(new_n284), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n293), .B1(new_n202), .B2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G13), .ZN(new_n297));
  NOR3_X1   g0097(.A1(new_n297), .A2(new_n284), .A3(G1), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(new_n202), .ZN(new_n299));
  XOR2_X1   g0099(.A(new_n299), .B(KEYINPUT12), .Z(new_n300));
  AOI21_X1  g0100(.A(KEYINPUT11), .B1(new_n290), .B2(new_n292), .ZN(new_n301));
  NOR3_X1   g0101(.A1(new_n296), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n280), .A2(new_n282), .A3(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(G169), .B1(new_n281), .B2(new_n277), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(KEYINPUT14), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n278), .A2(G179), .A3(new_n279), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT14), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n308), .B(G169), .C1(new_n281), .C2(new_n277), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n306), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n302), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n304), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  XNOR2_X1  g0112(.A(KEYINPUT8), .B(G58), .ZN(new_n313));
  INV_X1    g0113(.A(G150), .ZN(new_n314));
  OAI22_X1  g0114(.A1(new_n313), .A2(new_n285), .B1(new_n314), .B2(new_n288), .ZN(new_n315));
  XNOR2_X1  g0115(.A(new_n315), .B(KEYINPUT70), .ZN(new_n316));
  OAI21_X1  g0116(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AOI22_X1  g0118(.A1(new_n318), .A2(new_n292), .B1(new_n289), .B2(new_n298), .ZN(new_n319));
  OR2_X1    g0119(.A1(new_n295), .A2(new_n289), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(G1698), .B1(new_n248), .B2(new_n249), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(G222), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n254), .A2(new_n255), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(G77), .ZN(new_n325));
  INV_X1    g0125(.A(G223), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n250), .A2(G1698), .ZN(new_n327));
  OAI211_X1 g0127(.A(new_n323), .B(new_n325), .C1(new_n326), .C2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT69), .ZN(new_n329));
  OR2_X1    g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(new_n329), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n330), .A2(new_n259), .A3(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n271), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n333), .B1(G226), .B2(new_n275), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n321), .B1(new_n335), .B2(G179), .ZN(new_n336));
  AOI21_X1  g0136(.A(G169), .B1(new_n332), .B2(new_n334), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT9), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n321), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n335), .A2(G200), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n319), .A2(KEYINPUT9), .A3(new_n320), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n332), .A2(G190), .A3(new_n334), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n340), .A2(new_n341), .A3(new_n342), .A4(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(KEYINPUT10), .ZN(new_n345));
  AOI22_X1  g0145(.A1(new_n321), .A2(new_n339), .B1(new_n335), .B2(G200), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT10), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n346), .A2(new_n347), .A3(new_n342), .A4(new_n343), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n338), .B1(new_n345), .B2(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n333), .B1(new_n208), .B2(new_n275), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n250), .A2(G232), .A3(new_n251), .ZN(new_n351));
  INV_X1    g0151(.A(G107), .ZN(new_n352));
  OAI221_X1 g0152(.A(new_n351), .B1(new_n352), .B2(new_n250), .C1(new_n327), .C2(new_n206), .ZN(new_n353));
  XNOR2_X1  g0153(.A(new_n353), .B(KEYINPUT71), .ZN(new_n354));
  INV_X1    g0154(.A(new_n259), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n350), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(G169), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  OAI22_X1  g0158(.A1(new_n313), .A2(new_n288), .B1(new_n284), .B2(new_n286), .ZN(new_n359));
  XNOR2_X1  g0159(.A(KEYINPUT15), .B(G87), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n360), .A2(new_n285), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n292), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n298), .A2(new_n286), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n362), .B(new_n363), .C1(new_n286), .C2(new_n295), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n358), .B(new_n364), .C1(G179), .C2(new_n356), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n356), .A2(G200), .B1(KEYINPUT72), .B2(new_n364), .ZN(new_n366));
  INV_X1    g0166(.A(G190), .ZN(new_n367));
  OAI221_X1 g0167(.A(new_n366), .B1(KEYINPUT72), .B2(new_n364), .C1(new_n367), .C2(new_n356), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n349), .A2(new_n365), .A3(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT73), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n349), .A2(KEYINPUT73), .A3(new_n365), .A4(new_n368), .ZN(new_n372));
  AOI21_X1  g0172(.A(KEYINPUT7), .B1(new_n324), .B2(new_n284), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT7), .ZN(new_n374));
  NOR4_X1   g0174(.A1(new_n254), .A2(new_n255), .A3(new_n374), .A4(G20), .ZN(new_n375));
  OAI21_X1  g0175(.A(G68), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(G159), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n288), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(G58), .A2(G68), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n284), .B1(new_n203), .B2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n376), .A2(new_n379), .A3(new_n382), .ZN(new_n383));
  AND3_X1   g0183(.A1(new_n383), .A2(KEYINPUT76), .A3(KEYINPUT16), .ZN(new_n384));
  AOI21_X1  g0184(.A(KEYINPUT16), .B1(new_n383), .B2(KEYINPUT76), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n292), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n295), .A2(new_n313), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n313), .ZN(new_n389));
  INV_X1    g0189(.A(new_n298), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n386), .A2(new_n388), .A3(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(G179), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n275), .A2(G232), .B1(new_n267), .B2(new_n270), .ZN(new_n395));
  OAI211_X1 g0195(.A(G226), .B(G1698), .C1(new_n254), .C2(new_n255), .ZN(new_n396));
  OAI211_X1 g0196(.A(G223), .B(new_n251), .C1(new_n254), .C2(new_n255), .ZN(new_n397));
  NAND2_X1  g0197(.A1(G33), .A2(G87), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n399), .A2(KEYINPUT77), .A3(new_n259), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(KEYINPUT77), .B1(new_n399), .B2(new_n259), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n394), .B(new_n395), .C1(new_n401), .C2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n399), .A2(new_n259), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(new_n395), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n357), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n403), .A2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n393), .A2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT18), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n393), .A2(KEYINPUT18), .A3(new_n408), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n367), .B(new_n395), .C1(new_n401), .C2(new_n402), .ZN(new_n413));
  INV_X1    g0213(.A(G200), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n405), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n386), .A2(new_n388), .A3(new_n392), .A4(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(KEYINPUT17), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT16), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n248), .A2(new_n284), .A3(new_n249), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n374), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n248), .A2(KEYINPUT7), .A3(new_n284), .A4(new_n249), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n202), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NOR3_X1   g0223(.A1(new_n423), .A2(new_n378), .A3(new_n381), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT76), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n419), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n383), .A2(KEYINPUT76), .A3(KEYINPUT16), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n391), .B1(new_n428), .B2(new_n292), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT17), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n429), .A2(new_n430), .A3(new_n388), .A4(new_n416), .ZN(new_n431));
  AOI22_X1  g0231(.A1(new_n411), .A2(new_n412), .B1(new_n418), .B2(new_n431), .ZN(new_n432));
  AND4_X1   g0232(.A1(new_n312), .A2(new_n371), .A3(new_n372), .A4(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT4), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n322), .A2(new_n434), .A3(G244), .ZN(new_n435));
  OAI211_X1 g0235(.A(G244), .B(new_n251), .C1(new_n254), .C2(new_n255), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(KEYINPUT4), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n250), .A2(G250), .A3(G1698), .ZN(new_n439));
  NAND2_X1  g0239(.A1(G33), .A2(G283), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT79), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n438), .A2(KEYINPUT79), .A3(new_n439), .A4(new_n440), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n443), .A2(new_n259), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n268), .A2(G45), .ZN(new_n446));
  OR2_X1    g0246(.A1(KEYINPUT5), .A2(G41), .ZN(new_n447));
  NAND2_X1  g0247(.A1(KEYINPUT5), .A2(G41), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n446), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n449), .A2(new_n259), .ZN(new_n450));
  AOI22_X1  g0250(.A1(new_n450), .A2(G257), .B1(G274), .B2(new_n449), .ZN(new_n451));
  XNOR2_X1  g0251(.A(new_n451), .B(KEYINPUT80), .ZN(new_n452));
  AND2_X1   g0252(.A1(new_n445), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n352), .A2(KEYINPUT6), .A3(G97), .ZN(new_n454));
  INV_X1    g0254(.A(G97), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n455), .A2(new_n352), .ZN(new_n456));
  NOR2_X1   g0256(.A1(G97), .A2(G107), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n454), .B1(new_n458), .B2(KEYINPUT6), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(G20), .ZN(new_n460));
  OAI21_X1  g0260(.A(G107), .B1(new_n373), .B2(new_n375), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n287), .A2(G77), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(new_n292), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n298), .A2(new_n455), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n268), .A2(G33), .ZN(new_n466));
  AND3_X1   g0266(.A1(new_n390), .A2(new_n294), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(G97), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n464), .A2(new_n465), .A3(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT78), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n464), .A2(KEYINPUT78), .A3(new_n465), .A4(new_n468), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n453), .A2(G190), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n445), .A2(new_n452), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(G200), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n445), .A2(new_n452), .A3(G179), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n476), .B1(new_n453), .B2(new_n357), .ZN(new_n477));
  XNOR2_X1  g0277(.A(new_n469), .B(KEYINPUT81), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n473), .A2(new_n475), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n284), .A2(G33), .A3(G116), .ZN(new_n480));
  XNOR2_X1  g0280(.A(new_n480), .B(KEYINPUT87), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n250), .A2(new_n284), .A3(G87), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(KEYINPUT22), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT22), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n250), .A2(new_n484), .A3(new_n284), .A4(G87), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n481), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT24), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n284), .A2(G107), .ZN(new_n488));
  XNOR2_X1  g0288(.A(new_n488), .B(KEYINPUT23), .ZN(new_n489));
  AND3_X1   g0289(.A1(new_n486), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n487), .B1(new_n486), .B2(new_n489), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n292), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n467), .A2(G107), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n298), .A2(new_n352), .ZN(new_n494));
  XOR2_X1   g0294(.A(new_n494), .B(KEYINPUT25), .Z(new_n495));
  NAND3_X1  g0295(.A1(new_n492), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  OAI211_X1 g0297(.A(G257), .B(G1698), .C1(new_n254), .C2(new_n255), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT88), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n322), .A2(G250), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n250), .A2(KEYINPUT88), .A3(G257), .A4(G1698), .ZN(new_n502));
  NAND2_X1  g0302(.A1(G33), .A2(G294), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n500), .A2(new_n501), .A3(new_n502), .A4(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n259), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n450), .A2(G264), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n507), .B1(G274), .B2(new_n449), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(G190), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n497), .B(new_n509), .C1(new_n414), .C2(new_n508), .ZN(new_n510));
  AND2_X1   g0310(.A1(new_n505), .A2(new_n506), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n449), .A2(G274), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(new_n357), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n508), .A2(new_n394), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n496), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  AND3_X1   g0316(.A1(new_n479), .A2(new_n510), .A3(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT19), .ZN(new_n518));
  INV_X1    g0318(.A(G87), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n457), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n253), .A2(new_n284), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n518), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NOR3_X1   g0322(.A1(new_n253), .A2(KEYINPUT19), .A3(G20), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n250), .A2(new_n284), .ZN(new_n524));
  OAI22_X1  g0324(.A1(new_n522), .A2(new_n523), .B1(new_n524), .B2(new_n202), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(KEYINPUT83), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT83), .ZN(new_n527));
  OAI221_X1 g0327(.A(new_n527), .B1(new_n524), .B2(new_n202), .C1(new_n522), .C2(new_n523), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n526), .A2(new_n528), .A3(new_n292), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n360), .A2(new_n298), .ZN(new_n530));
  INV_X1    g0330(.A(new_n467), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n529), .B(new_n530), .C1(new_n360), .C2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n322), .A2(G238), .ZN(new_n533));
  NAND2_X1  g0333(.A1(G33), .A2(G116), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n250), .A2(G244), .A3(G1698), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n259), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n355), .A2(G250), .A3(new_n446), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT82), .ZN(new_n539));
  INV_X1    g0339(.A(G274), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n539), .B1(new_n446), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n355), .A2(new_n539), .A3(G250), .A4(new_n446), .ZN(new_n543));
  AND3_X1   g0343(.A1(new_n537), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n394), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n532), .A2(new_n545), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n544), .A2(G169), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n544), .A2(new_n414), .ZN(new_n548));
  AND2_X1   g0348(.A1(new_n542), .A2(new_n543), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n549), .A2(G190), .A3(new_n537), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n467), .A2(G87), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n550), .A2(new_n529), .A3(new_n530), .A4(new_n551), .ZN(new_n552));
  OAI22_X1  g0352(.A1(new_n546), .A2(new_n547), .B1(new_n548), .B2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n447), .A2(new_n448), .ZN(new_n555));
  INV_X1    g0355(.A(new_n446), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n557), .A2(new_n355), .A3(G270), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n512), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(KEYINPUT84), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n322), .A2(G257), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n250), .A2(G264), .A3(G1698), .ZN(new_n562));
  INV_X1    g0362(.A(G303), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n561), .B(new_n562), .C1(new_n563), .C2(new_n250), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n259), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT84), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n558), .A2(new_n566), .A3(new_n512), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n560), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n467), .A2(G116), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n298), .A2(new_n244), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n440), .B(new_n284), .C1(G33), .C2(new_n455), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n571), .B(new_n292), .C1(new_n284), .C2(G116), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT20), .ZN(new_n573));
  AND2_X1   g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n572), .A2(new_n573), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n569), .B(new_n570), .C1(new_n574), .C2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n568), .A2(G169), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(KEYINPUT85), .A2(KEYINPUT21), .ZN(new_n578));
  OR2_X1    g0378(.A1(KEYINPUT85), .A2(KEYINPUT21), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT86), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n577), .A2(KEYINPUT86), .A3(new_n578), .A4(new_n579), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n568), .A2(KEYINPUT21), .A3(G169), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n560), .A2(new_n565), .A3(G179), .A4(new_n567), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n576), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n568), .A2(G200), .ZN(new_n589));
  INV_X1    g0389(.A(new_n576), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n589), .B(new_n590), .C1(new_n367), .C2(new_n568), .ZN(new_n591));
  AND4_X1   g0391(.A1(new_n554), .A2(new_n584), .A3(new_n588), .A4(new_n591), .ZN(new_n592));
  AND3_X1   g0392(.A1(new_n433), .A2(new_n517), .A3(new_n592), .ZN(G372));
  NAND3_X1  g0393(.A1(new_n584), .A2(new_n516), .A3(new_n588), .ZN(new_n594));
  INV_X1    g0394(.A(new_n552), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT89), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n537), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n536), .A2(KEYINPUT89), .A3(new_n259), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n414), .B1(new_n599), .B2(new_n549), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n595), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n479), .A2(new_n594), .A3(new_n510), .A4(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT26), .ZN(new_n604));
  AND2_X1   g0404(.A1(new_n471), .A2(new_n472), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n477), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(G169), .B1(new_n599), .B2(new_n549), .ZN(new_n607));
  OAI22_X1  g0407(.A1(new_n546), .A2(new_n607), .B1(new_n552), .B2(new_n600), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n604), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  XOR2_X1   g0409(.A(KEYINPUT90), .B(KEYINPUT26), .Z(new_n610));
  NAND4_X1  g0410(.A1(new_n554), .A2(new_n477), .A3(new_n478), .A4(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  AND2_X1   g0412(.A1(new_n532), .A2(new_n545), .ZN(new_n613));
  INV_X1    g0413(.A(new_n607), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n603), .A2(new_n612), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n433), .A2(new_n616), .ZN(new_n617));
  AND2_X1   g0417(.A1(new_n418), .A2(new_n431), .ZN(new_n618));
  OR2_X1    g0418(.A1(new_n618), .A2(new_n304), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n310), .A2(new_n311), .ZN(new_n620));
  AND2_X1   g0420(.A1(new_n620), .A2(new_n365), .ZN(new_n621));
  AOI21_X1  g0421(.A(KEYINPUT18), .B1(new_n393), .B2(new_n408), .ZN(new_n622));
  AND3_X1   g0422(.A1(new_n393), .A2(KEYINPUT18), .A3(new_n408), .ZN(new_n623));
  OAI22_X1  g0423(.A1(new_n619), .A2(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n345), .A2(new_n348), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n338), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n617), .A2(new_n626), .ZN(G369));
  NOR2_X1   g0427(.A1(new_n297), .A2(G20), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n268), .ZN(new_n629));
  OR2_X1    g0429(.A1(new_n629), .A2(KEYINPUT27), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(KEYINPUT27), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n630), .A2(G213), .A3(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(G343), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n516), .A2(new_n635), .ZN(new_n636));
  XOR2_X1   g0436(.A(new_n636), .B(KEYINPUT91), .Z(new_n637));
  OAI211_X1 g0437(.A(new_n510), .B(new_n516), .C1(new_n497), .C2(new_n635), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT92), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n637), .A2(KEYINPUT92), .A3(new_n638), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n584), .A2(new_n588), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n576), .A2(new_n634), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n645), .A2(new_n591), .A3(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n647), .B1(new_n645), .B2(new_n646), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(G330), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n644), .A2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n645), .A2(new_n634), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n653), .B1(new_n641), .B2(new_n642), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n516), .A2(new_n634), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n651), .A2(new_n656), .ZN(G399));
  INV_X1    g0457(.A(new_n224), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n658), .A2(G41), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n520), .A2(G116), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n660), .A2(G1), .A3(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n662), .B1(new_n219), .B2(new_n660), .ZN(new_n663));
  XNOR2_X1  g0463(.A(new_n663), .B(KEYINPUT28), .ZN(new_n664));
  AOI21_X1  g0464(.A(KEYINPUT29), .B1(new_n616), .B2(new_n635), .ZN(new_n665));
  OR2_X1    g0465(.A1(new_n665), .A2(KEYINPUT94), .ZN(new_n666));
  INV_X1    g0466(.A(new_n610), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n477), .A2(new_n478), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n667), .B1(new_n668), .B2(new_n553), .ZN(new_n669));
  AOI22_X1  g0469(.A1(new_n613), .A2(new_n614), .B1(new_n595), .B2(new_n601), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n670), .A2(KEYINPUT26), .A3(new_n477), .A4(new_n605), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n603), .A2(new_n672), .A3(new_n615), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n673), .A2(KEYINPUT29), .A3(new_n635), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n665), .A2(KEYINPUT94), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n666), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n549), .A2(new_n537), .ZN(new_n677));
  NOR3_X1   g0477(.A1(new_n586), .A2(new_n677), .A3(new_n507), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n453), .A2(KEYINPUT30), .A3(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT30), .ZN(new_n680));
  AND3_X1   g0480(.A1(new_n560), .A2(new_n565), .A3(new_n567), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n681), .A2(new_n511), .A3(G179), .A4(new_n544), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n680), .B1(new_n682), .B2(new_n474), .ZN(new_n683));
  AOI21_X1  g0483(.A(G179), .B1(new_n599), .B2(new_n549), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n474), .A2(new_n684), .A3(new_n513), .A4(new_n568), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n679), .A2(new_n683), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(new_n634), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT31), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n686), .A2(KEYINPUT31), .A3(new_n634), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT93), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n517), .A2(new_n592), .A3(new_n635), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n689), .A2(KEYINPUT93), .A3(new_n690), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n693), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(G330), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n676), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n664), .B1(new_n699), .B2(G1), .ZN(G364));
  INV_X1    g0500(.A(new_n649), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n268), .B1(new_n628), .B2(G45), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n659), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n705), .B1(G330), .B2(new_n648), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n658), .A2(new_n250), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n220), .A2(new_n264), .ZN(new_n708));
  OAI211_X1 g0508(.A(new_n707), .B(new_n708), .C1(new_n241), .C2(new_n264), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n250), .A2(G355), .A3(new_n224), .ZN(new_n710));
  OAI211_X1 g0510(.A(new_n709), .B(new_n710), .C1(G116), .C2(new_n224), .ZN(new_n711));
  NOR2_X1   g0511(.A1(G13), .A2(G33), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n713), .A2(G20), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n221), .B1(G20), .B2(new_n357), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n284), .A2(G179), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n414), .A2(G190), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(G190), .A2(G200), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n717), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  AOI22_X1  g0523(.A1(new_n720), .A2(G283), .B1(new_n723), .B2(G329), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n284), .A2(new_n394), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(new_n718), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(G317), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(KEYINPUT33), .ZN(new_n729));
  OR2_X1    g0529(.A1(new_n728), .A2(KEYINPUT33), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n727), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n724), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n725), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n733), .A2(new_n367), .A3(G200), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(G322), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n324), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n367), .A2(new_n414), .ZN(new_n738));
  AND2_X1   g0538(.A1(new_n738), .A2(new_n717), .ZN(new_n739));
  OR2_X1    g0539(.A1(new_n739), .A2(KEYINPUT95), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(KEYINPUT95), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  AOI211_X1 g0543(.A(new_n732), .B(new_n737), .C1(new_n743), .C2(G303), .ZN(new_n744));
  NOR3_X1   g0544(.A1(new_n367), .A2(G179), .A3(G200), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(new_n284), .ZN(new_n746));
  INV_X1    g0546(.A(G294), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n725), .A2(new_n738), .ZN(new_n748));
  INV_X1    g0548(.A(G326), .ZN(new_n749));
  OAI22_X1  g0549(.A1(new_n746), .A2(new_n747), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  XOR2_X1   g0550(.A(new_n750), .B(KEYINPUT96), .Z(new_n751));
  INV_X1    g0551(.A(G311), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n725), .A2(new_n721), .ZN(new_n753));
  OAI211_X1 g0553(.A(new_n744), .B(new_n751), .C1(new_n752), .C2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n748), .ZN(new_n755));
  AOI22_X1  g0555(.A1(G50), .A2(new_n755), .B1(new_n720), .B2(G107), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n756), .B1(new_n286), .B2(new_n753), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n757), .B1(G87), .B2(new_n743), .ZN(new_n758));
  OAI21_X1  g0558(.A(KEYINPUT32), .B1(new_n722), .B2(new_n377), .ZN(new_n759));
  OR3_X1    g0559(.A1(new_n722), .A2(KEYINPUT32), .A3(new_n377), .ZN(new_n760));
  OAI211_X1 g0560(.A(new_n759), .B(new_n760), .C1(new_n735), .C2(new_n201), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n746), .A2(new_n455), .ZN(new_n762));
  NOR3_X1   g0562(.A1(new_n761), .A2(new_n324), .A3(new_n762), .ZN(new_n763));
  OAI211_X1 g0563(.A(new_n758), .B(new_n763), .C1(new_n202), .C2(new_n726), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n754), .A2(new_n764), .ZN(new_n765));
  AOI22_X1  g0565(.A1(new_n711), .A2(new_n716), .B1(new_n715), .B2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n714), .ZN(new_n767));
  OAI211_X1 g0567(.A(new_n704), .B(new_n766), .C1(new_n648), .C2(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n706), .A2(new_n768), .ZN(G396));
  NOR2_X1   g0569(.A1(new_n365), .A2(new_n634), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n364), .A2(new_n634), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n368), .A2(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n770), .B1(new_n772), .B2(new_n365), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n616), .A2(new_n635), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(KEYINPUT100), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n773), .B1(new_n616), .B2(new_n635), .ZN(new_n776));
  XOR2_X1   g0576(.A(new_n775), .B(new_n776), .Z(new_n777));
  XOR2_X1   g0577(.A(new_n777), .B(new_n697), .Z(new_n778));
  INV_X1    g0578(.A(new_n704), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n324), .B1(new_n723), .B2(G132), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n781), .B1(new_n742), .B2(new_n289), .ZN(new_n782));
  AOI22_X1  g0582(.A1(G137), .A2(new_n755), .B1(new_n727), .B2(G150), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n783), .B1(new_n377), .B2(new_n753), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n784), .B1(G143), .B2(new_n734), .ZN(new_n785));
  XOR2_X1   g0585(.A(new_n785), .B(KEYINPUT34), .Z(new_n786));
  XOR2_X1   g0586(.A(KEYINPUT97), .B(KEYINPUT98), .Z(new_n787));
  AOI21_X1  g0587(.A(new_n782), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n746), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n789), .A2(G58), .B1(new_n720), .B2(G68), .ZN(new_n790));
  OAI211_X1 g0590(.A(new_n788), .B(new_n790), .C1(new_n787), .C2(new_n786), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n722), .A2(new_n752), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n720), .A2(G87), .ZN(new_n793));
  INV_X1    g0593(.A(G283), .ZN(new_n794));
  OAI211_X1 g0594(.A(new_n793), .B(new_n324), .C1(new_n794), .C2(new_n726), .ZN(new_n795));
  AOI211_X1 g0595(.A(new_n762), .B(new_n795), .C1(G303), .C2(new_n755), .ZN(new_n796));
  INV_X1    g0596(.A(new_n753), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n734), .A2(G294), .B1(G116), .B2(new_n797), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n796), .B(new_n798), .C1(new_n352), .C2(new_n742), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n791), .B1(new_n792), .B2(new_n799), .ZN(new_n800));
  XOR2_X1   g0600(.A(new_n800), .B(KEYINPUT99), .Z(new_n801));
  AOI21_X1  g0601(.A(new_n779), .B1(new_n801), .B2(new_n715), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n715), .A2(new_n712), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n802), .B1(G77), .B2(new_n804), .C1(new_n713), .C2(new_n773), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n780), .A2(new_n805), .ZN(G384));
  INV_X1    g0606(.A(KEYINPUT106), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n687), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n686), .A2(KEYINPUT106), .A3(new_n634), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n808), .A2(new_n688), .A3(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(KEYINPUT107), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND4_X1  g0612(.A1(new_n808), .A2(KEYINPUT107), .A3(new_n688), .A4(new_n809), .ZN(new_n813));
  NAND4_X1  g0613(.A1(new_n812), .A2(new_n694), .A3(new_n690), .A4(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n772), .A2(new_n365), .ZN(new_n815));
  INV_X1    g0615(.A(new_n770), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n311), .A2(new_n634), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n620), .A2(new_n303), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(KEYINPUT101), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT101), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n312), .A2(new_n821), .A3(new_n818), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n620), .A2(new_n635), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n817), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n814), .A2(new_n826), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n429), .A2(new_n388), .B1(new_n407), .B2(new_n632), .ZN(new_n828));
  INV_X1    g0628(.A(new_n417), .ZN(new_n829));
  OAI21_X1  g0629(.A(KEYINPUT37), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n632), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n393), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT37), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n409), .A2(new_n832), .A3(new_n833), .A4(new_n417), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n830), .A2(new_n834), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n835), .B1(new_n432), .B2(new_n832), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT38), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n835), .B(KEYINPUT38), .C1(new_n432), .C2(new_n832), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n838), .A2(KEYINPUT104), .A3(new_n839), .ZN(new_n840));
  OR3_X1    g0640(.A1(new_n836), .A2(KEYINPUT104), .A3(new_n837), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT40), .ZN(new_n843));
  NOR3_X1   g0643(.A1(new_n827), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n839), .ZN(new_n845));
  INV_X1    g0645(.A(new_n832), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n623), .A2(new_n622), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n846), .B1(new_n847), .B2(new_n618), .ZN(new_n848));
  AOI21_X1  g0648(.A(KEYINPUT38), .B1(new_n848), .B2(new_n835), .ZN(new_n849));
  OAI21_X1  g0649(.A(KEYINPUT102), .B1(new_n845), .B2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT102), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n838), .A2(new_n851), .A3(new_n839), .ZN(new_n852));
  NAND4_X1  g0652(.A1(new_n850), .A2(new_n852), .A3(new_n814), .A4(new_n826), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(new_n843), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT108), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n853), .A2(KEYINPUT108), .A3(new_n843), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n844), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n433), .A2(new_n814), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n858), .B(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(G330), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n310), .A2(new_n311), .A3(new_n635), .ZN(new_n862));
  XNOR2_X1  g0662(.A(new_n862), .B(KEYINPUT103), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(KEYINPUT39), .B1(new_n840), .B2(new_n841), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT39), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n866), .B1(new_n838), .B2(new_n839), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n864), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n847), .A2(new_n632), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n774), .A2(new_n816), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n819), .A2(KEYINPUT101), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n821), .B1(new_n312), .B2(new_n818), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n825), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n870), .A2(new_n850), .A3(new_n873), .A4(new_n852), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n868), .A2(new_n869), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(KEYINPUT105), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT105), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n868), .A2(new_n877), .A3(new_n869), .A4(new_n874), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g0679(.A(new_n861), .B(new_n879), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n666), .A2(new_n433), .A3(new_n674), .A4(new_n675), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(new_n626), .ZN(new_n882));
  XNOR2_X1  g0682(.A(new_n880), .B(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n883), .B1(new_n268), .B2(new_n628), .ZN(new_n884));
  OAI211_X1 g0684(.A(G20), .B(new_n222), .C1(new_n459), .C2(KEYINPUT35), .ZN(new_n885));
  AOI211_X1 g0685(.A(new_n244), .B(new_n885), .C1(KEYINPUT35), .C2(new_n459), .ZN(new_n886));
  XOR2_X1   g0686(.A(new_n886), .B(KEYINPUT36), .Z(new_n887));
  NAND2_X1  g0687(.A1(new_n380), .A2(G77), .ZN(new_n888));
  OAI22_X1  g0688(.A1(new_n219), .A2(new_n888), .B1(G50), .B2(new_n202), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n889), .A2(G1), .A3(new_n297), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n884), .A2(new_n887), .A3(new_n890), .ZN(G367));
  INV_X1    g0691(.A(KEYINPUT109), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n605), .A2(new_n634), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n479), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n477), .A2(new_n605), .A3(new_n634), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n654), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n892), .B1(new_n897), .B2(KEYINPUT42), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(KEYINPUT42), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT42), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n654), .A2(KEYINPUT109), .A3(new_n900), .A4(new_n896), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n516), .B1(new_n894), .B2(new_n895), .ZN(new_n902));
  INV_X1    g0702(.A(new_n668), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n635), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND4_X1  g0704(.A1(new_n898), .A2(new_n899), .A3(new_n901), .A4(new_n904), .ZN(new_n905));
  AND3_X1   g0705(.A1(new_n529), .A2(new_n530), .A3(new_n551), .ZN(new_n906));
  OR2_X1    g0706(.A1(new_n906), .A2(new_n635), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n670), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n908), .B1(new_n615), .B2(new_n907), .ZN(new_n909));
  OR2_X1    g0709(.A1(new_n909), .A2(KEYINPUT43), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(KEYINPUT43), .ZN(new_n911));
  AND3_X1   g0711(.A1(new_n905), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n910), .B1(new_n905), .B2(new_n911), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n650), .A2(new_n896), .ZN(new_n914));
  OAI22_X1  g0714(.A1(new_n912), .A2(new_n913), .B1(KEYINPUT110), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(KEYINPUT110), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  OR2_X1    g0717(.A1(new_n915), .A2(new_n916), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n659), .B(KEYINPUT41), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT112), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n644), .A2(new_n649), .A3(new_n653), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n701), .B1(new_n643), .B2(new_n652), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n654), .A2(KEYINPUT111), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n924), .B(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n921), .B1(new_n926), .B2(new_n698), .ZN(new_n927));
  INV_X1    g0727(.A(new_n925), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n924), .B(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n929), .A2(KEYINPUT112), .A3(new_n699), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n656), .A2(new_n896), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n931), .A2(KEYINPUT44), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT44), .ZN(new_n933));
  NOR3_X1   g0733(.A1(new_n656), .A2(new_n933), .A3(new_n896), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n656), .A2(new_n896), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT45), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(KEYINPUT45), .B1(new_n656), .B2(new_n896), .ZN(new_n938));
  OAI22_X1  g0738(.A1(new_n932), .A2(new_n934), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n650), .ZN(new_n940));
  OAI221_X1 g0740(.A(new_n651), .B1(new_n937), .B2(new_n938), .C1(new_n932), .C2(new_n934), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n927), .A2(new_n930), .A3(new_n940), .A4(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n920), .B1(new_n942), .B2(new_n699), .ZN(new_n943));
  OAI211_X1 g0743(.A(new_n917), .B(new_n918), .C1(new_n943), .C2(new_n703), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n746), .A2(new_n202), .ZN(new_n945));
  OAI221_X1 g0745(.A(new_n250), .B1(new_n753), .B2(new_n289), .C1(new_n377), .C2(new_n726), .ZN(new_n946));
  AOI211_X1 g0746(.A(new_n945), .B(new_n946), .C1(G143), .C2(new_n755), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n734), .A2(G150), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n743), .A2(G58), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n719), .A2(new_n286), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n950), .B1(G137), .B2(new_n723), .ZN(new_n951));
  NAND4_X1  g0751(.A1(new_n947), .A2(new_n948), .A3(new_n949), .A4(new_n951), .ZN(new_n952));
  OAI22_X1  g0752(.A1(new_n735), .A2(new_n563), .B1(new_n753), .B2(new_n794), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n953), .B1(G294), .B2(new_n727), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n743), .A2(KEYINPUT46), .A3(G116), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT46), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(new_n742), .B2(new_n244), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n748), .A2(new_n752), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n324), .B1(new_n719), .B2(new_n455), .ZN(new_n959));
  AOI211_X1 g0759(.A(new_n958), .B(new_n959), .C1(G107), .C2(new_n789), .ZN(new_n960));
  NAND4_X1  g0760(.A1(new_n954), .A2(new_n955), .A3(new_n957), .A4(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n722), .A2(new_n728), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n952), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT47), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n779), .B1(new_n964), .B2(new_n715), .ZN(new_n965));
  INV_X1    g0765(.A(new_n707), .ZN(new_n966));
  OAI221_X1 g0766(.A(new_n716), .B1(new_n224), .B2(new_n360), .C1(new_n236), .C2(new_n966), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n965), .B(new_n967), .C1(new_n767), .C2(new_n909), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n944), .A2(new_n968), .ZN(G387));
  NAND2_X1  g0769(.A1(new_n927), .A2(new_n930), .ZN(new_n970));
  OAI211_X1 g0770(.A(new_n970), .B(new_n659), .C1(new_n699), .C2(new_n929), .ZN(new_n971));
  OAI22_X1  g0771(.A1(new_n753), .A2(new_n202), .B1(new_n722), .B2(new_n314), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n972), .B1(new_n743), .B2(G77), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n734), .A2(G50), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n755), .A2(G159), .ZN(new_n975));
  OAI221_X1 g0775(.A(new_n250), .B1(new_n719), .B2(new_n455), .C1(new_n313), .C2(new_n726), .ZN(new_n976));
  INV_X1    g0776(.A(new_n360), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n976), .B1(new_n977), .B2(new_n789), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n973), .A2(new_n974), .A3(new_n975), .A4(new_n978), .ZN(new_n979));
  OAI22_X1  g0779(.A1(new_n735), .A2(new_n728), .B1(new_n753), .B2(new_n563), .ZN(new_n980));
  AOI22_X1  g0780(.A1(new_n980), .A2(KEYINPUT113), .B1(G311), .B2(new_n727), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n981), .B1(KEYINPUT113), .B2(new_n980), .C1(new_n736), .C2(new_n748), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT48), .ZN(new_n983));
  OAI221_X1 g0783(.A(new_n983), .B1(new_n794), .B2(new_n746), .C1(new_n747), .C2(new_n742), .ZN(new_n984));
  XOR2_X1   g0784(.A(new_n984), .B(KEYINPUT49), .Z(new_n985));
  OAI221_X1 g0785(.A(new_n324), .B1(new_n722), .B2(new_n749), .C1(new_n244), .C2(new_n719), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT114), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n979), .B1(new_n985), .B2(new_n987), .ZN(new_n988));
  AOI211_X1 g0788(.A(G116), .B(new_n520), .C1(G68), .C2(G77), .ZN(new_n989));
  OAI21_X1  g0789(.A(KEYINPUT50), .B1(new_n313), .B2(G50), .ZN(new_n990));
  OR3_X1    g0790(.A1(new_n313), .A2(KEYINPUT50), .A3(G50), .ZN(new_n991));
  NAND4_X1  g0791(.A1(new_n989), .A2(new_n990), .A3(new_n991), .A4(new_n264), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n966), .B1(new_n233), .B2(G45), .ZN(new_n993));
  NOR3_X1   g0793(.A1(new_n661), .A2(new_n324), .A3(new_n658), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n992), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(G107), .B2(new_n224), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n988), .A2(new_n715), .B1(new_n716), .B2(new_n996), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n997), .B(new_n704), .C1(new_n643), .C2(new_n767), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(new_n926), .B2(new_n702), .ZN(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n971), .A2(new_n1000), .ZN(G393));
  OAI221_X1 g0801(.A(new_n716), .B1(new_n455), .B2(new_n224), .C1(new_n245), .C2(new_n966), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n746), .A2(new_n286), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(G50), .A2(new_n727), .B1(new_n723), .B2(G143), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(new_n313), .B2(new_n753), .ZN(new_n1005));
  AOI211_X1 g0805(.A(new_n1003), .B(new_n1005), .C1(G68), .C2(new_n743), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n734), .A2(G159), .B1(new_n755), .B2(G150), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n1007), .B(KEYINPUT51), .Z(new_n1008));
  NAND4_X1  g0808(.A1(new_n1006), .A2(new_n250), .A3(new_n793), .A4(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n250), .B1(new_n723), .B2(G322), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n1010), .B1(new_n352), .B2(new_n719), .C1(new_n742), .C2(new_n794), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n1011), .B(KEYINPUT115), .Z(new_n1012));
  AOI22_X1  g0812(.A1(new_n734), .A2(G311), .B1(new_n755), .B2(G317), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n1013), .B(KEYINPUT52), .Z(new_n1014));
  AOI22_X1  g0814(.A1(new_n789), .A2(G116), .B1(new_n727), .B2(G303), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1012), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n753), .A2(new_n747), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1009), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n779), .B1(new_n1018), .B2(new_n715), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n1002), .B(new_n1019), .C1(new_n896), .C2(new_n767), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n940), .A2(new_n941), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1020), .B1(new_n1021), .B2(new_n702), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n660), .B1(new_n970), .B2(new_n1021), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1022), .B1(new_n1023), .B2(new_n942), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n1024), .ZN(G390));
  AND2_X1   g0825(.A1(new_n773), .A2(G330), .ZN(new_n1026));
  AND2_X1   g0826(.A1(new_n814), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1027), .A2(KEYINPUT117), .A3(new_n873), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n864), .B1(new_n870), .B2(new_n873), .ZN(new_n1029));
  NOR3_X1   g0829(.A1(new_n1029), .A2(new_n865), .A3(new_n867), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n673), .A2(new_n635), .A3(new_n815), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1031), .A2(new_n816), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT116), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n873), .A2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n824), .B1(new_n820), .B2(new_n822), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(KEYINPUT116), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1032), .A2(new_n1034), .A3(new_n1036), .ZN(new_n1037));
  AND2_X1   g0837(.A1(new_n840), .A2(new_n841), .ZN(new_n1038));
  AND3_X1   g0838(.A1(new_n1037), .A2(new_n1038), .A3(new_n863), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1028), .B1(new_n1030), .B2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n867), .B1(new_n842), .B2(new_n866), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n870), .A2(new_n873), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(new_n863), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1037), .A2(new_n1038), .A3(new_n863), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n696), .A2(new_n1026), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n1046), .A2(new_n1035), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT117), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1027), .A2(new_n1048), .ZN(new_n1049));
  NAND4_X1  g0849(.A1(new_n1044), .A2(new_n1045), .A3(new_n1047), .A4(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1040), .A2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n433), .A2(G330), .A3(new_n814), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n881), .A2(new_n626), .A3(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n873), .B1(new_n696), .B2(new_n1026), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT118), .ZN(new_n1055));
  AND2_X1   g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n814), .A2(new_n873), .A3(new_n1026), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n870), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1032), .ZN(new_n1060));
  AND2_X1   g0860(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n1060), .B1(new_n1035), .B2(new_n1046), .C1(new_n1061), .C2(new_n1027), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1053), .B1(new_n1059), .B2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n660), .B1(new_n1051), .B2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(new_n1051), .B2(new_n1063), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1051), .A2(new_n703), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1041), .A2(new_n712), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n324), .B1(new_n722), .B2(new_n747), .C1(new_n202), .C2(new_n719), .ZN(new_n1068));
  AOI211_X1 g0868(.A(new_n1003), .B(new_n1068), .C1(G97), .C2(new_n797), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n743), .A2(G87), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n734), .A2(G116), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(G283), .A2(new_n755), .B1(new_n727), .B2(G107), .ZN(new_n1072));
  NAND4_X1  g0872(.A1(new_n1069), .A2(new_n1070), .A3(new_n1071), .A4(new_n1072), .ZN(new_n1073));
  OR3_X1    g0873(.A1(new_n742), .A2(KEYINPUT53), .A3(new_n314), .ZN(new_n1074));
  OAI21_X1  g0874(.A(KEYINPUT53), .B1(new_n742), .B2(new_n314), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(KEYINPUT54), .B(G143), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n753), .A2(new_n1076), .B1(new_n719), .B2(new_n289), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(G125), .B2(new_n723), .ZN(new_n1078));
  INV_X1    g0878(.A(G137), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n250), .B1(new_n726), .B2(new_n1079), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n746), .A2(new_n377), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n1080), .B(new_n1081), .C1(G132), .C2(new_n734), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n1074), .A2(new_n1075), .A3(new_n1078), .A4(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(G128), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n748), .A2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1073), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n1086), .A2(new_n715), .B1(new_n313), .B2(new_n803), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1067), .A2(new_n704), .A3(new_n1087), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1065), .A2(new_n1066), .A3(new_n1088), .ZN(G378));
  AND2_X1   g0889(.A1(new_n876), .A2(new_n878), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT56), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT55), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n632), .B1(new_n319), .B2(new_n320), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  OR2_X1    g0894(.A1(new_n349), .A2(new_n1094), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n338), .B(new_n1093), .C1(new_n345), .C2(new_n348), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1092), .B1(new_n1095), .B2(new_n1097), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n349), .A2(new_n1094), .ZN(new_n1099));
  NOR3_X1   g0899(.A1(new_n1099), .A2(new_n1096), .A3(KEYINPUT55), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1091), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1095), .A2(new_n1097), .A3(new_n1092), .ZN(new_n1102));
  OAI21_X1  g0902(.A(KEYINPUT55), .B1(new_n1099), .B2(new_n1096), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1102), .A2(new_n1103), .A3(KEYINPUT56), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1101), .A2(KEYINPUT120), .A3(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(new_n858), .B2(G330), .ZN(new_n1106));
  NAND4_X1  g0906(.A1(new_n1038), .A2(KEYINPUT40), .A3(new_n814), .A4(new_n826), .ZN(new_n1107));
  AND3_X1   g0907(.A1(new_n853), .A2(KEYINPUT108), .A3(new_n843), .ZN(new_n1108));
  AOI21_X1  g0908(.A(KEYINPUT108), .B1(new_n853), .B2(new_n843), .ZN(new_n1109));
  OAI211_X1 g0909(.A(G330), .B(new_n1107), .C1(new_n1108), .C2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT119), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n1111), .A2(KEYINPUT120), .ZN(new_n1112));
  AOI21_X1  g0912(.A(KEYINPUT119), .B1(new_n1101), .B2(new_n1104), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1101), .A2(KEYINPUT119), .A3(new_n1104), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1112), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n1110), .A2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1090), .B1(new_n1106), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n856), .A2(new_n857), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1104), .ZN(new_n1120));
  AOI21_X1  g0920(.A(KEYINPUT56), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1121));
  NOR3_X1   g0921(.A1(new_n1120), .A2(new_n1121), .A3(new_n1111), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n1122), .A2(new_n1113), .B1(new_n1111), .B2(KEYINPUT120), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n1119), .A2(new_n1123), .A3(G330), .A4(new_n1107), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1105), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1110), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1124), .A2(new_n1126), .A3(new_n879), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1118), .A2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1053), .B1(new_n1051), .B2(new_n1063), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(KEYINPUT57), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT57), .ZN(new_n1132));
  AOI211_X1 g0932(.A(new_n1132), .B(new_n1129), .C1(new_n1118), .C2(new_n1127), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT121), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n702), .B1(new_n1118), .B2(new_n1127), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n713), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n742), .A2(new_n1076), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(G132), .A2(new_n727), .B1(new_n797), .B2(G137), .ZN(new_n1139));
  OAI221_X1 g0939(.A(new_n1139), .B1(new_n314), .B2(new_n746), .C1(new_n1084), .C2(new_n735), .ZN(new_n1140));
  AOI211_X1 g0940(.A(new_n1138), .B(new_n1140), .C1(G125), .C2(new_n755), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(new_n1141), .B(KEYINPUT59), .ZN(new_n1142));
  AOI21_X1  g0942(.A(G41), .B1(new_n723), .B2(G124), .ZN(new_n1143));
  AOI21_X1  g0943(.A(G33), .B1(new_n720), .B2(G159), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1142), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n289), .B1(new_n254), .B2(G41), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n734), .A2(G107), .B1(G283), .B2(new_n723), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1147), .B1(new_n244), .B2(new_n748), .ZN(new_n1148));
  NOR4_X1   g0948(.A1(new_n1148), .A2(G41), .A3(new_n250), .A4(new_n945), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n720), .A2(G58), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n455), .A2(new_n726), .B1(new_n753), .B2(new_n360), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(new_n743), .B2(G77), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1149), .A2(new_n1150), .A3(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1153), .B(KEYINPUT58), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1145), .A2(new_n1146), .A3(new_n1154), .ZN(new_n1155));
  AOI211_X1 g0955(.A(new_n779), .B(new_n1137), .C1(new_n715), .C2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n803), .A2(new_n289), .ZN(new_n1157));
  AND2_X1   g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1135), .B1(new_n1136), .B2(new_n1158), .ZN(new_n1159));
  AND3_X1   g0959(.A1(new_n1124), .A2(new_n1126), .A3(new_n879), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n879), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n703), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1162), .A2(KEYINPUT121), .A3(new_n1163), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n1134), .A2(new_n659), .B1(new_n1159), .B2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(G375));
  NAND2_X1  g0966(.A1(new_n755), .A2(G132), .ZN(new_n1167));
  OAI221_X1 g0967(.A(new_n1167), .B1(new_n726), .B2(new_n1076), .C1(new_n735), .C2(new_n1079), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n324), .B1(new_n1168), .B2(KEYINPUT122), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n1169), .B(new_n1150), .C1(KEYINPUT122), .C2(new_n1168), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n742), .A2(new_n377), .B1(new_n1084), .B2(new_n722), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(new_n1171), .B(KEYINPUT124), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n746), .A2(new_n289), .B1(new_n753), .B2(new_n314), .ZN(new_n1173));
  XOR2_X1   g0973(.A(new_n1173), .B(KEYINPUT123), .Z(new_n1174));
  NOR3_X1   g0974(.A1(new_n1170), .A2(new_n1172), .A3(new_n1174), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(G107), .A2(new_n797), .B1(new_n727), .B2(G116), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1176), .B1(new_n742), .B2(new_n455), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n250), .B(new_n950), .C1(G294), .C2(new_n755), .ZN(new_n1178));
  OAI221_X1 g0978(.A(new_n1178), .B1(new_n563), .B2(new_n722), .C1(new_n360), .C2(new_n746), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n1177), .B(new_n1179), .C1(G283), .C2(new_n734), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n715), .B1(new_n1175), .B2(new_n1180), .ZN(new_n1181));
  OAI221_X1 g0981(.A(new_n1181), .B1(G68), .B2(new_n804), .C1(new_n1061), .C2(new_n713), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1182), .A2(new_n779), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1059), .A2(new_n1062), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1183), .B1(new_n1184), .B2(new_n703), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1059), .A2(new_n1062), .A3(new_n1053), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1186), .A2(new_n919), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1185), .B1(new_n1187), .B2(new_n1063), .ZN(G381));
  OR2_X1    g0988(.A1(G393), .A2(G396), .ZN(new_n1189));
  NOR3_X1   g0989(.A1(G387), .A2(new_n1189), .A3(G390), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  AND3_X1   g0991(.A1(new_n1065), .A2(new_n1066), .A3(new_n1088), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1165), .A2(new_n1192), .ZN(new_n1193));
  OR4_X1    g0993(.A1(G384), .A2(new_n1191), .A3(G381), .A4(new_n1193), .ZN(G407));
  OAI211_X1 g0994(.A(G407), .B(G213), .C1(G343), .C2(new_n1193), .ZN(G409));
  INV_X1    g0995(.A(KEYINPUT62), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1159), .A2(new_n1164), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1130), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1198), .A2(new_n1132), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1128), .A2(KEYINPUT57), .A3(new_n1130), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1199), .A2(new_n1200), .A3(new_n659), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1192), .B1(new_n1197), .B2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT60), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n660), .B1(new_n1186), .B2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1063), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n1204), .B(new_n1205), .C1(new_n1203), .C2(new_n1186), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1206), .A2(G384), .A3(new_n1185), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(G384), .B1(new_n1206), .B2(new_n1185), .ZN(new_n1209));
  OR2_X1    g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1136), .A2(new_n1158), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1129), .B1(new_n1118), .B2(new_n1127), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(new_n919), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1211), .A2(new_n1192), .A3(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n633), .A2(G213), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  NOR3_X1   g1016(.A1(new_n1202), .A2(new_n1210), .A3(new_n1216), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1196), .B1(new_n1217), .B2(KEYINPUT126), .ZN(new_n1218));
  AOI21_X1  g1018(.A(G378), .B1(new_n919), .B2(new_n1212), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n1219), .A2(new_n1211), .B1(G213), .B2(new_n633), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1220), .B1(new_n1165), .B2(new_n1192), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n633), .A2(G213), .A3(G2897), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(new_n1210), .B(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(KEYINPUT61), .B1(new_n1221), .B2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1210), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1225), .B(new_n1220), .C1(new_n1165), .C2(new_n1192), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT126), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1226), .A2(new_n1227), .A3(KEYINPUT62), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1218), .A2(new_n1224), .A3(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT127), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(G390), .A2(new_n944), .A3(new_n968), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1232), .A2(KEYINPUT125), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(G387), .A2(new_n1024), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(new_n1232), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(G393), .A2(G396), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1189), .A2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1233), .B1(new_n1235), .B2(new_n1238), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1234), .A2(new_n1232), .A3(KEYINPUT125), .A4(new_n1237), .ZN(new_n1240));
  AND2_X1   g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1218), .A2(new_n1224), .A3(new_n1228), .A4(KEYINPUT127), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1231), .A2(new_n1241), .A3(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(KEYINPUT61), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1217), .A2(KEYINPUT63), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT63), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1246), .B1(new_n1221), .B2(new_n1223), .ZN(new_n1247));
  OAI211_X1 g1047(.A(new_n1244), .B(new_n1245), .C1(new_n1217), .C2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1243), .A2(new_n1248), .ZN(G405));
  INV_X1    g1049(.A(new_n1202), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1193), .A2(new_n1250), .ZN(new_n1251));
  XNOR2_X1  g1051(.A(new_n1251), .B(new_n1210), .ZN(new_n1252));
  XNOR2_X1  g1052(.A(new_n1241), .B(new_n1252), .ZN(G402));
endmodule


