//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 1 1 1 0 0 0 1 1 0 0 0 1 0 1 0 1 1 0 0 0 0 1 1 0 1 1 1 0 0 0 0 1 1 1 1 0 0 1 1 1 1 1 0 1 0 1 0 1 0 0 0 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:28:08 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n890, new_n891,
    new_n892, new_n893, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966;
  INV_X1    g000(.A(KEYINPUT30), .ZN(new_n187));
  XNOR2_X1  g001(.A(G143), .B(G146), .ZN(new_n188));
  XNOR2_X1  g002(.A(KEYINPUT0), .B(G128), .ZN(new_n189));
  OR2_X1    g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n188), .A2(KEYINPUT0), .A3(G128), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  NAND2_X1  g006(.A1(KEYINPUT65), .A2(G131), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT11), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT64), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n196), .A2(G134), .ZN(new_n197));
  INV_X1    g011(.A(G134), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n198), .A2(KEYINPUT64), .ZN(new_n199));
  OAI21_X1  g013(.A(G137), .B1(new_n197), .B2(new_n199), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n198), .A2(G137), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n195), .B1(new_n200), .B2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n198), .A2(KEYINPUT64), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n196), .A2(G134), .ZN(new_n205));
  INV_X1    g019(.A(G137), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n204), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(new_n195), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n194), .B1(new_n203), .B2(new_n209), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n206), .B1(new_n204), .B2(new_n205), .ZN(new_n211));
  OAI21_X1  g025(.A(KEYINPUT11), .B1(new_n211), .B2(new_n201), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n212), .A2(new_n193), .A3(new_n208), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n192), .B1(new_n210), .B2(new_n213), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n207), .B1(G134), .B2(new_n206), .ZN(new_n215));
  INV_X1    g029(.A(G146), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G143), .ZN(new_n217));
  INV_X1    g031(.A(G143), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G146), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT1), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n221), .B1(G143), .B2(new_n216), .ZN(new_n222));
  INV_X1    g036(.A(G128), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n220), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n217), .A2(new_n219), .A3(new_n221), .A4(G128), .ZN(new_n225));
  AOI22_X1  g039(.A1(new_n215), .A2(G131), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G131), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n212), .A2(new_n227), .A3(new_n208), .ZN(new_n228));
  AND2_X1   g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n187), .B1(new_n214), .B2(new_n229), .ZN(new_n230));
  XNOR2_X1  g044(.A(G116), .B(G119), .ZN(new_n231));
  XNOR2_X1  g045(.A(KEYINPUT2), .B(G113), .ZN(new_n232));
  XNOR2_X1  g046(.A(new_n231), .B(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n192), .ZN(new_n235));
  AND3_X1   g049(.A1(new_n212), .A2(new_n193), .A3(new_n208), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n193), .B1(new_n212), .B2(new_n208), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n235), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n226), .A2(new_n228), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n238), .A2(KEYINPUT30), .A3(new_n239), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n230), .A2(new_n234), .A3(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G237), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(KEYINPUT66), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT66), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G237), .ZN(new_n245));
  AOI21_X1  g059(.A(G953), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G210), .ZN(new_n247));
  XOR2_X1   g061(.A(KEYINPUT26), .B(G101), .Z(new_n248));
  XNOR2_X1  g062(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g063(.A(KEYINPUT67), .B(KEYINPUT27), .ZN(new_n250));
  XNOR2_X1  g064(.A(new_n249), .B(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n238), .A2(new_n233), .A3(new_n239), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n241), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(KEYINPUT31), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT31), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n241), .A2(new_n255), .A3(new_n251), .A4(new_n252), .ZN(new_n256));
  INV_X1    g070(.A(new_n251), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT28), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n252), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n234), .B1(new_n214), .B2(new_n229), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n258), .B1(new_n261), .B2(new_n252), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n257), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n254), .A2(new_n256), .A3(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(G472), .ZN(new_n265));
  INV_X1    g079(.A(G902), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n264), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(KEYINPUT32), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT32), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n267), .A2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT68), .ZN(new_n272));
  NOR3_X1   g086(.A1(new_n260), .A2(new_n262), .A3(new_n257), .ZN(new_n273));
  AOI21_X1  g087(.A(G902), .B1(new_n273), .B2(KEYINPUT29), .ZN(new_n274));
  INV_X1    g088(.A(new_n262), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n275), .A2(new_n251), .A3(new_n259), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT29), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n241), .A2(new_n252), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(new_n257), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n276), .A2(new_n277), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n274), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n272), .B1(new_n281), .B2(G472), .ZN(new_n282));
  AOI211_X1 g096(.A(KEYINPUT68), .B(new_n265), .C1(new_n274), .C2(new_n280), .ZN(new_n283));
  OAI211_X1 g097(.A(new_n269), .B(new_n271), .C1(new_n282), .C2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G217), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n285), .B1(G234), .B2(new_n266), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT16), .ZN(new_n287));
  NAND2_X1  g101(.A1(KEYINPUT70), .A2(G125), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(G140), .ZN(new_n289));
  INV_X1    g103(.A(G140), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n290), .A2(KEYINPUT70), .A3(G125), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n287), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(KEYINPUT16), .B1(new_n290), .B2(G125), .ZN(new_n293));
  OR3_X1    g107(.A1(new_n292), .A2(G146), .A3(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(G146), .B1(new_n292), .B2(new_n293), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(G119), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(G128), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n223), .A2(G119), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  XNOR2_X1  g114(.A(KEYINPUT24), .B(G110), .ZN(new_n301));
  OR2_X1    g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  OR2_X1    g116(.A1(new_n302), .A2(KEYINPUT69), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT23), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n304), .B1(G119), .B2(new_n223), .ZN(new_n305));
  NOR3_X1   g119(.A1(new_n297), .A2(KEYINPUT23), .A3(G128), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n298), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(G110), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n302), .A2(KEYINPUT69), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n296), .A2(new_n303), .A3(new_n308), .A4(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(G110), .ZN(new_n311));
  OAI211_X1 g125(.A(new_n311), .B(new_n298), .C1(new_n305), .C2(new_n306), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n300), .A2(new_n301), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n290), .A2(G125), .ZN(new_n314));
  INV_X1    g128(.A(G125), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G140), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n314), .A2(new_n316), .A3(new_n216), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(KEYINPUT71), .ZN(new_n318));
  XNOR2_X1  g132(.A(G125), .B(G140), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT71), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n319), .A2(new_n320), .A3(new_n216), .ZN(new_n321));
  AOI22_X1  g135(.A1(new_n312), .A2(new_n313), .B1(new_n318), .B2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT72), .ZN(new_n323));
  AND3_X1   g137(.A1(new_n322), .A2(new_n323), .A3(new_n295), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n323), .B1(new_n322), .B2(new_n295), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n310), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT73), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  OAI211_X1 g142(.A(new_n310), .B(KEYINPUT73), .C1(new_n324), .C2(new_n325), .ZN(new_n329));
  XNOR2_X1  g143(.A(KEYINPUT22), .B(G137), .ZN(new_n330));
  INV_X1    g144(.A(G953), .ZN(new_n331));
  AND3_X1   g145(.A1(new_n331), .A2(G221), .A3(G234), .ZN(new_n332));
  XOR2_X1   g146(.A(new_n330), .B(new_n332), .Z(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n328), .A2(new_n329), .A3(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n326), .A2(new_n327), .A3(new_n333), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(KEYINPUT25), .B1(new_n337), .B2(new_n266), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT25), .ZN(new_n339));
  AOI211_X1 g153(.A(new_n339), .B(G902), .C1(new_n335), .C2(new_n336), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n286), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n286), .A2(G902), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n342), .B(KEYINPUT74), .ZN(new_n343));
  INV_X1    g157(.A(new_n337), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n341), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  AND2_X1   g160(.A1(new_n284), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT81), .ZN(new_n348));
  OR2_X1    g162(.A1(KEYINPUT75), .A2(KEYINPUT3), .ZN(new_n349));
  NAND2_X1  g163(.A1(KEYINPUT75), .A2(KEYINPUT3), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(G107), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(G104), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(G101), .ZN(new_n356));
  INV_X1    g170(.A(G104), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(G107), .ZN(new_n358));
  OAI22_X1  g172(.A1(new_n357), .A2(G107), .B1(KEYINPUT75), .B2(KEYINPUT3), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n355), .A2(new_n356), .A3(new_n358), .A4(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n231), .A2(KEYINPUT5), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n297), .A2(G116), .ZN(new_n362));
  OR2_X1    g176(.A1(new_n362), .A2(KEYINPUT5), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n361), .A2(G113), .A3(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(G116), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(G119), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n362), .A2(new_n366), .ZN(new_n367));
  OR2_X1    g181(.A1(new_n367), .A2(new_n232), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n356), .B1(new_n353), .B2(new_n358), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n360), .A2(new_n364), .A3(new_n368), .A4(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n353), .B1(new_n349), .B2(new_n350), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n359), .A2(new_n358), .ZN(new_n374));
  OAI21_X1  g188(.A(G101), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n360), .A2(new_n375), .A3(KEYINPUT4), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT4), .ZN(new_n377));
  OAI211_X1 g191(.A(new_n377), .B(G101), .C1(new_n373), .C2(new_n374), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n376), .A2(new_n234), .A3(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n372), .B1(new_n379), .B2(KEYINPUT79), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT79), .ZN(new_n381));
  NAND4_X1  g195(.A1(new_n376), .A2(new_n381), .A3(new_n234), .A4(new_n378), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  XNOR2_X1  g197(.A(G110), .B(G122), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n380), .A2(new_n384), .A3(new_n382), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n386), .A2(KEYINPUT6), .A3(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT6), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n383), .A2(new_n389), .A3(new_n385), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n192), .A2(G125), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n224), .A2(new_n315), .A3(new_n225), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(G224), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n394), .A2(G953), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n393), .B(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n388), .A2(new_n390), .A3(new_n396), .ZN(new_n397));
  XOR2_X1   g211(.A(new_n384), .B(KEYINPUT8), .Z(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  AOI22_X1  g213(.A1(new_n360), .A2(new_n370), .B1(new_n364), .B2(new_n368), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n399), .B1(new_n372), .B2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n392), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n315), .B1(new_n190), .B2(new_n191), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT7), .ZN(new_n404));
  OAI22_X1  g218(.A1(new_n402), .A2(new_n403), .B1(new_n404), .B2(new_n395), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n395), .A2(new_n404), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n391), .A2(new_n392), .A3(new_n406), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n401), .A2(KEYINPUT80), .A3(new_n405), .A4(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT80), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n405), .A2(new_n407), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n360), .A2(new_n370), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n364), .A2(new_n368), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n398), .B1(new_n413), .B2(new_n371), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n409), .B1(new_n410), .B2(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n387), .A2(new_n408), .A3(new_n415), .ZN(new_n416));
  AND2_X1   g230(.A1(new_n416), .A2(new_n266), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n397), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g232(.A(G210), .B1(G237), .B2(G902), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n348), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  AOI211_X1 g235(.A(KEYINPUT81), .B(new_n419), .C1(new_n397), .C2(new_n417), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n397), .A2(new_n417), .A3(new_n419), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(KEYINPUT82), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT82), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n397), .A2(new_n417), .A3(new_n426), .A4(new_n419), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n423), .A2(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(G214), .B1(G237), .B2(G902), .ZN(new_n430));
  XOR2_X1   g244(.A(new_n430), .B(KEYINPUT78), .Z(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(G475), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n244), .A2(G237), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n242), .A2(KEYINPUT66), .ZN(new_n436));
  OAI211_X1 g250(.A(G214), .B(new_n331), .C1(new_n435), .C2(new_n436), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n437), .A2(new_n218), .ZN(new_n438));
  AOI21_X1  g252(.A(G143), .B1(new_n246), .B2(G214), .ZN(new_n439));
  OAI21_X1  g253(.A(G131), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT17), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n437), .A2(new_n218), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n246), .A2(G143), .A3(G214), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n442), .A2(new_n227), .A3(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n440), .A2(new_n441), .A3(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT87), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n296), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n294), .A2(KEYINPUT87), .A3(new_n295), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n227), .B1(new_n442), .B2(new_n443), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(KEYINPUT17), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n445), .A2(new_n447), .A3(new_n448), .A4(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n318), .A2(new_n321), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n289), .A2(new_n291), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n452), .B1(new_n216), .B2(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n442), .A2(KEYINPUT83), .A3(new_n443), .ZN(new_n456));
  NAND2_X1  g270(.A1(KEYINPUT18), .A2(G131), .ZN(new_n457));
  AND2_X1   g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n456), .A2(new_n457), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n455), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n451), .A2(new_n460), .ZN(new_n461));
  XNOR2_X1  g275(.A(G113), .B(G122), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n462), .B(new_n357), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n451), .A2(new_n460), .A3(new_n463), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n434), .B1(new_n467), .B2(new_n266), .ZN(new_n468));
  NOR2_X1   g282(.A1(G475), .A2(G902), .ZN(new_n469));
  AND3_X1   g283(.A1(new_n442), .A2(new_n227), .A3(new_n443), .ZN(new_n470));
  OAI21_X1  g284(.A(KEYINPUT84), .B1(new_n470), .B2(new_n449), .ZN(new_n471));
  INV_X1    g285(.A(new_n295), .ZN(new_n472));
  AOI21_X1  g286(.A(KEYINPUT85), .B1(new_n453), .B2(KEYINPUT19), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n453), .A2(KEYINPUT19), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT19), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n319), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n473), .B1(new_n477), .B2(KEYINPUT85), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n472), .B1(new_n478), .B2(new_n216), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT84), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n440), .A2(new_n480), .A3(new_n444), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n471), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n463), .B1(new_n482), .B2(new_n460), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n466), .B1(new_n483), .B2(KEYINPUT86), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT86), .ZN(new_n485));
  AOI211_X1 g299(.A(new_n485), .B(new_n463), .C1(new_n482), .C2(new_n460), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n469), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(KEYINPUT20), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT20), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n489), .B(new_n469), .C1(new_n484), .C2(new_n486), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n468), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  XNOR2_X1  g305(.A(KEYINPUT21), .B(G898), .ZN(new_n492));
  NAND2_X1  g306(.A1(G234), .A2(G237), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n492), .A2(G902), .A3(G953), .A4(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n493), .A2(G952), .A3(new_n331), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  XOR2_X1   g310(.A(new_n496), .B(KEYINPUT90), .Z(new_n497));
  INV_X1    g311(.A(G122), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(G116), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n365), .A2(G122), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n499), .B1(new_n500), .B2(KEYINPUT14), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(KEYINPUT14), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n501), .B1(KEYINPUT88), .B2(new_n502), .ZN(new_n503));
  OR2_X1    g317(.A1(new_n502), .A2(KEYINPUT88), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n352), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  AND2_X1   g319(.A1(new_n499), .A2(new_n500), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(new_n352), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n204), .A2(new_n205), .ZN(new_n508));
  XNOR2_X1  g322(.A(G128), .B(G143), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n508), .A2(new_n509), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n507), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  OR2_X1    g327(.A1(new_n505), .A2(new_n513), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n506), .B(new_n352), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n218), .A2(G128), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT13), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n518), .B1(G128), .B2(new_n218), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n516), .A2(new_n517), .ZN(new_n520));
  OAI21_X1  g334(.A(G134), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n515), .A2(new_n521), .A3(new_n510), .ZN(new_n522));
  XOR2_X1   g336(.A(KEYINPUT9), .B(G234), .Z(new_n523));
  NAND3_X1  g337(.A1(new_n523), .A2(G217), .A3(new_n331), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  AND3_X1   g339(.A1(new_n514), .A2(new_n522), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n525), .B1(new_n514), .B2(new_n522), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n266), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n528), .A2(KEYINPUT89), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT15), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(G478), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  AOI22_X1  g346(.A1(new_n528), .A2(KEYINPUT89), .B1(new_n530), .B2(G478), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n532), .B1(new_n533), .B2(new_n529), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n491), .A2(new_n497), .A3(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT91), .ZN(new_n537));
  XNOR2_X1  g351(.A(new_n536), .B(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(G469), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n539), .A2(new_n266), .ZN(new_n540));
  XOR2_X1   g354(.A(KEYINPUT77), .B(KEYINPUT10), .Z(new_n541));
  NAND2_X1  g355(.A1(new_n224), .A2(new_n225), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NOR3_X1   g357(.A1(new_n411), .A2(new_n543), .A3(KEYINPUT76), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT76), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n373), .A2(new_n374), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n369), .B1(new_n546), .B2(new_n356), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n545), .B1(new_n547), .B2(new_n542), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n541), .B1(new_n544), .B2(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n376), .A2(new_n235), .A3(new_n378), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n547), .A2(KEYINPUT10), .A3(new_n542), .ZN(new_n551));
  AND2_X1   g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n236), .A2(new_n237), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n549), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n553), .ZN(new_n555));
  INV_X1    g369(.A(new_n541), .ZN(new_n556));
  OAI21_X1  g370(.A(KEYINPUT76), .B1(new_n411), .B2(new_n543), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n547), .A2(new_n545), .A3(new_n542), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n550), .A2(new_n551), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n555), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n554), .A2(new_n561), .ZN(new_n562));
  XNOR2_X1  g376(.A(G110), .B(G140), .ZN(new_n563));
  INV_X1    g377(.A(G227), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n564), .A2(G953), .ZN(new_n565));
  XOR2_X1   g379(.A(new_n563), .B(new_n565), .Z(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n562), .A2(new_n567), .ZN(new_n568));
  AOI22_X1  g382(.A1(new_n557), .A2(new_n558), .B1(new_n543), .B2(new_n411), .ZN(new_n569));
  OAI21_X1  g383(.A(KEYINPUT12), .B1(new_n569), .B2(new_n553), .ZN(new_n570));
  OAI22_X1  g384(.A1(new_n544), .A2(new_n548), .B1(new_n542), .B2(new_n547), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT12), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n571), .A2(new_n572), .A3(new_n555), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n570), .A2(new_n573), .A3(new_n554), .A4(new_n566), .ZN(new_n574));
  AOI21_X1  g388(.A(G902), .B1(new_n568), .B2(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n540), .B1(new_n575), .B2(new_n539), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n554), .A2(new_n561), .A3(new_n566), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n570), .A2(new_n573), .A3(new_n554), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n578), .B1(new_n567), .B2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n576), .B1(new_n539), .B2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(G221), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n583), .B1(new_n523), .B2(new_n266), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n347), .A2(new_n433), .A3(new_n538), .A4(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(KEYINPUT92), .B(G101), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n588), .B(new_n589), .ZN(G3));
  INV_X1    g404(.A(KEYINPUT33), .ZN(new_n591));
  OR3_X1    g405(.A1(new_n526), .A2(new_n527), .A3(new_n591), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n591), .B1(new_n526), .B2(new_n527), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n592), .A2(G478), .A3(new_n266), .A4(new_n593), .ZN(new_n594));
  NOR2_X1   g408(.A1(KEYINPUT93), .A2(G478), .ZN(new_n595));
  AND2_X1   g409(.A1(KEYINPUT93), .A2(G478), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n528), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n488), .A2(new_n490), .ZN(new_n600));
  INV_X1    g414(.A(new_n468), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n599), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT94), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n430), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n419), .B1(new_n397), .B2(new_n417), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n605), .B1(new_n607), .B2(new_n424), .ZN(new_n608));
  OAI21_X1  g422(.A(KEYINPUT94), .B1(new_n491), .B2(new_n599), .ZN(new_n609));
  AND4_X1   g423(.A1(new_n497), .A2(new_n604), .A3(new_n608), .A4(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n264), .A2(new_n266), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(G472), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n267), .ZN(new_n613));
  NOR3_X1   g427(.A1(new_n586), .A2(new_n345), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n610), .A2(new_n614), .ZN(new_n615));
  XOR2_X1   g429(.A(KEYINPUT34), .B(G104), .Z(new_n616));
  XNOR2_X1  g430(.A(new_n615), .B(new_n616), .ZN(G6));
  INV_X1    g431(.A(KEYINPUT95), .ZN(new_n618));
  AND3_X1   g432(.A1(new_n488), .A2(new_n618), .A3(new_n490), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n618), .B1(new_n488), .B2(new_n490), .ZN(new_n620));
  OAI211_X1 g434(.A(new_n601), .B(new_n534), .C1(new_n619), .C2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n424), .ZN(new_n622));
  OAI211_X1 g436(.A(new_n430), .B(new_n497), .C1(new_n622), .C2(new_n606), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n614), .A2(new_n624), .ZN(new_n625));
  XOR2_X1   g439(.A(KEYINPUT35), .B(G107), .Z(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G9));
  NAND3_X1  g441(.A1(new_n538), .A2(new_n433), .A3(new_n587), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT97), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n334), .A2(KEYINPUT36), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n326), .B(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n343), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  AND3_X1   g447(.A1(new_n341), .A2(KEYINPUT96), .A3(new_n633), .ZN(new_n634));
  AOI21_X1  g448(.A(KEYINPUT96), .B1(new_n341), .B2(new_n633), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n629), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n341), .A2(new_n633), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT96), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n341), .A2(KEYINPUT96), .A3(new_n633), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n639), .A2(KEYINPUT97), .A3(new_n640), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n636), .A2(new_n641), .A3(new_n267), .A4(new_n612), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n628), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(KEYINPUT37), .B(G110), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G12));
  INV_X1    g459(.A(KEYINPUT98), .ZN(new_n646));
  INV_X1    g460(.A(G900), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n493), .A2(new_n647), .A3(G902), .A4(G953), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n495), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n646), .B1(new_n621), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n600), .A2(KEYINPUT95), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n488), .A2(new_n618), .A3(new_n490), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n468), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n654), .A2(KEYINPUT98), .A3(new_n534), .A4(new_n649), .ZN(new_n655));
  AND3_X1   g469(.A1(new_n651), .A2(new_n655), .A3(new_n608), .ZN(new_n656));
  AND4_X1   g470(.A1(new_n284), .A2(new_n636), .A3(new_n641), .A4(new_n587), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(G128), .ZN(G30));
  XOR2_X1   g473(.A(new_n649), .B(KEYINPUT39), .Z(new_n660));
  NOR2_X1   g474(.A1(new_n586), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(KEYINPUT40), .ZN(new_n662));
  XNOR2_X1  g476(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n429), .B(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n253), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n251), .B1(new_n261), .B2(new_n252), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n266), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(G472), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n269), .A2(new_n271), .A3(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n634), .A2(new_n635), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n491), .A2(new_n535), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NOR3_X1   g486(.A1(new_n670), .A2(new_n672), .A3(new_n605), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n662), .A2(new_n664), .A3(new_n669), .A4(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G143), .ZN(G45));
  NAND3_X1  g489(.A1(new_n608), .A2(new_n602), .A3(new_n649), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(KEYINPUT100), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n657), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G146), .ZN(G48));
  NAND2_X1  g493(.A1(new_n568), .A2(new_n574), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n680), .A2(new_n539), .A3(new_n266), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n575), .A2(new_n539), .ZN(new_n683));
  NOR3_X1   g497(.A1(new_n682), .A2(new_n683), .A3(new_n584), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n610), .A2(new_n347), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(KEYINPUT41), .B(G113), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(G15));
  NAND3_X1  g501(.A1(new_n347), .A2(new_n624), .A3(new_n684), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G116), .ZN(G18));
  AND3_X1   g503(.A1(new_n636), .A2(new_n641), .A3(new_n284), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n684), .A2(new_n608), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n690), .A2(new_n538), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(KEYINPUT101), .B(G119), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n693), .B(new_n694), .ZN(G21));
  AOI21_X1  g509(.A(KEYINPUT102), .B1(new_n264), .B2(new_n266), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n613), .A2(new_n697), .ZN(new_n698));
  AOI211_X1 g512(.A(KEYINPUT102), .B(G472), .C1(new_n264), .C2(new_n266), .ZN(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n698), .A2(new_n346), .A3(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT103), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n696), .B1(new_n612), .B2(new_n267), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n704), .A2(new_n699), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n705), .A2(KEYINPUT103), .A3(new_n346), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(new_n684), .ZN(new_n708));
  NOR3_X1   g522(.A1(new_n672), .A2(new_n708), .A3(new_n623), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(KEYINPUT104), .B(G122), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(G24));
  INV_X1    g526(.A(KEYINPUT106), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT105), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n714), .B1(new_n602), .B2(new_n649), .ZN(new_n715));
  NOR4_X1   g529(.A1(new_n491), .A2(new_n599), .A3(KEYINPUT105), .A4(new_n650), .ZN(new_n716));
  OAI211_X1 g530(.A(new_n705), .B(new_n670), .C1(new_n715), .C2(new_n716), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n713), .B1(new_n717), .B2(new_n691), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n602), .A2(new_n649), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(KEYINPUT105), .ZN(new_n720));
  INV_X1    g534(.A(new_n716), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NOR4_X1   g536(.A1(new_n704), .A2(new_n634), .A3(new_n635), .A4(new_n699), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n722), .A2(new_n723), .A3(KEYINPUT106), .A4(new_n692), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n718), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G125), .ZN(G27));
  INV_X1    g540(.A(KEYINPUT107), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n579), .A2(new_n567), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n727), .B1(new_n728), .B2(new_n577), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n577), .A2(new_n727), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  NOR3_X1   g545(.A1(new_n729), .A2(new_n539), .A3(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n540), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n681), .A2(new_n733), .ZN(new_n734));
  OAI21_X1  g548(.A(KEYINPUT108), .B1(new_n732), .B2(new_n734), .ZN(new_n735));
  OAI211_X1 g549(.A(G469), .B(new_n730), .C1(new_n580), .C2(new_n727), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT108), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n736), .A2(new_n737), .A3(new_n576), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n584), .B1(new_n735), .B2(new_n738), .ZN(new_n739));
  NOR3_X1   g553(.A1(new_n423), .A2(new_n605), .A3(new_n428), .ZN(new_n740));
  AND2_X1   g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n741), .A2(new_n347), .A3(KEYINPUT42), .A4(new_n722), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT42), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n739), .A2(new_n740), .A3(new_n284), .A4(new_n346), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n715), .A2(new_n716), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n743), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n742), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G131), .ZN(G33));
  NAND4_X1  g562(.A1(new_n741), .A2(new_n347), .A3(new_n651), .A4(new_n655), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G134), .ZN(G36));
  INV_X1    g564(.A(KEYINPUT45), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n539), .B1(new_n581), .B2(new_n751), .ZN(new_n752));
  OAI211_X1 g566(.A(KEYINPUT45), .B(new_n730), .C1(new_n580), .C2(new_n727), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n540), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  OR2_X1    g568(.A1(new_n754), .A2(KEYINPUT46), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n682), .B1(new_n754), .B2(KEYINPUT46), .ZN(new_n756));
  AOI211_X1 g570(.A(new_n584), .B(new_n660), .C1(new_n755), .C2(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n670), .A2(new_n613), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(KEYINPUT109), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT109), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n670), .A2(new_n760), .A3(new_n613), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n491), .A2(new_n598), .ZN(new_n762));
  XOR2_X1   g576(.A(new_n762), .B(KEYINPUT43), .Z(new_n763));
  NAND3_X1  g577(.A1(new_n759), .A2(new_n761), .A3(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT44), .ZN(new_n765));
  OAI211_X1 g579(.A(new_n757), .B(new_n740), .C1(new_n764), .C2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(new_n764), .ZN(new_n767));
  OAI21_X1  g581(.A(KEYINPUT110), .B1(new_n767), .B2(KEYINPUT44), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT110), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n764), .A2(new_n769), .A3(new_n765), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n766), .B1(new_n768), .B2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(new_n206), .ZN(G39));
  NAND2_X1  g586(.A1(new_n755), .A2(new_n756), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n585), .ZN(new_n774));
  OR2_X1    g588(.A1(new_n774), .A2(KEYINPUT47), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(KEYINPUT47), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n429), .A2(new_n430), .ZN(new_n777));
  NOR4_X1   g591(.A1(new_n777), .A2(new_n284), .A3(new_n346), .A4(new_n719), .ZN(new_n778));
  AND3_X1   g592(.A1(new_n775), .A2(new_n776), .A3(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(new_n290), .ZN(G42));
  NOR2_X1   g594(.A1(new_n682), .A2(new_n683), .ZN(new_n781));
  INV_X1    g595(.A(new_n781), .ZN(new_n782));
  OR2_X1    g596(.A1(new_n782), .A2(KEYINPUT49), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(KEYINPUT49), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n783), .A2(new_n431), .A3(new_n585), .A4(new_n784), .ZN(new_n785));
  NOR3_X1   g599(.A1(new_n664), .A2(new_n785), .A3(new_n762), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n669), .A2(new_n345), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n657), .B1(new_n656), .B2(new_n677), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n649), .B(KEYINPUT113), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n341), .A2(new_n633), .A3(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(KEYINPUT114), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n671), .A2(new_n608), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n792), .A2(new_n669), .A3(new_n739), .A4(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n789), .A2(new_n725), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(KEYINPUT52), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT52), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n789), .A2(new_n725), .A3(new_n797), .A4(new_n794), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n742), .A2(new_n746), .ZN(new_n799));
  OAI211_X1 g613(.A(new_n347), .B(new_n684), .C1(new_n610), .C2(new_n624), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n710), .A2(new_n800), .A3(new_n693), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT112), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n534), .A2(KEYINPUT111), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT111), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n532), .B(new_n805), .C1(new_n533), .C2(new_n529), .ZN(new_n806));
  AND3_X1   g620(.A1(new_n804), .A2(new_n649), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n654), .A2(new_n807), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n803), .B1(new_n777), .B2(new_n808), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n740), .A2(KEYINPUT112), .A3(new_n654), .A4(new_n807), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n657), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n741), .A2(new_n723), .A3(new_n722), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n811), .A2(new_n749), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n804), .A2(new_n806), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(new_n491), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n815), .B1(new_n491), .B2(new_n599), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n433), .A2(new_n614), .A3(new_n497), .A4(new_n816), .ZN(new_n817));
  OAI211_X1 g631(.A(new_n588), .B(new_n817), .C1(new_n628), .C2(new_n642), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n813), .A2(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n796), .A2(new_n798), .A3(new_n802), .A4(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT53), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n820), .B(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(KEYINPUT54), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT115), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n796), .A2(new_n824), .A3(new_n802), .A4(new_n798), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n820), .A2(new_n825), .A3(KEYINPUT53), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n820), .B1(KEYINPUT53), .B2(new_n825), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n823), .B1(new_n828), .B2(KEYINPUT54), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n777), .A2(new_n495), .A3(new_n708), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n830), .A2(new_n347), .A3(new_n763), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT48), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n830), .A2(new_n787), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n604), .A2(new_n609), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n831), .A2(new_n832), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n836), .A2(G952), .A3(new_n331), .A4(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(new_n495), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n707), .A2(new_n839), .A3(new_n763), .ZN(new_n840));
  AOI211_X1 g654(.A(new_n833), .B(new_n838), .C1(new_n692), .C2(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n834), .A2(new_n491), .A3(new_n599), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n830), .A2(new_n723), .A3(new_n763), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n775), .A2(new_n776), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n845), .B1(new_n585), .B2(new_n782), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n840), .A2(new_n740), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n844), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT51), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n664), .A2(new_n430), .A3(new_n708), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n840), .A2(new_n850), .ZN(new_n851));
  NOR2_X1   g665(.A1(KEYINPUT116), .A2(KEYINPUT50), .ZN(new_n852));
  AND2_X1   g666(.A1(KEYINPUT116), .A2(KEYINPUT50), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n851), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n854), .B1(new_n851), .B2(new_n852), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n848), .A2(new_n849), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n849), .B1(new_n848), .B2(new_n855), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n841), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n829), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(G952), .A2(G953), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n860), .B(KEYINPUT117), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n788), .B1(new_n859), .B2(new_n861), .ZN(G75));
  AND3_X1   g676(.A1(new_n796), .A2(new_n798), .A3(new_n802), .ZN(new_n863));
  OAI211_X1 g677(.A(new_n863), .B(new_n819), .C1(new_n824), .C2(new_n821), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n820), .A2(new_n825), .A3(KEYINPUT53), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n864), .A2(G210), .A3(G902), .A4(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n388), .A2(new_n390), .ZN(new_n867));
  XOR2_X1   g681(.A(new_n867), .B(new_n396), .Z(new_n868));
  XNOR2_X1  g682(.A(new_n868), .B(KEYINPUT55), .ZN(new_n869));
  XOR2_X1   g683(.A(KEYINPUT119), .B(KEYINPUT56), .Z(new_n870));
  NOR2_X1   g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n866), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n331), .A2(G952), .ZN(new_n873));
  INV_X1    g687(.A(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT56), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n866), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(new_n869), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT118), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n877), .A2(KEYINPUT118), .A3(new_n869), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n875), .B1(new_n880), .B2(new_n881), .ZN(G51));
  XNOR2_X1  g696(.A(new_n540), .B(KEYINPUT57), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n864), .A2(KEYINPUT54), .A3(new_n865), .ZN(new_n884));
  AOI21_X1  g698(.A(KEYINPUT54), .B1(new_n864), .B2(new_n865), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n883), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(new_n680), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n828), .A2(G902), .A3(new_n753), .A4(new_n752), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n873), .B1(new_n887), .B2(new_n888), .ZN(G54));
  NAND4_X1  g703(.A1(new_n828), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n484), .A2(new_n486), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n890), .A2(new_n891), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n892), .A2(new_n893), .A3(new_n873), .ZN(G60));
  NAND2_X1  g708(.A1(new_n592), .A2(new_n593), .ZN(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(G478), .A2(G902), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(KEYINPUT59), .ZN(new_n898));
  OAI211_X1 g712(.A(new_n896), .B(new_n898), .C1(new_n884), .C2(new_n885), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(new_n874), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n896), .B1(new_n829), .B2(new_n898), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n900), .A2(new_n901), .ZN(G63));
  NAND2_X1  g716(.A1(G217), .A2(G902), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(KEYINPUT121), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT60), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n864), .A2(new_n865), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n873), .B1(new_n906), .B2(new_n344), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT122), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n828), .A2(new_n908), .A3(new_n631), .A4(new_n905), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n864), .A2(new_n631), .A3(new_n865), .A4(new_n905), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(KEYINPUT122), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n907), .A2(new_n909), .A3(new_n911), .ZN(new_n912));
  XNOR2_X1  g726(.A(KEYINPUT120), .B(KEYINPUT61), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n907), .A2(KEYINPUT61), .A3(new_n910), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(G66));
  OAI21_X1  g730(.A(G953), .B1(new_n492), .B2(new_n394), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n801), .A2(new_n818), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n917), .B1(new_n918), .B2(G953), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n867), .B1(G898), .B2(new_n331), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n919), .B(new_n920), .ZN(G69));
  NAND2_X1  g735(.A1(new_n230), .A2(new_n240), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n922), .B(new_n478), .Z(new_n923));
  NOR2_X1   g737(.A1(new_n331), .A2(G900), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(KEYINPUT125), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  AND3_X1   g740(.A1(new_n757), .A2(new_n347), .A3(new_n793), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n771), .A2(new_n779), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n789), .A2(new_n725), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(KEYINPUT124), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT124), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n789), .A2(new_n725), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n747), .A2(new_n749), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT126), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n928), .A2(new_n930), .A3(new_n932), .A4(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n926), .B1(new_n935), .B2(new_n331), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n930), .A2(new_n674), .A3(new_n932), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT62), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n930), .A2(KEYINPUT62), .A3(new_n674), .A4(new_n932), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  AND4_X1   g755(.A1(new_n347), .A2(new_n661), .A3(new_n740), .A4(new_n816), .ZN(new_n942));
  NOR3_X1   g756(.A1(new_n771), .A2(new_n779), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(G953), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT123), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n936), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(new_n923), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n947), .B1(new_n944), .B2(KEYINPUT123), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  OAI21_X1  g763(.A(G953), .B1(new_n564), .B2(new_n647), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(new_n950), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n946), .A2(new_n948), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n951), .A2(new_n953), .ZN(G72));
  NAND2_X1  g768(.A1(G472), .A2(G902), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n955), .B(KEYINPUT63), .Z(new_n956));
  INV_X1    g770(.A(new_n918), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n956), .B1(new_n935), .B2(new_n957), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n278), .A2(new_n251), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n873), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n941), .A2(new_n918), .A3(new_n943), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n956), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n962), .A2(new_n251), .A3(new_n278), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n253), .A2(KEYINPUT127), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(new_n279), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n822), .A2(new_n956), .A3(new_n965), .ZN(new_n966));
  AND3_X1   g780(.A1(new_n960), .A2(new_n963), .A3(new_n966), .ZN(G57));
endmodule


