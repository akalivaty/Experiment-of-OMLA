//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 1 0 0 0 0 1 0 0 1 1 0 1 0 1 1 0 1 1 1 1 0 0 1 1 0 0 1 1 1 1 0 1 0 0 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:17 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1268, new_n1269, new_n1270, new_n1271, new_n1272, new_n1273,
    new_n1274, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1333, new_n1334, new_n1335,
    new_n1336;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  OAI21_X1  g0013(.A(G50), .B1(G58), .B2(G68), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  NAND3_X1  g0017(.A1(new_n215), .A2(G20), .A3(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  AND2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OR2_X1    g0021(.A1(new_n221), .A2(KEYINPUT64), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(KEYINPUT64), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n225));
  NAND4_X1  g0025(.A1(new_n222), .A2(new_n223), .A3(new_n224), .A4(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n226), .A2(new_n210), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n213), .B(new_n218), .C1(new_n227), .C2(KEYINPUT1), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XNOR2_X1  g0037(.A(G50), .B(G68), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G58), .B(G77), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n238), .B(new_n239), .Z(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  INV_X1    g0044(.A(G169), .ZN(new_n245));
  NAND2_X1  g0045(.A1(G33), .A2(G41), .ZN(new_n246));
  INV_X1    g0046(.A(KEYINPUT65), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g0048(.A1(KEYINPUT65), .A2(G33), .A3(G41), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n248), .A2(new_n217), .A3(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G41), .ZN(new_n251));
  INV_X1    g0051(.A(G45), .ZN(new_n252));
  AOI21_X1  g0052(.A(G1), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n250), .A2(G274), .A3(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(new_n253), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n250), .A2(new_n255), .A3(G232), .ZN(new_n256));
  AND2_X1   g0056(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT76), .ZN(new_n258));
  INV_X1    g0058(.A(G33), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n258), .B1(new_n259), .B2(KEYINPUT3), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(KEYINPUT3), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT3), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n262), .A2(KEYINPUT76), .A3(G33), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n260), .A2(new_n261), .A3(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G226), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G1698), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n266), .B1(G223), .B2(G1698), .ZN(new_n267));
  INV_X1    g0067(.A(G87), .ZN(new_n268));
  OAI22_X1  g0068(.A1(new_n264), .A2(new_n267), .B1(new_n259), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n217), .A2(new_n246), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n245), .B1(new_n257), .B2(new_n272), .ZN(new_n273));
  AND2_X1   g0073(.A1(new_n257), .A2(new_n272), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n273), .B1(new_n274), .B2(G179), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT16), .ZN(new_n276));
  XNOR2_X1  g0076(.A(G58), .B(G68), .ZN(new_n277));
  NOR2_X1   g0077(.A1(G20), .A2(G33), .ZN(new_n278));
  AOI22_X1  g0078(.A1(new_n277), .A2(G20), .B1(G159), .B2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT7), .ZN(new_n280));
  XNOR2_X1  g0080(.A(KEYINPUT3), .B(G33), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n280), .B1(new_n281), .B2(G20), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n262), .A2(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n261), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n284), .A2(KEYINPUT7), .A3(new_n208), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n203), .B1(new_n282), .B2(new_n285), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n279), .B1(new_n286), .B2(KEYINPUT77), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT77), .ZN(new_n288));
  AOI211_X1 g0088(.A(new_n288), .B(new_n203), .C1(new_n282), .C2(new_n285), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n276), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(new_n216), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n264), .A2(new_n280), .A3(new_n208), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(G68), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n280), .B1(new_n264), .B2(new_n208), .ZN(new_n295));
  OAI211_X1 g0095(.A(KEYINPUT16), .B(new_n279), .C1(new_n294), .C2(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n290), .A2(new_n292), .A3(new_n296), .ZN(new_n297));
  XNOR2_X1  g0097(.A(KEYINPUT8), .B(G58), .ZN(new_n298));
  XNOR2_X1  g0098(.A(new_n298), .B(KEYINPUT68), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n208), .A2(G1), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n292), .A2(KEYINPUT67), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT67), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n291), .A2(new_n303), .A3(new_n216), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n302), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n305), .ZN(new_n308));
  AOI22_X1  g0108(.A1(new_n301), .A2(new_n307), .B1(new_n308), .B2(new_n299), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n275), .B1(new_n297), .B2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT18), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  AOI211_X1 g0112(.A(KEYINPUT18), .B(new_n275), .C1(new_n297), .C2(new_n309), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G190), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n257), .A2(new_n272), .A3(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n316), .B1(new_n274), .B2(G200), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n297), .A2(new_n309), .A3(new_n317), .ZN(new_n318));
  XNOR2_X1  g0118(.A(new_n318), .B(KEYINPUT17), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n314), .A2(new_n319), .ZN(new_n320));
  NOR3_X1   g0120(.A1(new_n306), .A2(new_n201), .A3(new_n300), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n321), .B1(new_n201), .B2(new_n308), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n302), .A2(new_n304), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n208), .A2(G33), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n299), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n204), .A2(G20), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT69), .ZN(new_n327));
  AOI22_X1  g0127(.A1(new_n326), .A2(new_n327), .B1(G150), .B2(new_n278), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n328), .B1(new_n327), .B2(new_n326), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n323), .B1(new_n325), .B2(new_n329), .ZN(new_n330));
  AND3_X1   g0130(.A1(new_n322), .A2(new_n330), .A3(KEYINPUT9), .ZN(new_n331));
  AOI21_X1  g0131(.A(KEYINPUT9), .B1(new_n322), .B2(new_n330), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT10), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n250), .A2(new_n255), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n254), .B1(new_n335), .B2(new_n265), .ZN(new_n336));
  OR2_X1    g0136(.A1(new_n336), .A2(KEYINPUT66), .ZN(new_n337));
  NOR2_X1   g0137(.A1(G222), .A2(G1698), .ZN(new_n338));
  INV_X1    g0138(.A(G1698), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n339), .A2(G223), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n281), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n341), .B(new_n271), .C1(G77), .C2(new_n281), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n336), .A2(KEYINPUT66), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n337), .A2(G190), .A3(new_n342), .A4(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n337), .A2(new_n342), .A3(new_n343), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(G200), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n333), .A2(new_n334), .A3(new_n344), .A4(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n322), .A2(new_n330), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT9), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n322), .A2(new_n330), .A3(KEYINPUT9), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n350), .A2(new_n346), .A3(new_n344), .A4(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(KEYINPUT10), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n347), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n345), .A2(new_n245), .ZN(new_n355));
  OAI211_X1 g0155(.A(new_n355), .B(new_n348), .C1(G179), .C2(new_n345), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  XNOR2_X1  g0157(.A(KEYINPUT15), .B(G87), .ZN(new_n358));
  OR3_X1    g0158(.A1(new_n358), .A2(KEYINPUT72), .A3(new_n324), .ZN(new_n359));
  OAI21_X1  g0159(.A(KEYINPUT72), .B1(new_n358), .B2(new_n324), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n208), .A2(new_n259), .ZN(new_n361));
  INV_X1    g0161(.A(G77), .ZN(new_n362));
  OAI22_X1  g0162(.A1(new_n298), .A2(new_n361), .B1(new_n208), .B2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT71), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n359), .B(new_n360), .C1(new_n363), .C2(new_n364), .ZN(new_n365));
  AND2_X1   g0165(.A1(new_n363), .A2(new_n364), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n292), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n308), .A2(new_n292), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n300), .A2(new_n362), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n368), .A2(new_n369), .B1(new_n362), .B2(new_n308), .ZN(new_n370));
  AND2_X1   g0170(.A1(new_n367), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(G244), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n254), .B1(new_n335), .B2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT70), .ZN(new_n374));
  OR2_X1    g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n281), .A2(G238), .A3(G1698), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n281), .A2(G232), .A3(new_n339), .ZN(new_n377));
  INV_X1    g0177(.A(G107), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n376), .B(new_n377), .C1(new_n378), .C2(new_n281), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(new_n271), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n373), .A2(new_n374), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n375), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n371), .B1(new_n245), .B2(new_n382), .ZN(new_n383));
  OR2_X1    g0183(.A1(new_n382), .A2(G179), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n382), .A2(G200), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n386), .B(new_n371), .C1(new_n315), .C2(new_n382), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  NOR3_X1   g0188(.A1(new_n320), .A2(new_n357), .A3(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n250), .A2(new_n255), .A3(G238), .ZN(new_n390));
  NAND2_X1  g0190(.A1(G33), .A2(G97), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  NOR2_X1   g0192(.A1(G226), .A2(G1698), .ZN(new_n393));
  INV_X1    g0193(.A(G232), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n393), .B1(new_n394), .B2(G1698), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n392), .B1(new_n395), .B2(new_n281), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n254), .B(new_n390), .C1(new_n396), .C2(new_n270), .ZN(new_n397));
  OAI21_X1  g0197(.A(KEYINPUT73), .B1(new_n397), .B2(KEYINPUT13), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n394), .A2(G1698), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n399), .B1(G226), .B2(G1698), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n391), .B1(new_n400), .B2(new_n284), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n216), .B1(new_n247), .B2(new_n246), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n253), .B1(new_n402), .B2(new_n249), .ZN(new_n403));
  AOI22_X1  g0203(.A1(new_n401), .A2(new_n271), .B1(new_n403), .B2(G238), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT73), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT13), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n404), .A2(new_n405), .A3(new_n406), .A4(new_n254), .ZN(new_n407));
  AND2_X1   g0207(.A1(new_n398), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n397), .A2(KEYINPUT13), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT74), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n397), .A2(KEYINPUT74), .A3(KEYINPUT13), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(G200), .B1(new_n408), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n308), .A2(new_n203), .ZN(new_n415));
  XNOR2_X1  g0215(.A(new_n415), .B(KEYINPUT12), .ZN(new_n416));
  AOI22_X1  g0216(.A1(new_n278), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n417), .B1(new_n362), .B2(new_n324), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n323), .A2(new_n418), .A3(KEYINPUT11), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n368), .B(G68), .C1(G1), .C2(new_n208), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n416), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(KEYINPUT11), .B1(new_n323), .B2(new_n418), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n404), .A2(new_n406), .A3(new_n254), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n424), .A2(G190), .A3(new_n409), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n414), .A2(new_n423), .A3(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  AND3_X1   g0227(.A1(new_n397), .A2(KEYINPUT74), .A3(KEYINPUT13), .ZN(new_n428));
  AOI21_X1  g0228(.A(KEYINPUT74), .B1(new_n397), .B2(KEYINPUT13), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n398), .A2(new_n407), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n245), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT14), .ZN(new_n433));
  OAI21_X1  g0233(.A(KEYINPUT75), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  AND3_X1   g0234(.A1(new_n424), .A2(G179), .A3(new_n409), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n435), .B1(new_n432), .B2(new_n433), .ZN(new_n436));
  OAI21_X1  g0236(.A(G169), .B1(new_n408), .B2(new_n413), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT75), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n437), .A2(new_n438), .A3(KEYINPUT14), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n434), .A2(new_n436), .A3(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n423), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n427), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  AND2_X1   g0242(.A1(new_n389), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n308), .A2(new_n378), .ZN(new_n445));
  XNOR2_X1  g0245(.A(new_n445), .B(KEYINPUT25), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n207), .A2(G33), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n302), .A2(new_n304), .A3(new_n305), .A4(new_n447), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n448), .A2(new_n378), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT83), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT24), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT22), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n208), .A2(G87), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n454), .B1(new_n284), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(G33), .A2(G116), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n457), .A2(G20), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT23), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n459), .B1(new_n208), .B2(G107), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n378), .A2(KEYINPUT23), .A3(G20), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n458), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n456), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(KEYINPUT22), .A2(G87), .ZN(new_n464));
  NOR3_X1   g0264(.A1(new_n264), .A2(G20), .A3(new_n464), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n452), .B(new_n453), .C1(new_n463), .C2(new_n465), .ZN(new_n466));
  AND2_X1   g0266(.A1(new_n466), .A2(new_n292), .ZN(new_n467));
  AND3_X1   g0267(.A1(new_n260), .A2(new_n261), .A3(new_n263), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n468), .A2(KEYINPUT22), .A3(new_n208), .A4(G87), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n469), .A2(KEYINPUT83), .A3(new_n456), .A4(new_n462), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n452), .B1(new_n463), .B2(new_n465), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n470), .A2(new_n471), .A3(KEYINPUT24), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n451), .B1(new_n467), .B2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(G250), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(new_n339), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n475), .B1(G257), .B2(new_n339), .ZN(new_n476));
  INV_X1    g0276(.A(G294), .ZN(new_n477));
  OAI22_X1  g0277(.A1(new_n264), .A2(new_n476), .B1(new_n259), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(new_n271), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n252), .A2(G1), .ZN(new_n480));
  AND2_X1   g0280(.A1(KEYINPUT5), .A2(G41), .ZN(new_n481));
  NOR2_X1   g0281(.A1(KEYINPUT5), .A2(G41), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  AND2_X1   g0283(.A1(new_n250), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(G264), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n207), .A2(G45), .ZN(new_n486));
  OR2_X1    g0286(.A1(KEYINPUT5), .A2(G41), .ZN(new_n487));
  NAND2_X1  g0287(.A1(KEYINPUT5), .A2(G41), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n489), .A2(new_n250), .A3(G274), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n479), .A2(new_n485), .A3(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT84), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n491), .A2(new_n492), .A3(G169), .ZN(new_n493));
  AOI22_X1  g0293(.A1(new_n271), .A2(new_n478), .B1(new_n484), .B2(G264), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n494), .A2(G179), .A3(new_n490), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n492), .B1(new_n491), .B2(G169), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n473), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(G200), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n491), .A2(new_n501), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n502), .B1(G190), .B2(new_n491), .ZN(new_n503));
  AND2_X1   g0303(.A1(new_n473), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n500), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n250), .A2(new_n483), .A3(G270), .ZN(new_n506));
  AND2_X1   g0306(.A1(new_n490), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n284), .A2(G303), .ZN(new_n508));
  INV_X1    g0308(.A(G264), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(G1698), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n510), .B1(G257), .B2(G1698), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n508), .B1(new_n264), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n271), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n507), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(G200), .ZN(new_n515));
  AND2_X1   g0315(.A1(new_n291), .A2(new_n216), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n516), .A2(G116), .A3(new_n305), .A4(new_n447), .ZN(new_n517));
  INV_X1    g0317(.A(G116), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n207), .A2(new_n518), .A3(G13), .A4(G20), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT82), .ZN(new_n520));
  AND2_X1   g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n519), .A2(new_n520), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n517), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n291), .A2(new_n216), .B1(G20), .B2(new_n518), .ZN(new_n524));
  NAND2_X1  g0324(.A1(G33), .A2(G283), .ZN(new_n525));
  INV_X1    g0325(.A(G97), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n525), .B(new_n208), .C1(G33), .C2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT20), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n524), .A2(KEYINPUT20), .A3(new_n527), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n523), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n515), .B(new_n532), .C1(new_n315), .C2(new_n514), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT21), .ZN(new_n534));
  NOR2_X1   g0334(.A1(G257), .A2(G1698), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n535), .B1(new_n509), .B2(G1698), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n536), .A2(new_n261), .A3(new_n260), .A4(new_n263), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n270), .B1(new_n537), .B2(new_n508), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n490), .A2(new_n506), .ZN(new_n539));
  OAI21_X1  g0339(.A(G169), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n534), .B1(new_n540), .B2(new_n532), .ZN(new_n541));
  INV_X1    g0341(.A(G179), .ZN(new_n542));
  NOR3_X1   g0342(.A1(new_n538), .A2(new_n539), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n530), .A2(new_n531), .ZN(new_n544));
  OR2_X1    g0344(.A1(new_n521), .A2(new_n522), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n544), .A2(new_n545), .A3(new_n517), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n514), .A2(new_n546), .A3(KEYINPUT21), .A4(G169), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n533), .A2(new_n541), .A3(new_n547), .A4(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n372), .A2(G1698), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n550), .B1(G238), .B2(G1698), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n457), .B1(new_n264), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(KEYINPUT81), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT81), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n554), .B(new_n457), .C1(new_n264), .C2(new_n551), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n553), .A2(new_n271), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n486), .A2(new_n474), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n250), .B(new_n557), .C1(G274), .C2(new_n486), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n556), .A2(G190), .A3(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n468), .A2(new_n208), .A3(G68), .ZN(new_n560));
  NOR2_X1   g0360(.A1(G97), .A2(G107), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n561), .A2(new_n268), .B1(new_n391), .B2(new_n208), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT19), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(G97), .ZN(new_n564));
  OAI22_X1  g0364(.A1(new_n562), .A2(new_n563), .B1(new_n324), .B2(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n516), .B1(new_n560), .B2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(new_n358), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n567), .A2(new_n305), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n448), .A2(new_n268), .ZN(new_n569));
  NOR3_X1   g0369(.A1(new_n566), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n559), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n501), .B1(new_n556), .B2(new_n558), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n448), .A2(new_n358), .ZN(new_n574));
  NOR3_X1   g0374(.A1(new_n566), .A2(new_n568), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n555), .A2(new_n271), .ZN(new_n576));
  NOR2_X1   g0376(.A1(G238), .A2(G1698), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n577), .B1(new_n372), .B2(G1698), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n578), .A2(new_n261), .A3(new_n260), .A4(new_n263), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n554), .B1(new_n579), .B2(new_n457), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n558), .B1(new_n576), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(G169), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n556), .A2(G179), .A3(new_n558), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n575), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NOR3_X1   g0384(.A1(new_n549), .A2(new_n573), .A3(new_n584), .ZN(new_n585));
  MUX2_X1   g0385(.A(new_n305), .B(new_n448), .S(G97), .Z(new_n586));
  INV_X1    g0386(.A(KEYINPUT79), .ZN(new_n587));
  AOI21_X1  g0387(.A(KEYINPUT7), .B1(new_n284), .B2(new_n208), .ZN(new_n588));
  AOI211_X1 g0388(.A(new_n280), .B(G20), .C1(new_n261), .C2(new_n283), .ZN(new_n589));
  OAI21_X1  g0389(.A(G107), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT6), .ZN(new_n591));
  AND2_X1   g0391(.A1(G97), .A2(G107), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n591), .B1(new_n592), .B2(new_n561), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n378), .A2(KEYINPUT6), .A3(G97), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n208), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  OAI21_X1  g0395(.A(KEYINPUT78), .B1(new_n361), .B2(new_n362), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT78), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n278), .A2(new_n597), .A3(G77), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n590), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n587), .B1(new_n601), .B2(new_n292), .ZN(new_n602));
  AOI211_X1 g0402(.A(KEYINPUT79), .B(new_n516), .C1(new_n590), .C2(new_n600), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n586), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n372), .A2(G1698), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n260), .A2(new_n263), .A3(new_n605), .A4(new_n261), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT4), .ZN(new_n607));
  AND2_X1   g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n261), .A2(new_n283), .A3(G250), .A4(G1698), .ZN(new_n609));
  AND2_X1   g0409(.A1(KEYINPUT4), .A2(G244), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n261), .A2(new_n283), .A3(new_n610), .A4(new_n339), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n609), .A2(new_n611), .A3(new_n525), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n271), .B1(new_n608), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n250), .A2(new_n483), .A3(G257), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n490), .A2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(G169), .B1(new_n613), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n606), .A2(new_n607), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n618), .A2(new_n609), .A3(new_n611), .A4(new_n525), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n615), .B1(new_n619), .B2(new_n271), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n617), .B1(new_n542), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n604), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n613), .A2(new_n616), .A3(new_n315), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n623), .B1(new_n620), .B2(G200), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n624), .B(new_n586), .C1(new_n603), .C2(new_n602), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n622), .A2(new_n625), .A3(KEYINPUT80), .ZN(new_n626));
  AOI21_X1  g0426(.A(KEYINPUT80), .B1(new_n622), .B2(new_n625), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n505), .B(new_n585), .C1(new_n626), .C2(new_n627), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n444), .A2(new_n628), .ZN(G372));
  INV_X1    g0429(.A(new_n319), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n440), .A2(new_n441), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n426), .A2(new_n384), .A3(new_n383), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n630), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n297), .A2(new_n309), .ZN(new_n634));
  INV_X1    g0434(.A(new_n275), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(KEYINPUT18), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n310), .A2(new_n311), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n637), .A2(KEYINPUT88), .A3(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT88), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n640), .B1(new_n312), .B2(new_n313), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n354), .B1(new_n633), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n356), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT26), .ZN(new_n646));
  NOR4_X1   g0446(.A1(new_n622), .A2(new_n573), .A3(new_n646), .A4(new_n584), .ZN(new_n647));
  INV_X1    g0447(.A(new_n575), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT85), .ZN(new_n649));
  AND3_X1   g0449(.A1(new_n582), .A2(new_n649), .A3(new_n583), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n649), .B1(new_n582), .B2(new_n583), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n648), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n622), .ZN(new_n653));
  OR2_X1    g0453(.A1(new_n572), .A2(KEYINPUT86), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n572), .A2(KEYINPUT86), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n654), .A2(new_n559), .A3(new_n570), .A4(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n652), .A2(new_n653), .A3(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n647), .B1(new_n657), .B2(new_n646), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT87), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n652), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n582), .A2(new_n583), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(KEYINPUT85), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n582), .A2(new_n649), .A3(new_n583), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n575), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(KEYINPUT87), .ZN(new_n665));
  AND3_X1   g0465(.A1(new_n541), .A2(new_n547), .A3(new_n548), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n496), .A2(new_n498), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n666), .B1(new_n667), .B2(new_n473), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n668), .A2(new_n652), .A3(new_n656), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n473), .A2(new_n503), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n670), .A2(new_n622), .A3(new_n625), .ZN(new_n671));
  OAI211_X1 g0471(.A(new_n660), .B(new_n665), .C1(new_n669), .C2(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n443), .B1(new_n658), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n645), .A2(new_n673), .ZN(G369));
  NAND3_X1  g0474(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n675));
  OR2_X1    g0475(.A1(new_n675), .A2(KEYINPUT27), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(KEYINPUT27), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n676), .A2(G213), .A3(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(G343), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n505), .B1(new_n473), .B2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n680), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n500), .A2(new_n682), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n666), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n532), .A2(new_n680), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n687), .B1(new_n549), .B2(new_n686), .ZN(new_n688));
  XNOR2_X1  g0488(.A(KEYINPUT89), .B(G330), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n684), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n666), .A2(new_n682), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n505), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n500), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n695), .B1(new_n696), .B2(new_n682), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n693), .A2(new_n698), .ZN(G399));
  INV_X1    g0499(.A(new_n211), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(G41), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n561), .A2(new_n268), .A3(new_n518), .ZN(new_n702));
  NOR3_X1   g0502(.A1(new_n701), .A2(new_n702), .A3(new_n207), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n703), .B1(new_n215), .B2(new_n701), .ZN(new_n704));
  XOR2_X1   g0504(.A(new_n704), .B(KEYINPUT28), .Z(new_n705));
  OAI21_X1  g0505(.A(new_n680), .B1(new_n672), .B2(new_n658), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(KEYINPUT91), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT29), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT91), .ZN(new_n709));
  OAI211_X1 g0509(.A(new_n709), .B(new_n680), .C1(new_n672), .C2(new_n658), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n707), .A2(new_n708), .A3(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n664), .A2(KEYINPUT87), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n652), .A2(new_n659), .ZN(new_n713));
  OAI21_X1  g0513(.A(KEYINPUT92), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT92), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n665), .A2(new_n660), .A3(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT93), .ZN(new_n717));
  AND3_X1   g0517(.A1(new_n622), .A2(new_n625), .A3(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n717), .B1(new_n622), .B2(new_n625), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n670), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  OAI211_X1 g0520(.A(new_n714), .B(new_n716), .C1(new_n720), .C2(new_n669), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n622), .A2(new_n573), .A3(new_n584), .ZN(new_n722));
  MUX2_X1   g0522(.A(new_n722), .B(new_n657), .S(KEYINPUT26), .Z(new_n723));
  OAI211_X1 g0523(.A(KEYINPUT29), .B(new_n680), .C1(new_n721), .C2(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(KEYINPUT90), .A2(KEYINPUT30), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n543), .A2(new_n620), .A3(new_n494), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n725), .B1(new_n726), .B2(new_n581), .ZN(new_n727));
  AND3_X1   g0527(.A1(new_n494), .A2(new_n613), .A3(new_n616), .ZN(new_n728));
  INV_X1    g0528(.A(new_n581), .ZN(new_n729));
  INV_X1    g0529(.A(new_n725), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n728), .A2(new_n729), .A3(new_n543), .A4(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n620), .ZN(new_n732));
  AOI21_X1  g0532(.A(G179), .B1(new_n507), .B2(new_n513), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n732), .A2(new_n491), .A3(new_n581), .A4(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n727), .A2(new_n731), .A3(new_n734), .ZN(new_n735));
  AND3_X1   g0535(.A1(new_n735), .A2(KEYINPUT31), .A3(new_n682), .ZN(new_n736));
  AOI21_X1  g0536(.A(KEYINPUT31), .B1(new_n735), .B2(new_n682), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n738), .B1(new_n628), .B2(new_n682), .ZN(new_n739));
  AOI22_X1  g0539(.A1(new_n711), .A2(new_n724), .B1(new_n690), .B2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT94), .ZN(new_n741));
  XNOR2_X1  g0541(.A(new_n740), .B(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n705), .B1(new_n742), .B2(G1), .ZN(new_n743));
  XNOR2_X1  g0543(.A(new_n743), .B(KEYINPUT95), .ZN(G364));
  INV_X1    g0544(.A(G13), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(G20), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n207), .B1(new_n746), .B2(G45), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n701), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g0549(.A(new_n749), .B(KEYINPUT96), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n700), .A2(new_n284), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G355), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n752), .B1(G116), .B2(new_n211), .ZN(new_n753));
  OR2_X1    g0553(.A1(new_n240), .A2(new_n252), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n211), .A2(new_n264), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n755), .B1(new_n252), .B2(new_n215), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n753), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(G13), .A2(G33), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(G20), .ZN(new_n760));
  XNOR2_X1  g0560(.A(new_n760), .B(KEYINPUT97), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n216), .B1(G20), .B2(new_n245), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n750), .B1(new_n757), .B2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n208), .A2(G179), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n767), .A2(new_n315), .A3(G200), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(new_n378), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n208), .A2(new_n542), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n770), .A2(G190), .A3(new_n501), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(G190), .A2(G200), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n770), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  AOI22_X1  g0575(.A1(new_n772), .A2(G58), .B1(new_n775), .B2(G77), .ZN(new_n776));
  INV_X1    g0576(.A(KEYINPUT98), .ZN(new_n777));
  AOI211_X1 g0577(.A(new_n284), .B(new_n769), .C1(new_n776), .C2(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n767), .A2(new_n773), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(KEYINPUT32), .B1(new_n780), .B2(G159), .ZN(new_n781));
  INV_X1    g0581(.A(KEYINPUT32), .ZN(new_n782));
  INV_X1    g0582(.A(G159), .ZN(new_n783));
  NOR3_X1   g0583(.A1(new_n779), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  OAI221_X1 g0584(.A(new_n778), .B1(new_n777), .B2(new_n776), .C1(new_n781), .C2(new_n784), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n767), .A2(G190), .A3(G200), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(G87), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n770), .A2(G200), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(G190), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n788), .B1(new_n791), .B2(new_n203), .ZN(new_n792));
  NOR3_X1   g0592(.A1(new_n315), .A2(G179), .A3(G200), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(new_n208), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(new_n526), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n789), .A2(new_n315), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(new_n201), .ZN(new_n798));
  NOR4_X1   g0598(.A1(new_n785), .A2(new_n792), .A3(new_n795), .A4(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  OR2_X1    g0600(.A1(new_n800), .A2(KEYINPUT99), .ZN(new_n801));
  INV_X1    g0601(.A(G322), .ZN(new_n802));
  INV_X1    g0602(.A(G311), .ZN(new_n803));
  OAI22_X1  g0603(.A1(new_n771), .A2(new_n802), .B1(new_n774), .B2(new_n803), .ZN(new_n804));
  AOI211_X1 g0604(.A(new_n281), .B(new_n804), .C1(G329), .C2(new_n780), .ZN(new_n805));
  INV_X1    g0605(.A(G317), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(KEYINPUT33), .ZN(new_n807));
  OR2_X1    g0607(.A1(new_n806), .A2(KEYINPUT33), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n790), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n794), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n810), .A2(G294), .B1(new_n787), .B2(G303), .ZN(new_n811));
  INV_X1    g0611(.A(new_n768), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n796), .A2(G326), .B1(new_n812), .B2(G283), .ZN(new_n813));
  NAND4_X1  g0613(.A1(new_n805), .A2(new_n809), .A3(new_n811), .A4(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n800), .A2(KEYINPUT99), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n801), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n766), .B1(new_n816), .B2(new_n763), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n817), .B1(new_n688), .B2(new_n761), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n749), .B1(new_n688), .B2(new_n690), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n819), .B1(new_n690), .B2(new_n688), .ZN(new_n820));
  AND2_X1   g0620(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(G396));
  OAI21_X1  g0622(.A(new_n387), .B1(new_n371), .B2(new_n680), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(new_n385), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n383), .A2(new_n384), .A3(new_n680), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n707), .A2(new_n710), .A3(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n826), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n828), .B(new_n680), .C1(new_n672), .C2(new_n658), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n739), .A2(new_n690), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n749), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n832), .B1(new_n831), .B2(new_n830), .ZN(new_n833));
  INV_X1    g0633(.A(G303), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n797), .A2(new_n834), .B1(new_n786), .B2(new_n378), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n835), .B1(G87), .B2(new_n812), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n281), .B1(new_n772), .B2(G294), .ZN(new_n837));
  AOI22_X1  g0637(.A1(G116), .A2(new_n775), .B1(new_n780), .B2(G311), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n795), .B1(G283), .B2(new_n790), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n836), .A2(new_n837), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n772), .A2(G143), .B1(new_n775), .B2(G159), .ZN(new_n841));
  INV_X1    g0641(.A(G150), .ZN(new_n842));
  INV_X1    g0642(.A(G137), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n841), .B1(new_n791), .B2(new_n842), .C1(new_n843), .C2(new_n797), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT34), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n264), .B1(new_n780), .B2(G132), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n768), .A2(new_n203), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n849), .B1(new_n202), .B2(new_n794), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n850), .B1(G50), .B2(new_n787), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n846), .A2(new_n847), .A3(new_n851), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n844), .A2(new_n845), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n840), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(new_n763), .ZN(new_n855));
  INV_X1    g0655(.A(new_n750), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n763), .A2(new_n758), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n856), .B1(new_n362), .B2(new_n857), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n855), .B(new_n858), .C1(new_n828), .C2(new_n759), .ZN(new_n859));
  AND2_X1   g0659(.A1(new_n833), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(G384));
  NOR3_X1   g0661(.A1(new_n216), .A2(new_n208), .A3(new_n518), .ZN(new_n862));
  AND2_X1   g0662(.A1(new_n593), .A2(new_n594), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n862), .B1(new_n864), .B2(KEYINPUT35), .ZN(new_n865));
  AOI22_X1  g0665(.A1(new_n865), .A2(KEYINPUT100), .B1(KEYINPUT35), .B2(new_n864), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n866), .B1(KEYINPUT100), .B2(new_n865), .ZN(new_n867));
  XNOR2_X1  g0667(.A(new_n867), .B(KEYINPUT36), .ZN(new_n868));
  OAI21_X1  g0668(.A(G77), .B1(new_n202), .B2(new_n203), .ZN(new_n869));
  OAI22_X1  g0669(.A1(new_n869), .A2(new_n214), .B1(G50), .B2(new_n203), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n870), .A2(G1), .A3(new_n745), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  XOR2_X1   g0672(.A(new_n872), .B(KEYINPUT101), .Z(new_n873));
  INV_X1    g0673(.A(KEYINPUT38), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n639), .A2(new_n641), .A3(new_n319), .ZN(new_n875));
  AOI21_X1  g0675(.A(KEYINPUT102), .B1(new_n634), .B2(new_n679), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT102), .ZN(new_n877));
  AOI211_X1 g0677(.A(new_n877), .B(new_n678), .C1(new_n297), .C2(new_n309), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  AND2_X1   g0679(.A1(new_n875), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT37), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n636), .A2(new_n881), .A3(new_n318), .ZN(new_n882));
  OAI21_X1  g0682(.A(KEYINPUT103), .B1(new_n879), .B2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n309), .ZN(new_n884));
  OAI21_X1  g0684(.A(G68), .B1(new_n588), .B2(new_n589), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n288), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n286), .A2(KEYINPUT77), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n886), .A2(new_n279), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n516), .B1(new_n888), .B2(new_n276), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n884), .B1(new_n889), .B2(new_n296), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n877), .B1(new_n890), .B2(new_n678), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n634), .A2(KEYINPUT102), .A3(new_n679), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT103), .ZN(new_n894));
  AND3_X1   g0694(.A1(new_n297), .A2(new_n309), .A3(new_n317), .ZN(new_n895));
  NOR3_X1   g0695(.A1(new_n895), .A2(new_n310), .A3(KEYINPUT37), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n893), .A2(new_n894), .A3(new_n896), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n636), .B(new_n318), .C1(new_n876), .C2(new_n878), .ZN(new_n898));
  AOI22_X1  g0698(.A1(new_n883), .A2(new_n897), .B1(new_n898), .B2(KEYINPUT37), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n874), .B1(new_n880), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n279), .B1(new_n294), .B2(new_n295), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(new_n276), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n902), .A2(new_n323), .A3(new_n296), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n309), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n635), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n679), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n905), .A2(new_n906), .A3(new_n318), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(KEYINPUT37), .ZN(new_n908));
  NOR3_X1   g0708(.A1(new_n879), .A2(KEYINPUT103), .A3(new_n882), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n894), .B1(new_n893), .B2(new_n896), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n908), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n906), .B1(new_n314), .B2(new_n319), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n911), .A2(KEYINPUT38), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n900), .A2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT39), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n631), .A2(new_n682), .ZN(new_n918));
  INV_X1    g0718(.A(new_n908), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n919), .B1(new_n883), .B2(new_n897), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n874), .B1(new_n920), .B2(new_n912), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n921), .A2(new_n914), .A3(KEYINPUT39), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n917), .A2(new_n918), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n829), .A2(new_n825), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n441), .A2(new_n682), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n631), .A2(new_n426), .A3(new_n925), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n441), .B(new_n682), .C1(new_n440), .C2(new_n427), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n924), .A2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n921), .A2(new_n914), .ZN(new_n931));
  AOI22_X1  g0731(.A1(new_n930), .A2(new_n931), .B1(new_n642), .B2(new_n678), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n923), .A2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  AND3_X1   g0734(.A1(new_n707), .A2(new_n708), .A3(new_n710), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n724), .A2(new_n443), .ZN(new_n936));
  OAI21_X1  g0736(.A(KEYINPUT104), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT104), .ZN(new_n938));
  NAND4_X1  g0738(.A1(new_n711), .A2(new_n938), .A3(new_n443), .A4(new_n724), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(new_n645), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n934), .B(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n826), .B1(new_n926), .B2(new_n927), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT105), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n739), .A2(new_n944), .ZN(new_n945));
  OAI211_X1 g0745(.A(KEYINPUT105), .B(new_n738), .C1(new_n628), .C2(new_n682), .ZN(new_n946));
  AND3_X1   g0746(.A1(new_n943), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n915), .A2(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(KEYINPUT40), .B1(new_n921), .B2(new_n914), .ZN(new_n949));
  AOI22_X1  g0749(.A1(new_n948), .A2(KEYINPUT40), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n443), .A2(new_n945), .A3(new_n946), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n950), .B(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n952), .A2(new_n689), .ZN(new_n953));
  OAI22_X1  g0753(.A1(new_n942), .A2(new_n953), .B1(new_n207), .B2(new_n746), .ZN(new_n954));
  AND2_X1   g0754(.A1(new_n942), .A2(new_n953), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n873), .B1(new_n954), .B2(new_n955), .ZN(G367));
  NOR2_X1   g0756(.A1(new_n236), .A2(new_n755), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n764), .B1(new_n211), .B2(new_n358), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n750), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n771), .A2(new_n842), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n794), .A2(new_n203), .ZN(new_n961));
  AOI211_X1 g0761(.A(new_n960), .B(new_n961), .C1(G143), .C2(new_n796), .ZN(new_n962));
  AND2_X1   g0762(.A1(new_n962), .A2(KEYINPUT111), .ZN(new_n963));
  OAI221_X1 g0763(.A(new_n281), .B1(new_n779), .B2(new_n843), .C1(new_n201), .C2(new_n774), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n812), .A2(G77), .ZN(new_n965));
  OAI221_X1 g0765(.A(new_n965), .B1(new_n202), .B2(new_n786), .C1(new_n791), .C2(new_n783), .ZN(new_n966));
  NOR3_X1   g0766(.A1(new_n963), .A2(new_n964), .A3(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(KEYINPUT111), .B2(new_n962), .ZN(new_n968));
  INV_X1    g0768(.A(G283), .ZN(new_n969));
  OAI22_X1  g0769(.A1(new_n771), .A2(new_n834), .B1(new_n774), .B2(new_n969), .ZN(new_n970));
  XOR2_X1   g0770(.A(KEYINPUT110), .B(G311), .Z(new_n971));
  OAI21_X1  g0771(.A(new_n264), .B1(new_n797), .B2(new_n971), .ZN(new_n972));
  AOI211_X1 g0772(.A(new_n970), .B(new_n972), .C1(G317), .C2(new_n780), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n787), .A2(G116), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT46), .ZN(new_n975));
  OAI22_X1  g0775(.A1(new_n794), .A2(new_n378), .B1(new_n768), .B2(new_n526), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n976), .B1(G294), .B2(new_n790), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n973), .A2(new_n975), .A3(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n968), .A2(new_n978), .ZN(new_n979));
  XOR2_X1   g0779(.A(KEYINPUT112), .B(KEYINPUT47), .Z(new_n980));
  XNOR2_X1  g0780(.A(new_n979), .B(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n959), .B1(new_n981), .B2(new_n763), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n570), .A2(new_n680), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n712), .B2(new_n713), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n652), .B(new_n656), .C1(new_n570), .C2(new_n680), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n982), .B1(new_n761), .B2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n684), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n695), .B1(new_n988), .B2(new_n694), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n989), .B(new_n691), .Z(new_n990));
  NAND2_X1  g0790(.A1(new_n742), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n604), .A2(new_n682), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n718), .B2(new_n719), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n653), .A2(new_n682), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT107), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n993), .A2(KEYINPUT107), .A3(new_n994), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n997), .A2(new_n697), .A3(new_n998), .ZN(new_n999));
  XOR2_X1   g0799(.A(KEYINPUT109), .B(KEYINPUT44), .Z(new_n1000));
  XNOR2_X1  g0800(.A(new_n999), .B(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n997), .A2(new_n998), .ZN(new_n1002));
  AND3_X1   g0802(.A1(new_n1002), .A2(KEYINPUT45), .A3(new_n698), .ZN(new_n1003));
  AOI21_X1  g0803(.A(KEYINPUT45), .B1(new_n1002), .B2(new_n698), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1001), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1005), .A2(new_n692), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n1001), .B(new_n693), .C1(new_n1003), .C2(new_n1004), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n742), .B1(new_n991), .B2(new_n1008), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n701), .B(KEYINPUT41), .Z(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n748), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT108), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1002), .A2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n997), .A2(KEYINPUT108), .A3(new_n998), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n696), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n680), .B1(new_n1016), .B2(new_n653), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n695), .B1(new_n997), .B2(new_n998), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT42), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  AND2_X1   g0820(.A1(new_n984), .A2(new_n985), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(KEYINPUT106), .B(KEYINPUT43), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(new_n1023));
  AND2_X1   g0823(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1024), .B1(KEYINPUT43), .B2(new_n986), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1020), .A2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1017), .A2(new_n1019), .A3(new_n1024), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n1030), .A2(new_n693), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1028), .B(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n987), .B1(new_n1012), .B2(new_n1033), .ZN(G387));
  NAND2_X1  g0834(.A1(new_n684), .A2(new_n762), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n298), .A2(G50), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT50), .ZN(new_n1037));
  AOI211_X1 g0837(.A(G45), .B(new_n702), .C1(G68), .C2(G77), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n755), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(new_n233), .B2(new_n252), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n751), .A2(new_n702), .B1(new_n378), .B2(new_n700), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1040), .A2(KEYINPUT113), .A3(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(new_n764), .ZN(new_n1043));
  AOI21_X1  g0843(.A(KEYINPUT113), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n750), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n772), .A2(G317), .B1(new_n775), .B2(G303), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1046), .B1(new_n791), .B2(new_n971), .C1(new_n802), .C2(new_n797), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT48), .ZN(new_n1048));
  OR2_X1    g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n794), .A2(new_n969), .B1(new_n786), .B2(new_n477), .ZN(new_n1051));
  XOR2_X1   g0851(.A(new_n1051), .B(KEYINPUT115), .Z(new_n1052));
  NAND3_X1  g0852(.A1(new_n1049), .A2(new_n1050), .A3(new_n1052), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT49), .ZN(new_n1054));
  OR2_X1    g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n768), .A2(new_n518), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n468), .B(new_n1057), .C1(G326), .C2(new_n780), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1055), .A2(new_n1056), .A3(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n264), .B1(new_n780), .B2(G150), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n1060), .B1(new_n362), .B2(new_n786), .C1(new_n526), .C2(new_n768), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT114), .Z(new_n1062));
  AOI22_X1  g0862(.A1(new_n772), .A2(G50), .B1(new_n775), .B2(G68), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n810), .A2(new_n567), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n1063), .B(new_n1064), .C1(new_n783), .C2(new_n797), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n299), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1065), .B1(new_n1066), .B2(new_n790), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1062), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1059), .A2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1045), .B1(new_n1069), .B2(new_n763), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n990), .A2(new_n748), .B1(new_n1035), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n991), .A2(new_n701), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n742), .A2(new_n990), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1071), .B1(new_n1072), .B2(new_n1073), .ZN(G393));
  INV_X1    g0874(.A(new_n1008), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1075), .A2(new_n742), .A3(new_n990), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n991), .A2(new_n1008), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1076), .A2(new_n701), .A3(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1075), .A2(new_n748), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n764), .B1(new_n526), .B2(new_n211), .C1(new_n243), .C2(new_n755), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n750), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n797), .A2(new_n806), .B1(new_n803), .B2(new_n771), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT52), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n284), .B1(new_n774), .B2(new_n477), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(G322), .B2(new_n780), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n769), .B1(G283), .B2(new_n787), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(G116), .A2(new_n810), .B1(new_n790), .B2(G303), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n1083), .A2(new_n1085), .A3(new_n1086), .A4(new_n1087), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n797), .A2(new_n842), .B1(new_n783), .B2(new_n771), .ZN(new_n1089));
  XOR2_X1   g0889(.A(new_n1089), .B(KEYINPUT51), .Z(new_n1090));
  NOR2_X1   g0890(.A1(new_n794), .A2(new_n362), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n203), .A2(new_n786), .B1(new_n768), .B2(new_n268), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n1091), .B(new_n1092), .C1(G50), .C2(new_n790), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n298), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n1094), .A2(new_n775), .B1(new_n780), .B2(G143), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1093), .A2(new_n468), .A3(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1088), .B1(new_n1090), .B2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1081), .B1(new_n1097), .B2(new_n763), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1098), .B1(new_n1029), .B2(new_n761), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1078), .A2(new_n1079), .A3(new_n1099), .ZN(G390));
  INV_X1    g0900(.A(new_n701), .ZN(new_n1101));
  NAND4_X1  g0901(.A1(new_n943), .A2(new_n945), .A3(G330), .A4(new_n946), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n918), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n917), .A2(new_n922), .B1(new_n1104), .B2(new_n929), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n928), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n680), .B(new_n824), .C1(new_n721), .C2(new_n723), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1106), .B1(new_n1107), .B2(new_n825), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n898), .A2(KEYINPUT37), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1109), .B1(new_n909), .B2(new_n910), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n875), .A2(new_n879), .ZN(new_n1111));
  AOI21_X1  g0911(.A(KEYINPUT38), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NOR3_X1   g0912(.A1(new_n920), .A2(new_n874), .A3(new_n912), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NOR3_X1   g0914(.A1(new_n1108), .A2(new_n1114), .A3(new_n918), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1103), .B1(new_n1105), .B2(new_n1115), .ZN(new_n1116));
  AND2_X1   g0916(.A1(new_n1107), .A2(new_n825), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1104), .B(new_n915), .C1(new_n1117), .C2(new_n1106), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n739), .A2(new_n690), .A3(new_n828), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT116), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1120), .A2(new_n1121), .A3(new_n928), .ZN(new_n1122));
  OAI21_X1  g0922(.A(KEYINPUT116), .B1(new_n1106), .B2(new_n1119), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n922), .ZN(new_n1125));
  AOI21_X1  g0925(.A(KEYINPUT39), .B1(new_n900), .B2(new_n914), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n930), .A2(new_n918), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n1118), .B(new_n1124), .C1(new_n1127), .C2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1116), .A2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n945), .A2(G330), .A3(new_n946), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n444), .A2(new_n1131), .ZN(new_n1132));
  AOI211_X1 g0932(.A(new_n644), .B(new_n1132), .C1(new_n937), .C2(new_n939), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1106), .B1(new_n1131), .B2(new_n826), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1124), .A2(new_n1117), .A3(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1106), .A2(new_n1119), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1102), .A2(new_n1136), .ZN(new_n1137));
  AND3_X1   g0937(.A1(new_n1137), .A2(KEYINPUT117), .A3(new_n924), .ZN(new_n1138));
  AOI21_X1  g0938(.A(KEYINPUT117), .B1(new_n1137), .B2(new_n924), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1135), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1133), .A2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1101), .B1(new_n1130), .B2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1142), .B1(new_n1130), .B2(new_n1141), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n857), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n750), .B1(new_n1066), .B2(new_n1144), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(G159), .A2(new_n810), .B1(new_n790), .B2(G137), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n796), .A2(G128), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n772), .A2(G132), .B1(new_n780), .B2(G125), .ZN(new_n1148));
  AND3_X1   g0948(.A1(new_n1146), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(KEYINPUT54), .B(G143), .ZN(new_n1150));
  XOR2_X1   g0950(.A(new_n1150), .B(KEYINPUT118), .Z(new_n1151));
  NAND2_X1  g0951(.A1(new_n787), .A2(G150), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n1151), .A2(new_n775), .B1(KEYINPUT53), .B2(new_n1152), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1149), .B(new_n1153), .C1(KEYINPUT53), .C2(new_n1152), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n281), .B1(new_n768), .B2(new_n201), .ZN(new_n1155));
  XOR2_X1   g0955(.A(new_n1155), .B(KEYINPUT119), .Z(new_n1156));
  AOI21_X1  g0956(.A(new_n1091), .B1(G283), .B2(new_n796), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1157), .B1(new_n378), .B2(new_n791), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n771), .A2(new_n518), .B1(new_n774), .B2(new_n526), .ZN(new_n1159));
  AOI211_X1 g0959(.A(new_n281), .B(new_n1159), .C1(G294), .C2(new_n780), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1160), .A2(new_n788), .A3(new_n849), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n1154), .A2(new_n1156), .B1(new_n1158), .B2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1145), .B1(new_n1162), .B2(new_n763), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1163), .B1(new_n1127), .B2(new_n759), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1164), .B1(new_n1130), .B2(new_n747), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT120), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  OAI211_X1 g0967(.A(KEYINPUT120), .B(new_n1164), .C1(new_n1130), .C2(new_n747), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1143), .A2(new_n1167), .A3(new_n1168), .ZN(G378));
  INV_X1    g0969(.A(G330), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n678), .B1(new_n322), .B2(new_n330), .ZN(new_n1171));
  AND2_X1   g0971(.A1(new_n357), .A2(new_n1171), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n357), .A2(new_n1171), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  OR3_X1    g0975(.A1(new_n1172), .A2(new_n1173), .A3(new_n1175), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1175), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n943), .A2(new_n945), .A3(new_n946), .ZN(new_n1180));
  OAI21_X1  g0980(.A(KEYINPUT40), .B1(new_n1114), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(KEYINPUT40), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n947), .A2(new_n931), .A3(new_n1182), .ZN(new_n1183));
  AOI211_X1 g0983(.A(new_n1170), .B(new_n1179), .C1(new_n1181), .C2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1180), .B1(new_n914), .B2(new_n900), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1183), .B1(new_n1185), .B2(new_n1182), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1178), .B1(new_n1186), .B2(G330), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n933), .B1(new_n1184), .B2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT122), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1179), .B1(new_n950), .B2(new_n1170), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1186), .A2(G330), .A3(new_n1178), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1190), .A2(new_n934), .A3(new_n1191), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1188), .A2(new_n1189), .A3(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1137), .A2(new_n924), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT117), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1137), .A2(KEYINPUT117), .A3(new_n924), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1107), .A2(new_n825), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n1196), .A2(new_n1197), .B1(new_n1134), .B2(new_n1199), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1133), .B1(new_n1130), .B2(new_n1200), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1190), .A2(KEYINPUT122), .A3(new_n934), .A4(new_n1191), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1193), .A2(new_n1201), .A3(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT57), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1204), .B1(new_n1188), .B2(new_n1192), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1101), .B1(new_n1206), .B2(new_n1201), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1205), .A2(new_n1207), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1193), .A2(new_n748), .A3(new_n1202), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1179), .A2(new_n758), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n749), .B1(G50), .B2(new_n1144), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n791), .A2(new_n526), .B1(new_n768), .B2(new_n202), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n961), .B(new_n1212), .C1(G116), .C2(new_n796), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n264), .A2(new_n251), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(G77), .B2(new_n787), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1215), .A2(KEYINPUT121), .ZN(new_n1216));
  OR2_X1    g1016(.A1(new_n1215), .A2(KEYINPUT121), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n771), .A2(new_n378), .B1(new_n779), .B2(new_n969), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(new_n567), .B2(new_n775), .ZN(new_n1219));
  NAND4_X1  g1019(.A1(new_n1213), .A2(new_n1216), .A3(new_n1217), .A4(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT58), .ZN(new_n1221));
  OR2_X1    g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1214), .B(new_n201), .C1(G33), .C2(G41), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1224));
  INV_X1    g1024(.A(G128), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n771), .A2(new_n1225), .B1(new_n774), .B2(new_n843), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(G132), .B2(new_n790), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(G150), .A2(new_n810), .B1(new_n796), .B2(G125), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1151), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n1227), .B(new_n1228), .C1(new_n1229), .C2(new_n786), .ZN(new_n1230));
  OR2_X1    g1030(.A1(new_n1230), .A2(KEYINPUT59), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1230), .A2(KEYINPUT59), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n812), .A2(G159), .ZN(new_n1233));
  AOI211_X1 g1033(.A(G33), .B(G41), .C1(new_n780), .C2(G124), .ZN(new_n1234));
  NAND4_X1  g1034(.A1(new_n1231), .A2(new_n1232), .A3(new_n1233), .A4(new_n1234), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1222), .A2(new_n1223), .A3(new_n1224), .A4(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1211), .B1(new_n1236), .B2(new_n763), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1210), .A2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1209), .A2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1208), .A2(new_n1240), .ZN(G375));
  INV_X1    g1041(.A(new_n1132), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n940), .A2(new_n645), .A3(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1200), .A2(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1244), .A2(new_n1141), .A3(new_n1011), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1106), .A2(new_n758), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n750), .B1(G68), .B2(new_n1144), .ZN(new_n1247));
  OAI22_X1  g1047(.A1(new_n518), .A2(new_n791), .B1(new_n797), .B2(new_n477), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1248), .B1(G97), .B2(new_n787), .ZN(new_n1249));
  OAI22_X1  g1049(.A1(new_n771), .A2(new_n969), .B1(new_n774), .B2(new_n378), .ZN(new_n1250));
  AOI211_X1 g1050(.A(new_n281), .B(new_n1250), .C1(G303), .C2(new_n780), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1249), .A2(new_n965), .A3(new_n1064), .A4(new_n1251), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(G50), .A2(new_n810), .B1(new_n796), .B2(G132), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1253), .B1(new_n783), .B2(new_n786), .ZN(new_n1254));
  OAI22_X1  g1054(.A1(new_n774), .A2(new_n842), .B1(new_n779), .B2(new_n1225), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1255), .B1(G137), .B2(new_n772), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n264), .B1(new_n812), .B2(G58), .ZN(new_n1257));
  OAI211_X1 g1057(.A(new_n1256), .B(new_n1257), .C1(new_n1229), .C2(new_n791), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1252), .B1(new_n1254), .B2(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1247), .B1(new_n1259), .B2(new_n763), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(new_n1140), .A2(new_n748), .B1(new_n1246), .B2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1245), .A2(new_n1261), .ZN(G381));
  NOR3_X1   g1062(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1263));
  XOR2_X1   g1063(.A(new_n1263), .B(KEYINPUT123), .Z(new_n1264));
  NOR4_X1   g1064(.A1(G387), .A2(G378), .A3(G390), .A4(G381), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1239), .B1(new_n1205), .B2(new_n1207), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1264), .A2(new_n1265), .A3(new_n1266), .ZN(G407));
  INV_X1    g1067(.A(G378), .ZN(new_n1268));
  INV_X1    g1068(.A(G213), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1269), .A2(G343), .ZN(new_n1270));
  AND3_X1   g1070(.A1(new_n1266), .A2(new_n1268), .A3(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT124), .ZN(new_n1272));
  AND2_X1   g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1274));
  OAI211_X1 g1074(.A(G213), .B(G407), .C1(new_n1273), .C2(new_n1274), .ZN(G409));
  NAND4_X1  g1075(.A1(new_n1193), .A2(new_n1201), .A3(new_n1202), .A4(new_n1011), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n747), .B1(new_n1188), .B2(new_n1192), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1277), .B1(new_n1210), .B2(new_n1237), .ZN(new_n1278));
  AOI21_X1  g1078(.A(G378), .B1(new_n1276), .B2(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1279), .B1(new_n1266), .B2(G378), .ZN(new_n1280));
  OAI21_X1  g1080(.A(KEYINPUT126), .B1(new_n1280), .B2(new_n1270), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1208), .A2(G378), .A3(new_n1240), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1278), .A2(new_n1276), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1268), .A2(new_n1283), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1270), .B1(new_n1282), .B2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT126), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT60), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1288), .B1(new_n1133), .B2(new_n1140), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1101), .B1(new_n1133), .B2(new_n1140), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1200), .A2(new_n1243), .A3(KEYINPUT60), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT125), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1200), .A2(new_n1243), .A3(KEYINPUT125), .A4(KEYINPUT60), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1291), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1261), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n860), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1298));
  AND2_X1   g1098(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1299));
  OAI211_X1 g1099(.A(G384), .B(new_n1261), .C1(new_n1299), .C2(new_n1291), .ZN(new_n1300));
  AND4_X1   g1100(.A1(G2897), .A2(new_n1298), .A3(new_n1270), .A4(new_n1300), .ZN(new_n1301));
  AOI22_X1  g1101(.A1(new_n1298), .A2(new_n1300), .B1(G2897), .B2(new_n1270), .ZN(new_n1302));
  OR2_X1    g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1281), .A2(new_n1287), .A3(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(G390), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(G387), .ZN(new_n1306));
  OAI211_X1 g1106(.A(G390), .B(new_n987), .C1(new_n1012), .C2(new_n1033), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  XNOR2_X1  g1108(.A(G393), .B(new_n821), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1308), .A2(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT61), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1306), .A2(new_n1307), .A3(new_n1309), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1311), .A2(new_n1312), .A3(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1298), .A2(new_n1300), .ZN(new_n1315));
  AOI211_X1 g1115(.A(new_n1270), .B(new_n1315), .C1(new_n1282), .C2(new_n1284), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1314), .B1(new_n1316), .B2(KEYINPUT63), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1315), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1285), .A2(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT63), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1304), .A2(new_n1317), .A3(new_n1321), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1312), .B1(new_n1323), .B2(new_n1285), .ZN(new_n1324));
  AND2_X1   g1124(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n1325));
  NOR2_X1   g1125(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1326), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1325), .B1(new_n1316), .B2(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1319), .A2(new_n1326), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1324), .B1(new_n1328), .B2(new_n1329), .ZN(new_n1330));
  AND2_X1   g1130(.A1(new_n1311), .A2(new_n1313), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n1322), .B1(new_n1330), .B2(new_n1331), .ZN(G405));
  NAND2_X1  g1132(.A1(G375), .A2(new_n1268), .ZN(new_n1333));
  AND3_X1   g1133(.A1(new_n1333), .A2(new_n1282), .A3(new_n1315), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1315), .B1(new_n1333), .B2(new_n1282), .ZN(new_n1335));
  NOR2_X1   g1135(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1336));
  XNOR2_X1  g1136(.A(new_n1336), .B(new_n1331), .ZN(G402));
endmodule


