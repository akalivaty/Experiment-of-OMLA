

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594;

  INV_X1 U324 ( .A(KEYINPUT26), .ZN(n464) );
  NOR2_X1 U325 ( .A1(n531), .A2(n457), .ZN(n572) );
  XOR2_X1 U326 ( .A(KEYINPUT45), .B(n390), .Z(n292) );
  XOR2_X1 U327 ( .A(KEYINPUT71), .B(G85GAT), .Z(n293) );
  XOR2_X1 U328 ( .A(KEYINPUT84), .B(G176GAT), .Z(n294) );
  XOR2_X1 U329 ( .A(n379), .B(n413), .Z(n295) );
  XNOR2_X1 U330 ( .A(G36GAT), .B(G190GAT), .ZN(n320) );
  NOR2_X1 U331 ( .A1(n543), .A2(n388), .ZN(n389) );
  XNOR2_X1 U332 ( .A(n320), .B(KEYINPUT75), .ZN(n415) );
  XNOR2_X1 U333 ( .A(n395), .B(n294), .ZN(n307) );
  NOR2_X1 U334 ( .A1(n453), .A2(n452), .ZN(n454) );
  XOR2_X1 U335 ( .A(KEYINPUT48), .B(n394), .Z(n453) );
  XNOR2_X1 U336 ( .A(n308), .B(n307), .ZN(n309) );
  NOR2_X1 U337 ( .A1(n463), .A2(n576), .ZN(n456) );
  XNOR2_X1 U338 ( .A(n464), .B(KEYINPUT92), .ZN(n465) );
  XNOR2_X1 U339 ( .A(n466), .B(n465), .ZN(n574) );
  XNOR2_X1 U340 ( .A(n383), .B(n382), .ZN(n582) );
  XNOR2_X1 U341 ( .A(n332), .B(n331), .ZN(n543) );
  INV_X1 U342 ( .A(G127GAT), .ZN(n448) );
  NOR2_X1 U343 ( .A1(n531), .A2(n447), .ZN(n544) );
  XOR2_X1 U344 ( .A(n313), .B(n312), .Z(n531) );
  XNOR2_X1 U345 ( .A(n480), .B(n479), .ZN(n510) );
  XNOR2_X1 U346 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n458) );
  XNOR2_X1 U347 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U348 ( .A(n487), .B(G50GAT), .ZN(n488) );
  XNOR2_X1 U349 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U350 ( .A(n459), .B(n458), .ZN(G1351GAT) );
  XNOR2_X1 U351 ( .A(n489), .B(n488), .ZN(G1331GAT) );
  XOR2_X1 U352 ( .A(KEYINPUT20), .B(KEYINPUT83), .Z(n297) );
  XNOR2_X1 U353 ( .A(G169GAT), .B(G190GAT), .ZN(n296) );
  XNOR2_X1 U354 ( .A(n297), .B(n296), .ZN(n313) );
  XOR2_X1 U355 ( .A(G120GAT), .B(G71GAT), .Z(n379) );
  INV_X1 U356 ( .A(KEYINPUT19), .ZN(n298) );
  NAND2_X1 U357 ( .A1(G183GAT), .A2(n298), .ZN(n301) );
  INV_X1 U358 ( .A(G183GAT), .ZN(n299) );
  NAND2_X1 U359 ( .A1(n299), .A2(KEYINPUT19), .ZN(n300) );
  NAND2_X1 U360 ( .A1(n301), .A2(n300), .ZN(n303) );
  XNOR2_X1 U361 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n302) );
  XNOR2_X1 U362 ( .A(n303), .B(n302), .ZN(n413) );
  NAND2_X1 U363 ( .A1(G227GAT), .A2(G233GAT), .ZN(n304) );
  XNOR2_X1 U364 ( .A(n295), .B(n304), .ZN(n308) );
  XOR2_X1 U365 ( .A(KEYINPUT0), .B(KEYINPUT82), .Z(n306) );
  XNOR2_X1 U366 ( .A(G113GAT), .B(G134GAT), .ZN(n305) );
  XNOR2_X1 U367 ( .A(n306), .B(n305), .ZN(n395) );
  XOR2_X1 U368 ( .A(G15GAT), .B(G127GAT), .Z(n341) );
  XOR2_X1 U369 ( .A(n309), .B(n341), .Z(n311) );
  XNOR2_X1 U370 ( .A(G43GAT), .B(G99GAT), .ZN(n310) );
  XNOR2_X1 U371 ( .A(n311), .B(n310), .ZN(n312) );
  INV_X1 U372 ( .A(KEYINPUT111), .ZN(n431) );
  XOR2_X1 U373 ( .A(KEYINPUT74), .B(G92GAT), .Z(n315) );
  XNOR2_X1 U374 ( .A(G134GAT), .B(G218GAT), .ZN(n314) );
  XNOR2_X1 U375 ( .A(n315), .B(n314), .ZN(n319) );
  XOR2_X1 U376 ( .A(KEYINPUT65), .B(KEYINPUT64), .Z(n317) );
  XNOR2_X1 U377 ( .A(KEYINPUT11), .B(KEYINPUT73), .ZN(n316) );
  XNOR2_X1 U378 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U379 ( .A(n319), .B(n318), .Z(n328) );
  XOR2_X1 U380 ( .A(G50GAT), .B(G162GAT), .Z(n444) );
  XOR2_X1 U381 ( .A(n444), .B(n415), .Z(n322) );
  NAND2_X1 U382 ( .A1(G232GAT), .A2(G233GAT), .ZN(n321) );
  XNOR2_X1 U383 ( .A(n322), .B(n321), .ZN(n326) );
  XOR2_X1 U384 ( .A(KEYINPUT7), .B(KEYINPUT8), .Z(n324) );
  XNOR2_X1 U385 ( .A(G43GAT), .B(G29GAT), .ZN(n323) );
  XNOR2_X1 U386 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U387 ( .A(KEYINPUT67), .B(n325), .Z(n368) );
  XNOR2_X1 U388 ( .A(n326), .B(n368), .ZN(n327) );
  XNOR2_X1 U389 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U390 ( .A(n329), .B(KEYINPUT10), .Z(n332) );
  XNOR2_X1 U391 ( .A(G99GAT), .B(G106GAT), .ZN(n330) );
  XNOR2_X1 U392 ( .A(n293), .B(n330), .ZN(n372) );
  XNOR2_X1 U393 ( .A(n372), .B(KEYINPUT9), .ZN(n331) );
  INV_X1 U394 ( .A(KEYINPUT110), .ZN(n387) );
  XOR2_X1 U395 ( .A(KEYINPUT15), .B(KEYINPUT77), .Z(n334) );
  XNOR2_X1 U396 ( .A(G64GAT), .B(KEYINPUT76), .ZN(n333) );
  XNOR2_X1 U397 ( .A(n334), .B(n333), .ZN(n338) );
  XOR2_X1 U398 ( .A(G78GAT), .B(G155GAT), .Z(n336) );
  XNOR2_X1 U399 ( .A(G8GAT), .B(G211GAT), .ZN(n335) );
  XNOR2_X1 U400 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U401 ( .A(n338), .B(n337), .ZN(n354) );
  XOR2_X1 U402 ( .A(KEYINPUT80), .B(KEYINPUT12), .Z(n340) );
  XNOR2_X1 U403 ( .A(KEYINPUT14), .B(KEYINPUT81), .ZN(n339) );
  XNOR2_X1 U404 ( .A(n340), .B(n339), .ZN(n345) );
  XOR2_X1 U405 ( .A(G183GAT), .B(G71GAT), .Z(n343) );
  XOR2_X1 U406 ( .A(G22GAT), .B(G1GAT), .Z(n355) );
  XNOR2_X1 U407 ( .A(n355), .B(n341), .ZN(n342) );
  XNOR2_X1 U408 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U409 ( .A(n345), .B(n344), .Z(n347) );
  NAND2_X1 U410 ( .A1(G231GAT), .A2(G233GAT), .ZN(n346) );
  XNOR2_X1 U411 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U412 ( .A(n348), .B(KEYINPUT78), .Z(n352) );
  XOR2_X1 U413 ( .A(KEYINPUT13), .B(KEYINPUT68), .Z(n350) );
  XNOR2_X1 U414 ( .A(G57GAT), .B(KEYINPUT69), .ZN(n349) );
  XNOR2_X1 U415 ( .A(n350), .B(n349), .ZN(n371) );
  XNOR2_X1 U416 ( .A(n371), .B(KEYINPUT79), .ZN(n351) );
  XNOR2_X1 U417 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U418 ( .A(n354), .B(n353), .ZN(n585) );
  XOR2_X1 U419 ( .A(n355), .B(KEYINPUT66), .Z(n357) );
  NAND2_X1 U420 ( .A1(G229GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U421 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U422 ( .A(G169GAT), .B(G8GAT), .Z(n421) );
  XOR2_X1 U423 ( .A(n358), .B(n421), .Z(n366) );
  XOR2_X1 U424 ( .A(G113GAT), .B(G15GAT), .Z(n360) );
  XNOR2_X1 U425 ( .A(G36GAT), .B(G50GAT), .ZN(n359) );
  XNOR2_X1 U426 ( .A(n360), .B(n359), .ZN(n364) );
  XOR2_X1 U427 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n362) );
  XNOR2_X1 U428 ( .A(G197GAT), .B(G141GAT), .ZN(n361) );
  XNOR2_X1 U429 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U430 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U431 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U432 ( .A(n368), .B(n367), .ZN(n577) );
  INV_X1 U433 ( .A(n577), .ZN(n550) );
  XOR2_X1 U434 ( .A(G64GAT), .B(G92GAT), .Z(n370) );
  XNOR2_X1 U435 ( .A(G176GAT), .B(G204GAT), .ZN(n369) );
  XNOR2_X1 U436 ( .A(n370), .B(n369), .ZN(n414) );
  XNOR2_X1 U437 ( .A(n414), .B(n371), .ZN(n383) );
  XOR2_X1 U438 ( .A(KEYINPUT32), .B(n372), .Z(n374) );
  NAND2_X1 U439 ( .A1(G230GAT), .A2(G233GAT), .ZN(n373) );
  XNOR2_X1 U440 ( .A(n374), .B(n373), .ZN(n378) );
  XOR2_X1 U441 ( .A(KEYINPUT72), .B(KEYINPUT33), .Z(n376) );
  XNOR2_X1 U442 ( .A(KEYINPUT31), .B(KEYINPUT70), .ZN(n375) );
  XNOR2_X1 U443 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U444 ( .A(n378), .B(n377), .ZN(n381) );
  XOR2_X1 U445 ( .A(G148GAT), .B(G78GAT), .Z(n441) );
  XOR2_X1 U446 ( .A(n379), .B(n441), .Z(n380) );
  XNOR2_X1 U447 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U448 ( .A(n582), .B(KEYINPUT41), .ZN(n555) );
  NOR2_X1 U449 ( .A1(n550), .A2(n555), .ZN(n384) );
  XNOR2_X1 U450 ( .A(n384), .B(KEYINPUT46), .ZN(n385) );
  NOR2_X1 U451 ( .A1(n585), .A2(n385), .ZN(n386) );
  XNOR2_X1 U452 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U453 ( .A(n389), .B(KEYINPUT47), .ZN(n393) );
  XOR2_X1 U454 ( .A(KEYINPUT36), .B(n543), .Z(n591) );
  INV_X1 U455 ( .A(n585), .ZN(n558) );
  NOR2_X1 U456 ( .A1(n591), .A2(n558), .ZN(n390) );
  NOR2_X1 U457 ( .A1(n582), .A2(n292), .ZN(n391) );
  NAND2_X1 U458 ( .A1(n391), .A2(n550), .ZN(n392) );
  NAND2_X1 U459 ( .A1(n393), .A2(n392), .ZN(n394) );
  XOR2_X1 U460 ( .A(n395), .B(G1GAT), .Z(n397) );
  NAND2_X1 U461 ( .A1(G225GAT), .A2(G233GAT), .ZN(n396) );
  XNOR2_X1 U462 ( .A(n397), .B(n396), .ZN(n412) );
  XOR2_X1 U463 ( .A(G85GAT), .B(G162GAT), .Z(n399) );
  XNOR2_X1 U464 ( .A(G29GAT), .B(G120GAT), .ZN(n398) );
  XNOR2_X1 U465 ( .A(n399), .B(n398), .ZN(n403) );
  XOR2_X1 U466 ( .A(KEYINPUT88), .B(KEYINPUT1), .Z(n401) );
  XNOR2_X1 U467 ( .A(KEYINPUT4), .B(G57GAT), .ZN(n400) );
  XNOR2_X1 U468 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U469 ( .A(n403), .B(n402), .Z(n410) );
  XOR2_X1 U470 ( .A(G155GAT), .B(KEYINPUT2), .Z(n405) );
  XNOR2_X1 U471 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n404) );
  XNOR2_X1 U472 ( .A(n405), .B(n404), .ZN(n443) );
  XOR2_X1 U473 ( .A(KEYINPUT6), .B(KEYINPUT5), .Z(n407) );
  XNOR2_X1 U474 ( .A(G127GAT), .B(G148GAT), .ZN(n406) );
  XNOR2_X1 U475 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U476 ( .A(n443), .B(n408), .ZN(n409) );
  XNOR2_X1 U477 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U478 ( .A(n412), .B(n411), .ZN(n525) );
  INV_X1 U479 ( .A(n525), .ZN(n506) );
  XNOR2_X1 U480 ( .A(n413), .B(n414), .ZN(n419) );
  XOR2_X1 U481 ( .A(n415), .B(KEYINPUT89), .Z(n417) );
  NAND2_X1 U482 ( .A1(G226GAT), .A2(G233GAT), .ZN(n416) );
  XNOR2_X1 U483 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U484 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U485 ( .A(n420), .B(KEYINPUT90), .Z(n423) );
  XNOR2_X1 U486 ( .A(n421), .B(KEYINPUT76), .ZN(n422) );
  XNOR2_X1 U487 ( .A(n423), .B(n422), .ZN(n429) );
  XNOR2_X1 U488 ( .A(G211GAT), .B(KEYINPUT21), .ZN(n424) );
  XNOR2_X1 U489 ( .A(n424), .B(KEYINPUT85), .ZN(n425) );
  XOR2_X1 U490 ( .A(n425), .B(KEYINPUT86), .Z(n427) );
  XNOR2_X1 U491 ( .A(G197GAT), .B(G218GAT), .ZN(n426) );
  XNOR2_X1 U492 ( .A(n427), .B(n426), .ZN(n438) );
  INV_X1 U493 ( .A(n438), .ZN(n428) );
  XOR2_X1 U494 ( .A(n429), .B(n428), .Z(n528) );
  INV_X1 U495 ( .A(n528), .ZN(n509) );
  XNOR2_X1 U496 ( .A(n509), .B(KEYINPUT27), .ZN(n467) );
  NAND2_X1 U497 ( .A1(n506), .A2(n467), .ZN(n473) );
  OR2_X1 U498 ( .A1(n453), .A2(n473), .ZN(n430) );
  XOR2_X1 U499 ( .A(n431), .B(n430), .Z(n549) );
  XOR2_X1 U500 ( .A(KEYINPUT24), .B(G204GAT), .Z(n433) );
  NAND2_X1 U501 ( .A1(G228GAT), .A2(G233GAT), .ZN(n432) );
  XNOR2_X1 U502 ( .A(n433), .B(n432), .ZN(n437) );
  XOR2_X1 U503 ( .A(KEYINPUT87), .B(KEYINPUT22), .Z(n435) );
  XNOR2_X1 U504 ( .A(G106GAT), .B(KEYINPUT23), .ZN(n434) );
  XNOR2_X1 U505 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U506 ( .A(n437), .B(n436), .Z(n440) );
  XNOR2_X1 U507 ( .A(G22GAT), .B(n438), .ZN(n439) );
  XNOR2_X1 U508 ( .A(n440), .B(n439), .ZN(n442) );
  XOR2_X1 U509 ( .A(n442), .B(n441), .Z(n446) );
  XNOR2_X1 U510 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U511 ( .A(n446), .B(n445), .ZN(n463) );
  XOR2_X1 U512 ( .A(n463), .B(KEYINPUT28), .Z(n534) );
  NAND2_X1 U513 ( .A1(n549), .A2(n534), .ZN(n447) );
  NAND2_X1 U514 ( .A1(n544), .A2(n585), .ZN(n451) );
  XOR2_X1 U515 ( .A(KEYINPUT50), .B(KEYINPUT114), .Z(n449) );
  XNOR2_X1 U516 ( .A(n451), .B(n450), .ZN(G1342GAT) );
  XOR2_X1 U517 ( .A(KEYINPUT120), .B(n509), .Z(n452) );
  XNOR2_X1 U518 ( .A(n454), .B(KEYINPUT54), .ZN(n455) );
  NAND2_X1 U519 ( .A1(n455), .A2(n525), .ZN(n576) );
  XNOR2_X1 U520 ( .A(n456), .B(KEYINPUT55), .ZN(n457) );
  NAND2_X1 U521 ( .A1(n572), .A2(n543), .ZN(n459) );
  INV_X1 U522 ( .A(KEYINPUT38), .ZN(n480) );
  INV_X1 U523 ( .A(n531), .ZN(n481) );
  NAND2_X1 U524 ( .A1(n509), .A2(n481), .ZN(n460) );
  XNOR2_X1 U525 ( .A(KEYINPUT93), .B(n460), .ZN(n461) );
  NOR2_X1 U526 ( .A1(n463), .A2(n461), .ZN(n462) );
  XNOR2_X1 U527 ( .A(n462), .B(KEYINPUT25), .ZN(n469) );
  NAND2_X1 U528 ( .A1(n463), .A2(n531), .ZN(n466) );
  NAND2_X1 U529 ( .A1(n574), .A2(n467), .ZN(n468) );
  NAND2_X1 U530 ( .A1(n469), .A2(n468), .ZN(n470) );
  XNOR2_X1 U531 ( .A(n470), .B(KEYINPUT94), .ZN(n471) );
  NAND2_X1 U532 ( .A1(n471), .A2(n525), .ZN(n476) );
  NAND2_X1 U533 ( .A1(n531), .A2(n534), .ZN(n472) );
  NOR2_X1 U534 ( .A1(n473), .A2(n472), .ZN(n474) );
  XNOR2_X1 U535 ( .A(n474), .B(KEYINPUT91), .ZN(n475) );
  NAND2_X1 U536 ( .A1(n476), .A2(n475), .ZN(n492) );
  NOR2_X1 U537 ( .A1(n591), .A2(n585), .ZN(n477) );
  NAND2_X1 U538 ( .A1(n492), .A2(n477), .ZN(n478) );
  XNOR2_X1 U539 ( .A(KEYINPUT37), .B(n478), .ZN(n524) );
  NOR2_X1 U540 ( .A1(n550), .A2(n582), .ZN(n493) );
  NAND2_X1 U541 ( .A1(n524), .A2(n493), .ZN(n479) );
  NAND2_X1 U542 ( .A1(n510), .A2(n481), .ZN(n485) );
  XOR2_X1 U543 ( .A(KEYINPUT102), .B(KEYINPUT101), .Z(n483) );
  XNOR2_X1 U544 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n482) );
  XNOR2_X1 U545 ( .A(n485), .B(n484), .ZN(G1330GAT) );
  INV_X1 U546 ( .A(n534), .ZN(n486) );
  NAND2_X1 U547 ( .A1(n510), .A2(n486), .ZN(n489) );
  XOR2_X1 U548 ( .A(KEYINPUT103), .B(KEYINPUT104), .Z(n487) );
  INV_X1 U549 ( .A(n543), .ZN(n561) );
  NAND2_X1 U550 ( .A1(n585), .A2(n561), .ZN(n490) );
  XOR2_X1 U551 ( .A(KEYINPUT16), .B(n490), .Z(n491) );
  AND2_X1 U552 ( .A1(n492), .A2(n491), .ZN(n513) );
  NAND2_X1 U553 ( .A1(n493), .A2(n513), .ZN(n502) );
  NOR2_X1 U554 ( .A1(n525), .A2(n502), .ZN(n495) );
  XNOR2_X1 U555 ( .A(KEYINPUT95), .B(KEYINPUT34), .ZN(n494) );
  XNOR2_X1 U556 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U557 ( .A(G1GAT), .B(n496), .ZN(G1324GAT) );
  NOR2_X1 U558 ( .A1(n528), .A2(n502), .ZN(n497) );
  XOR2_X1 U559 ( .A(KEYINPUT96), .B(n497), .Z(n498) );
  XNOR2_X1 U560 ( .A(G8GAT), .B(n498), .ZN(G1325GAT) );
  NOR2_X1 U561 ( .A1(n531), .A2(n502), .ZN(n500) );
  XNOR2_X1 U562 ( .A(KEYINPUT35), .B(KEYINPUT97), .ZN(n499) );
  XNOR2_X1 U563 ( .A(n500), .B(n499), .ZN(n501) );
  XOR2_X1 U564 ( .A(G15GAT), .B(n501), .Z(G1326GAT) );
  NOR2_X1 U565 ( .A1(n534), .A2(n502), .ZN(n504) );
  XNOR2_X1 U566 ( .A(KEYINPUT98), .B(KEYINPUT99), .ZN(n503) );
  XNOR2_X1 U567 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U568 ( .A(G22GAT), .B(n505), .ZN(G1327GAT) );
  XOR2_X1 U569 ( .A(G29GAT), .B(KEYINPUT39), .Z(n508) );
  NAND2_X1 U570 ( .A1(n506), .A2(n510), .ZN(n507) );
  XNOR2_X1 U571 ( .A(n508), .B(n507), .ZN(G1328GAT) );
  NAND2_X1 U572 ( .A1(n510), .A2(n509), .ZN(n511) );
  XNOR2_X1 U573 ( .A(n511), .B(KEYINPUT100), .ZN(n512) );
  XNOR2_X1 U574 ( .A(G36GAT), .B(n512), .ZN(G1329GAT) );
  NOR2_X1 U575 ( .A1(n577), .A2(n555), .ZN(n523) );
  NAND2_X1 U576 ( .A1(n523), .A2(n513), .ZN(n519) );
  NOR2_X1 U577 ( .A1(n525), .A2(n519), .ZN(n514) );
  XOR2_X1 U578 ( .A(G57GAT), .B(n514), .Z(n515) );
  XNOR2_X1 U579 ( .A(KEYINPUT42), .B(n515), .ZN(G1332GAT) );
  NOR2_X1 U580 ( .A1(n528), .A2(n519), .ZN(n517) );
  XNOR2_X1 U581 ( .A(G64GAT), .B(KEYINPUT105), .ZN(n516) );
  XNOR2_X1 U582 ( .A(n517), .B(n516), .ZN(G1333GAT) );
  NOR2_X1 U583 ( .A1(n531), .A2(n519), .ZN(n518) );
  XOR2_X1 U584 ( .A(G71GAT), .B(n518), .Z(G1334GAT) );
  NOR2_X1 U585 ( .A1(n534), .A2(n519), .ZN(n521) );
  XNOR2_X1 U586 ( .A(KEYINPUT106), .B(KEYINPUT43), .ZN(n520) );
  XNOR2_X1 U587 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U588 ( .A(G78GAT), .B(n522), .ZN(G1335GAT) );
  NAND2_X1 U589 ( .A1(n524), .A2(n523), .ZN(n533) );
  NOR2_X1 U590 ( .A1(n525), .A2(n533), .ZN(n527) );
  XNOR2_X1 U591 ( .A(G85GAT), .B(KEYINPUT107), .ZN(n526) );
  XNOR2_X1 U592 ( .A(n527), .B(n526), .ZN(G1336GAT) );
  NOR2_X1 U593 ( .A1(n528), .A2(n533), .ZN(n529) );
  XOR2_X1 U594 ( .A(KEYINPUT108), .B(n529), .Z(n530) );
  XNOR2_X1 U595 ( .A(G92GAT), .B(n530), .ZN(G1337GAT) );
  NOR2_X1 U596 ( .A1(n531), .A2(n533), .ZN(n532) );
  XOR2_X1 U597 ( .A(G99GAT), .B(n532), .Z(G1338GAT) );
  NOR2_X1 U598 ( .A1(n534), .A2(n533), .ZN(n536) );
  XNOR2_X1 U599 ( .A(KEYINPUT109), .B(KEYINPUT44), .ZN(n535) );
  XNOR2_X1 U600 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U601 ( .A(G106GAT), .B(n537), .ZN(G1339GAT) );
  XNOR2_X1 U602 ( .A(G113GAT), .B(KEYINPUT112), .ZN(n539) );
  NAND2_X1 U603 ( .A1(n544), .A2(n577), .ZN(n538) );
  XNOR2_X1 U604 ( .A(n539), .B(n538), .ZN(G1340GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT49), .B(KEYINPUT113), .Z(n541) );
  INV_X1 U606 ( .A(n555), .ZN(n569) );
  NAND2_X1 U607 ( .A1(n544), .A2(n569), .ZN(n540) );
  XNOR2_X1 U608 ( .A(n541), .B(n540), .ZN(n542) );
  XOR2_X1 U609 ( .A(G120GAT), .B(n542), .Z(G1341GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n546) );
  NAND2_X1 U611 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(n548) );
  XOR2_X1 U613 ( .A(G134GAT), .B(KEYINPUT116), .Z(n547) );
  XNOR2_X1 U614 ( .A(n548), .B(n547), .ZN(G1343GAT) );
  NAND2_X1 U615 ( .A1(n574), .A2(n549), .ZN(n560) );
  NOR2_X1 U616 ( .A1(n550), .A2(n560), .ZN(n552) );
  XNOR2_X1 U617 ( .A(G141GAT), .B(KEYINPUT117), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n552), .B(n551), .ZN(G1344GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT118), .B(KEYINPUT52), .Z(n554) );
  XNOR2_X1 U620 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n553) );
  XNOR2_X1 U621 ( .A(n554), .B(n553), .ZN(n557) );
  NOR2_X1 U622 ( .A1(n555), .A2(n560), .ZN(n556) );
  XOR2_X1 U623 ( .A(n557), .B(n556), .Z(G1345GAT) );
  NOR2_X1 U624 ( .A1(n558), .A2(n560), .ZN(n559) );
  XOR2_X1 U625 ( .A(G155GAT), .B(n559), .Z(G1346GAT) );
  NOR2_X1 U626 ( .A1(n561), .A2(n560), .ZN(n563) );
  XNOR2_X1 U627 ( .A(G162GAT), .B(KEYINPUT119), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n563), .B(n562), .ZN(G1347GAT) );
  XOR2_X1 U629 ( .A(G169GAT), .B(KEYINPUT121), .Z(n565) );
  NAND2_X1 U630 ( .A1(n572), .A2(n577), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(G1348GAT) );
  XOR2_X1 U632 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n567) );
  XNOR2_X1 U633 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n566) );
  XNOR2_X1 U634 ( .A(n567), .B(n566), .ZN(n568) );
  XOR2_X1 U635 ( .A(KEYINPUT56), .B(n568), .Z(n571) );
  NAND2_X1 U636 ( .A1(n572), .A2(n569), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(G1349GAT) );
  NAND2_X1 U638 ( .A1(n572), .A2(n585), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n573), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U640 ( .A(KEYINPUT59), .B(KEYINPUT124), .ZN(n581) );
  XOR2_X1 U641 ( .A(G197GAT), .B(KEYINPUT60), .Z(n579) );
  INV_X1 U642 ( .A(n574), .ZN(n575) );
  NOR2_X1 U643 ( .A1(n576), .A2(n575), .ZN(n589) );
  NAND2_X1 U644 ( .A1(n589), .A2(n577), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1352GAT) );
  XOR2_X1 U647 ( .A(G204GAT), .B(KEYINPUT61), .Z(n584) );
  NAND2_X1 U648 ( .A1(n589), .A2(n582), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(G1353GAT) );
  XOR2_X1 U650 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n587) );
  NAND2_X1 U651 ( .A1(n589), .A2(n585), .ZN(n586) );
  XNOR2_X1 U652 ( .A(n587), .B(n586), .ZN(n588) );
  XNOR2_X1 U653 ( .A(G211GAT), .B(n588), .ZN(G1354GAT) );
  INV_X1 U654 ( .A(n589), .ZN(n590) );
  NOR2_X1 U655 ( .A1(n591), .A2(n590), .ZN(n593) );
  XNOR2_X1 U656 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n592) );
  XNOR2_X1 U657 ( .A(n593), .B(n592), .ZN(n594) );
  XNOR2_X1 U658 ( .A(G218GAT), .B(n594), .ZN(G1355GAT) );
endmodule

