

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748;

  INV_X1 U368 ( .A(G902), .ZN(n465) );
  INV_X1 U369 ( .A(G237), .ZN(n464) );
  XNOR2_X1 U370 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n453) );
  XNOR2_X1 U371 ( .A(G107), .B(G104), .ZN(n452) );
  INV_X1 U372 ( .A(G140), .ZN(n413) );
  NAND2_X1 U373 ( .A1(G234), .A2(G237), .ZN(n469) );
  XNOR2_X1 U374 ( .A(G119), .B(KEYINPUT24), .ZN(n498) );
  XNOR2_X1 U375 ( .A(G122), .B(KEYINPUT12), .ZN(n435) );
  INV_X2 U376 ( .A(n716), .ZN(n399) );
  INV_X2 U377 ( .A(KEYINPUT66), .ZN(n617) );
  XOR2_X2 U378 ( .A(n630), .B(n633), .Z(n362) );
  INV_X2 U379 ( .A(KEYINPUT73), .ZN(n425) );
  XOR2_X2 U380 ( .A(KEYINPUT62), .B(n618), .Z(n363) );
  XOR2_X1 U381 ( .A(KEYINPUT101), .B(KEYINPUT11), .Z(n436) );
  XOR2_X1 U382 ( .A(KEYINPUT100), .B(KEYINPUT99), .Z(n439) );
  AND2_X1 U383 ( .A1(n736), .A2(KEYINPUT2), .ZN(n401) );
  XOR2_X1 U384 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n427) );
  NOR2_X2 U385 ( .A1(n624), .A2(G902), .ZN(n445) );
  XNOR2_X2 U386 ( .A(n445), .B(n444), .ZN(n545) );
  INV_X2 U387 ( .A(G953), .ZN(n740) );
  INV_X1 U388 ( .A(n579), .ZN(n569) );
  XNOR2_X1 U389 ( .A(n579), .B(n516), .ZN(n560) );
  INV_X1 U390 ( .A(KEYINPUT110), .ZN(n347) );
  INV_X1 U391 ( .A(KEYINPUT109), .ZN(n348) );
  OR2_X1 U392 ( .A1(n698), .A2(n424), .ZN(n699) );
  NOR2_X1 U393 ( .A1(n605), .A2(n412), .ZN(n411) );
  NOR2_X1 U394 ( .A1(n532), .A2(KEYINPUT44), .ZN(n528) );
  XNOR2_X1 U395 ( .A(n365), .B(KEYINPUT32), .ZN(n747) );
  NOR2_X1 U396 ( .A1(n606), .A2(n609), .ZN(n567) );
  XNOR2_X1 U397 ( .A(n521), .B(KEYINPUT33), .ZN(n685) );
  NOR2_X1 U398 ( .A1(n563), .A2(n562), .ZN(n564) );
  NAND2_X1 U399 ( .A1(n417), .A2(n416), .ZN(n415) );
  XNOR2_X1 U400 ( .A(n561), .B(n347), .ZN(n562) );
  XNOR2_X1 U401 ( .A(n537), .B(n348), .ZN(n520) );
  NOR2_X2 U402 ( .A1(n581), .A2(n582), .ZN(n407) );
  NOR2_X1 U403 ( .A1(n570), .A2(n569), .ZN(n571) );
  NOR2_X1 U404 ( .A1(n570), .A2(n560), .ZN(n561) );
  XNOR2_X1 U405 ( .A(n383), .B(G469), .ZN(n573) );
  NOR2_X1 U406 ( .A1(n710), .A2(G902), .ZN(n544) );
  NOR2_X1 U407 ( .A1(n707), .A2(G902), .ZN(n383) );
  XNOR2_X1 U408 ( .A(n369), .B(n367), .ZN(n710) );
  XNOR2_X1 U409 ( .A(n378), .B(n495), .ZN(n707) );
  XNOR2_X1 U410 ( .A(n732), .B(G101), .ZN(n349) );
  XNOR2_X1 U411 ( .A(n431), .B(n430), .ZN(n460) );
  XNOR2_X1 U412 ( .A(n731), .B(G146), .ZN(n504) );
  XNOR2_X1 U413 ( .A(n429), .B(KEYINPUT79), .ZN(n431) );
  XNOR2_X1 U414 ( .A(n414), .B(n413), .ZN(n731) );
  XNOR2_X1 U415 ( .A(n427), .B(n426), .ZN(n370) );
  XNOR2_X1 U416 ( .A(KEYINPUT10), .B(G125), .ZN(n414) );
  NOR2_X2 U417 ( .A1(G953), .A2(G237), .ZN(n484) );
  XNOR2_X2 U418 ( .A(G128), .B(G137), .ZN(n500) );
  XNOR2_X2 U419 ( .A(KEYINPUT16), .B(G122), .ZN(n450) );
  XNOR2_X2 U420 ( .A(G134), .B(G116), .ZN(n428) );
  INV_X1 U421 ( .A(KEYINPUT65), .ZN(n429) );
  XNOR2_X1 U422 ( .A(KEYINPUT23), .B(KEYINPUT78), .ZN(n497) );
  XNOR2_X1 U423 ( .A(G107), .B(KEYINPUT104), .ZN(n426) );
  XNOR2_X1 U424 ( .A(G143), .B(G128), .ZN(n430) );
  XNOR2_X1 U425 ( .A(n346), .B(n480), .ZN(n618) );
  XNOR2_X1 U426 ( .A(n487), .B(n732), .ZN(n346) );
  XNOR2_X1 U427 ( .A(n423), .B(n477), .ZN(n522) );
  XNOR2_X1 U428 ( .A(n735), .B(n349), .ZN(n378) );
  XNOR2_X2 U429 ( .A(n350), .B(n494), .ZN(n724) );
  XNOR2_X2 U430 ( .A(n481), .B(n450), .ZN(n350) );
  XNOR2_X2 U431 ( .A(n352), .B(n351), .ZN(n481) );
  XNOR2_X2 U432 ( .A(G119), .B(KEYINPUT3), .ZN(n351) );
  XNOR2_X2 U433 ( .A(G116), .B(G113), .ZN(n352) );
  BUF_X1 U434 ( .A(n384), .Z(n353) );
  XNOR2_X1 U435 ( .A(n478), .B(n385), .ZN(n384) );
  BUF_X1 U436 ( .A(n622), .Z(n354) );
  BUF_X1 U437 ( .A(n616), .Z(n355) );
  BUF_X1 U438 ( .A(n373), .Z(n356) );
  XNOR2_X1 U439 ( .A(n366), .B(KEYINPUT108), .ZN(n622) );
  INV_X1 U440 ( .A(KEYINPUT107), .ZN(n420) );
  INV_X1 U441 ( .A(KEYINPUT81), .ZN(n402) );
  NAND2_X1 U442 ( .A1(n520), .A2(n519), .ZN(n521) );
  INV_X1 U443 ( .A(KEYINPUT111), .ZN(n574) );
  XNOR2_X1 U444 ( .A(n583), .B(KEYINPUT39), .ZN(n611) );
  INV_X1 U445 ( .A(KEYINPUT22), .ZN(n385) );
  NAND2_X1 U446 ( .A1(n522), .A2(n422), .ZN(n478) );
  NAND2_X1 U447 ( .A1(n418), .A2(n415), .ZN(n422) );
  XNOR2_X1 U448 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U449 ( .A(n460), .B(n368), .ZN(n367) );
  XNOR2_X1 U450 ( .A(n371), .B(n370), .ZN(n369) );
  XNOR2_X1 U451 ( .A(n428), .B(G122), .ZN(n368) );
  XOR2_X1 U452 ( .A(KEYINPUT97), .B(KEYINPUT5), .Z(n483) );
  AND2_X1 U453 ( .A1(n659), .A2(n420), .ZN(n416) );
  XOR2_X1 U454 ( .A(KEYINPUT25), .B(KEYINPUT77), .Z(n510) );
  INV_X1 U455 ( .A(KEYINPUT48), .ZN(n408) );
  XNOR2_X1 U456 ( .A(n500), .B(G110), .ZN(n501) );
  XNOR2_X1 U457 ( .A(n432), .B(n372), .ZN(n505) );
  INV_X1 U458 ( .A(KEYINPUT8), .ZN(n372) );
  NAND2_X1 U459 ( .A1(n505), .A2(G217), .ZN(n371) );
  XNOR2_X2 U460 ( .A(G137), .B(G134), .ZN(n479) );
  XOR2_X1 U461 ( .A(G125), .B(KEYINPUT92), .Z(n456) );
  INV_X1 U462 ( .A(KEYINPUT74), .ZN(n403) );
  INV_X1 U463 ( .A(n625), .ZN(n392) );
  XNOR2_X1 U464 ( .A(KEYINPUT42), .B(n379), .ZN(n748) );
  NAND2_X1 U465 ( .A1(n353), .A2(n361), .ZN(n365) );
  XNOR2_X1 U466 ( .A(n714), .B(n715), .ZN(n390) );
  XNOR2_X1 U467 ( .A(n709), .B(n397), .ZN(n711) );
  XNOR2_X1 U468 ( .A(n710), .B(KEYINPUT122), .ZN(n397) );
  XNOR2_X1 U469 ( .A(n704), .B(n395), .ZN(G75) );
  XNOR2_X1 U470 ( .A(n396), .B(KEYINPUT120), .ZN(n395) );
  INV_X1 U471 ( .A(KEYINPUT53), .ZN(n396) );
  XOR2_X1 U472 ( .A(KEYINPUT76), .B(KEYINPUT19), .Z(n357) );
  NOR2_X1 U473 ( .A1(n666), .A2(n607), .ZN(n358) );
  XOR2_X1 U474 ( .A(KEYINPUT30), .B(n580), .Z(n359) );
  OR2_X1 U475 ( .A1(n659), .A2(n420), .ZN(n360) );
  AND2_X1 U476 ( .A1(n518), .A2(n607), .ZN(n361) );
  NOR2_X1 U477 ( .A1(n740), .A2(G952), .ZN(n716) );
  XNOR2_X2 U478 ( .A(n364), .B(KEYINPUT88), .ZN(n533) );
  NAND2_X1 U479 ( .A1(n622), .A2(n747), .ZN(n364) );
  NAND2_X1 U480 ( .A1(n514), .A2(n517), .ZN(n366) );
  NAND2_X1 U481 ( .A1(n373), .A2(n476), .ZN(n423) );
  NAND2_X1 U482 ( .A1(n588), .A2(n356), .ZN(n593) );
  XNOR2_X1 U483 ( .A(n468), .B(n357), .ZN(n373) );
  INV_X1 U484 ( .A(n607), .ZN(n374) );
  XNOR2_X1 U485 ( .A(n573), .B(KEYINPUT1), .ZN(n662) );
  XNOR2_X1 U486 ( .A(n463), .B(n376), .ZN(n565) );
  XNOR2_X2 U487 ( .A(n387), .B(n617), .ZN(n375) );
  NAND2_X2 U488 ( .A1(n616), .A2(n388), .ZN(n387) );
  AND2_X1 U489 ( .A1(n466), .A2(G210), .ZN(n376) );
  NAND2_X1 U490 ( .A1(n391), .A2(n399), .ZN(n628) );
  XNOR2_X1 U491 ( .A(n626), .B(n392), .ZN(n391) );
  NAND2_X1 U492 ( .A1(n393), .A2(n399), .ZN(n636) );
  XNOR2_X1 U493 ( .A(n634), .B(n362), .ZN(n393) );
  XNOR2_X1 U494 ( .A(n377), .B(n437), .ZN(n441) );
  XOR2_X1 U495 ( .A(n434), .B(n433), .Z(n377) );
  BUF_X1 U496 ( .A(n522), .Z(n543) );
  NOR2_X2 U497 ( .A1(n609), .A2(n601), .ZN(n621) );
  AND2_X1 U498 ( .A1(n673), .A2(n588), .ZN(n379) );
  INV_X1 U499 ( .A(n353), .ZN(n515) );
  NAND2_X1 U500 ( .A1(n595), .A2(n594), .ZN(n381) );
  NAND2_X1 U501 ( .A1(n380), .A2(KEYINPUT83), .ZN(n382) );
  NAND2_X1 U502 ( .A1(n381), .A2(n382), .ZN(n598) );
  INV_X1 U503 ( .A(n595), .ZN(n380) );
  BUF_X1 U504 ( .A(n579), .Z(n666) );
  BUF_X1 U505 ( .A(n724), .Z(n726) );
  AND2_X2 U506 ( .A1(n386), .A2(n615), .ZN(n388) );
  NAND2_X1 U507 ( .A1(n614), .A2(n693), .ZN(n386) );
  XNOR2_X2 U508 ( .A(n387), .B(n617), .ZN(n712) );
  XNOR2_X2 U509 ( .A(n389), .B(n425), .ZN(n616) );
  NAND2_X1 U510 ( .A1(n401), .A2(n717), .ZN(n389) );
  BUF_X2 U511 ( .A(n375), .Z(n713) );
  NOR2_X1 U512 ( .A1(n390), .A2(n716), .ZN(G66) );
  XNOR2_X1 U513 ( .A(n394), .B(n363), .ZN(n400) );
  NAND2_X1 U514 ( .A1(n375), .A2(G472), .ZN(n394) );
  XNOR2_X1 U515 ( .A(n409), .B(n408), .ZN(n613) );
  XNOR2_X1 U516 ( .A(n706), .B(n398), .ZN(n708) );
  XNOR2_X1 U517 ( .A(n707), .B(n705), .ZN(n398) );
  NAND2_X1 U518 ( .A1(n400), .A2(n399), .ZN(n619) );
  XNOR2_X2 U519 ( .A(n554), .B(KEYINPUT45), .ZN(n717) );
  NAND2_X1 U520 ( .A1(n717), .A2(n736), .ZN(n614) );
  NAND2_X1 U521 ( .A1(n614), .A2(n402), .ZN(n694) );
  XNOR2_X2 U522 ( .A(n404), .B(n403), .ZN(n599) );
  NAND2_X1 U523 ( .A1(n359), .A2(n405), .ZN(n404) );
  XNOR2_X1 U524 ( .A(n407), .B(n406), .ZN(n405) );
  INV_X1 U525 ( .A(KEYINPUT75), .ZN(n406) );
  NAND2_X1 U526 ( .A1(n411), .A2(n410), .ZN(n409) );
  XNOR2_X1 U527 ( .A(n591), .B(n590), .ZN(n410) );
  INV_X1 U528 ( .A(n592), .ZN(n412) );
  INV_X1 U529 ( .A(n678), .ZN(n417) );
  INV_X1 U530 ( .A(n419), .ZN(n418) );
  NAND2_X1 U531 ( .A1(n421), .A2(n360), .ZN(n419) );
  NAND2_X1 U532 ( .A1(n678), .A2(KEYINPUT107), .ZN(n421) );
  INV_X1 U533 ( .A(n355), .ZN(n424) );
  INV_X1 U534 ( .A(KEYINPUT83), .ZN(n594) );
  BUF_X1 U535 ( .A(n540), .Z(n663) );
  XNOR2_X1 U536 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U537 ( .A(n575), .B(n574), .ZN(n588) );
  BUF_X1 U538 ( .A(n532), .Z(n746) );
  NAND2_X1 U539 ( .A1(G234), .A2(n740), .ZN(n432) );
  XNOR2_X1 U540 ( .A(n544), .B(G478), .ZN(n525) );
  XOR2_X1 U541 ( .A(G104), .B(G113), .Z(n434) );
  XNOR2_X1 U542 ( .A(G143), .B(G131), .ZN(n433) );
  XNOR2_X1 U543 ( .A(n436), .B(n435), .ZN(n437) );
  NAND2_X1 U544 ( .A1(G214), .A2(n484), .ZN(n438) );
  XNOR2_X1 U545 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U546 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U547 ( .A(n504), .B(n442), .ZN(n624) );
  XOR2_X1 U548 ( .A(G475), .B(KEYINPUT102), .Z(n443) );
  XNOR2_X1 U549 ( .A(KEYINPUT13), .B(n443), .ZN(n444) );
  NAND2_X1 U550 ( .A1(n525), .A2(n545), .ZN(n446) );
  XNOR2_X2 U551 ( .A(n446), .B(KEYINPUT106), .ZN(n678) );
  XNOR2_X1 U552 ( .A(G902), .B(KEYINPUT90), .ZN(n447) );
  XNOR2_X1 U553 ( .A(n447), .B(KEYINPUT15), .ZN(n462) );
  NAND2_X1 U554 ( .A1(n462), .A2(G234), .ZN(n448) );
  XNOR2_X1 U555 ( .A(KEYINPUT20), .B(n448), .ZN(n508) );
  NAND2_X1 U556 ( .A1(n508), .A2(G221), .ZN(n449) );
  XOR2_X1 U557 ( .A(KEYINPUT21), .B(n449), .Z(n659) );
  XNOR2_X1 U558 ( .A(KEYINPUT91), .B(G110), .ZN(n451) );
  XNOR2_X1 U559 ( .A(n452), .B(n451), .ZN(n494) );
  NAND2_X1 U560 ( .A1(G224), .A2(n740), .ZN(n454) );
  XNOR2_X1 U561 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U562 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U563 ( .A(n724), .B(n457), .ZN(n461) );
  XNOR2_X2 U564 ( .A(KEYINPUT4), .B(G146), .ZN(n458) );
  XNOR2_X1 U565 ( .A(n458), .B(KEYINPUT69), .ZN(n459) );
  XNOR2_X2 U566 ( .A(n460), .B(n459), .ZN(n735) );
  XNOR2_X2 U567 ( .A(n735), .B(G101), .ZN(n480) );
  XNOR2_X1 U568 ( .A(n461), .B(n480), .ZN(n629) );
  INV_X1 U569 ( .A(n462), .ZN(n615) );
  NOR2_X1 U570 ( .A1(n629), .A2(n615), .ZN(n463) );
  NAND2_X1 U571 ( .A1(n465), .A2(n464), .ZN(n466) );
  NAND2_X1 U572 ( .A1(n466), .A2(G214), .ZN(n680) );
  INV_X1 U573 ( .A(n680), .ZN(n467) );
  NOR2_X2 U574 ( .A1(n565), .A2(n467), .ZN(n468) );
  XNOR2_X1 U575 ( .A(n469), .B(KEYINPUT14), .ZN(n473) );
  NAND2_X1 U576 ( .A1(n473), .A2(G902), .ZN(n470) );
  XNOR2_X1 U577 ( .A(KEYINPUT94), .B(n470), .ZN(n555) );
  NOR2_X1 U578 ( .A1(G898), .A2(n740), .ZN(n471) );
  XNOR2_X1 U579 ( .A(KEYINPUT93), .B(n471), .ZN(n727) );
  NOR2_X1 U580 ( .A1(n555), .A2(n727), .ZN(n472) );
  XNOR2_X1 U581 ( .A(n472), .B(KEYINPUT95), .ZN(n475) );
  NAND2_X1 U582 ( .A1(G952), .A2(n473), .ZN(n692) );
  NOR2_X1 U583 ( .A1(n692), .A2(G953), .ZN(n558) );
  INV_X1 U584 ( .A(n558), .ZN(n474) );
  NAND2_X1 U585 ( .A1(n475), .A2(n474), .ZN(n476) );
  INV_X1 U586 ( .A(KEYINPUT0), .ZN(n477) );
  XNOR2_X1 U587 ( .A(n479), .B(G131), .ZN(n732) );
  BUF_X1 U588 ( .A(n481), .Z(n482) );
  XNOR2_X1 U589 ( .A(n482), .B(n483), .ZN(n486) );
  NAND2_X1 U590 ( .A1(n484), .A2(G210), .ZN(n485) );
  NOR2_X1 U591 ( .A1(n618), .A2(G902), .ZN(n491) );
  XNOR2_X1 U592 ( .A(KEYINPUT72), .B(KEYINPUT98), .ZN(n489) );
  INV_X1 U593 ( .A(G472), .ZN(n488) );
  XNOR2_X1 U594 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X2 U595 ( .A(n491), .B(n490), .ZN(n579) );
  NAND2_X1 U596 ( .A1(G227), .A2(n740), .ZN(n492) );
  XNOR2_X1 U597 ( .A(n492), .B(G140), .ZN(n493) );
  XNOR2_X1 U598 ( .A(n494), .B(n493), .ZN(n495) );
  INV_X1 U599 ( .A(n662), .ZN(n607) );
  NAND2_X1 U600 ( .A1(n384), .A2(n358), .ZN(n496) );
  XNOR2_X1 U601 ( .A(n496), .B(KEYINPUT67), .ZN(n514) );
  INV_X1 U602 ( .A(n497), .ZN(n499) );
  XNOR2_X1 U603 ( .A(n499), .B(n498), .ZN(n502) );
  XNOR2_X1 U604 ( .A(n504), .B(n503), .ZN(n507) );
  NAND2_X1 U605 ( .A1(G221), .A2(n505), .ZN(n506) );
  XNOR2_X1 U606 ( .A(n507), .B(n506), .ZN(n715) );
  NOR2_X1 U607 ( .A1(n715), .A2(G902), .ZN(n513) );
  NAND2_X1 U608 ( .A1(n508), .A2(G217), .ZN(n509) );
  XNOR2_X1 U609 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U610 ( .A(n511), .B(KEYINPUT96), .ZN(n512) );
  XNOR2_X2 U611 ( .A(n513), .B(n512), .ZN(n658) );
  INV_X1 U612 ( .A(n658), .ZN(n517) );
  XOR2_X1 U613 ( .A(KEYINPUT6), .B(KEYINPUT105), .Z(n516) );
  AND2_X1 U614 ( .A1(n560), .A2(n517), .ZN(n518) );
  XNOR2_X1 U615 ( .A(n533), .B(KEYINPUT87), .ZN(n530) );
  NAND2_X1 U616 ( .A1(n659), .A2(n658), .ZN(n540) );
  NOR2_X2 U617 ( .A1(n662), .A2(n663), .ZN(n537) );
  INV_X1 U618 ( .A(n560), .ZN(n519) );
  NAND2_X1 U619 ( .A1(n685), .A2(n543), .ZN(n524) );
  XNOR2_X1 U620 ( .A(KEYINPUT71), .B(KEYINPUT34), .ZN(n523) );
  XNOR2_X1 U621 ( .A(n524), .B(n523), .ZN(n526) );
  NOR2_X1 U622 ( .A1(n525), .A2(n545), .ZN(n600) );
  NAND2_X1 U623 ( .A1(n526), .A2(n600), .ZN(n527) );
  XNOR2_X1 U624 ( .A(n527), .B(KEYINPUT35), .ZN(n532) );
  XNOR2_X1 U625 ( .A(n528), .B(KEYINPUT68), .ZN(n529) );
  NAND2_X1 U626 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U627 ( .A(n531), .B(KEYINPUT70), .ZN(n553) );
  OR2_X1 U628 ( .A1(n746), .A2(n533), .ZN(n534) );
  NAND2_X1 U629 ( .A1(n534), .A2(KEYINPUT44), .ZN(n551) );
  AND2_X1 U630 ( .A1(n560), .A2(n658), .ZN(n535) );
  NAND2_X1 U631 ( .A1(n535), .A2(n374), .ZN(n536) );
  OR2_X1 U632 ( .A1(n515), .A2(n536), .ZN(n637) );
  NAND2_X1 U633 ( .A1(n666), .A2(n537), .ZN(n669) );
  INV_X1 U634 ( .A(n543), .ZN(n538) );
  OR2_X1 U635 ( .A1(n669), .A2(n538), .ZN(n539) );
  XNOR2_X1 U636 ( .A(n539), .B(KEYINPUT31), .ZN(n653) );
  OR2_X2 U637 ( .A1(n573), .A2(n540), .ZN(n581) );
  OR2_X1 U638 ( .A1(n666), .A2(n581), .ZN(n541) );
  INV_X1 U639 ( .A(n541), .ZN(n542) );
  AND2_X1 U640 ( .A1(n543), .A2(n542), .ZN(n639) );
  OR2_X1 U641 ( .A1(n653), .A2(n639), .ZN(n548) );
  XOR2_X1 U642 ( .A(n544), .B(G478), .Z(n547) );
  XOR2_X1 U643 ( .A(n545), .B(KEYINPUT103), .Z(n546) );
  NOR2_X1 U644 ( .A1(n547), .A2(n546), .ZN(n649) );
  AND2_X1 U645 ( .A1(n547), .A2(n546), .ZN(n652) );
  OR2_X1 U646 ( .A1(n649), .A2(n652), .ZN(n677) );
  NAND2_X1 U647 ( .A1(n548), .A2(n677), .ZN(n549) );
  AND2_X1 U648 ( .A1(n637), .A2(n549), .ZN(n550) );
  AND2_X1 U649 ( .A1(n551), .A2(n550), .ZN(n552) );
  NAND2_X1 U650 ( .A1(n553), .A2(n552), .ZN(n554) );
  INV_X1 U651 ( .A(n649), .ZN(n563) );
  OR2_X1 U652 ( .A1(n555), .A2(n740), .ZN(n556) );
  NOR2_X1 U653 ( .A1(G900), .A2(n556), .ZN(n557) );
  NOR2_X1 U654 ( .A1(n558), .A2(n557), .ZN(n582) );
  NOR2_X1 U655 ( .A1(n658), .A2(n582), .ZN(n559) );
  NAND2_X1 U656 ( .A1(n559), .A2(n659), .ZN(n570) );
  NAND2_X1 U657 ( .A1(n564), .A2(n680), .ZN(n606) );
  BUF_X1 U658 ( .A(n565), .Z(n609) );
  INV_X1 U659 ( .A(KEYINPUT36), .ZN(n566) );
  XNOR2_X1 U660 ( .A(n567), .B(n566), .ZN(n568) );
  NOR2_X1 U661 ( .A1(n374), .A2(n568), .ZN(n655) );
  XNOR2_X1 U662 ( .A(n655), .B(KEYINPUT86), .ZN(n578) );
  XOR2_X1 U663 ( .A(KEYINPUT28), .B(n571), .Z(n572) );
  NOR2_X1 U664 ( .A1(n573), .A2(n572), .ZN(n575) );
  INV_X1 U665 ( .A(n593), .ZN(n646) );
  NAND2_X1 U666 ( .A1(n646), .A2(n677), .ZN(n576) );
  NOR2_X1 U667 ( .A1(n576), .A2(KEYINPUT47), .ZN(n577) );
  NOR2_X1 U668 ( .A1(n578), .A2(n577), .ZN(n592) );
  XOR2_X1 U669 ( .A(KEYINPUT40), .B(KEYINPUT112), .Z(n585) );
  NAND2_X1 U670 ( .A1(n579), .A2(n680), .ZN(n580) );
  XNOR2_X1 U671 ( .A(n609), .B(KEYINPUT38), .ZN(n676) );
  NAND2_X1 U672 ( .A1(n599), .A2(n676), .ZN(n583) );
  NAND2_X1 U673 ( .A1(n611), .A2(n649), .ZN(n584) );
  XNOR2_X1 U674 ( .A(n585), .B(n584), .ZN(n745) );
  INV_X1 U675 ( .A(n676), .ZN(n586) );
  NOR2_X1 U676 ( .A1(n678), .A2(n586), .ZN(n675) );
  NAND2_X1 U677 ( .A1(n680), .A2(n675), .ZN(n587) );
  XNOR2_X1 U678 ( .A(n587), .B(KEYINPUT41), .ZN(n673) );
  NOR2_X1 U679 ( .A1(n745), .A2(n748), .ZN(n591) );
  XOR2_X1 U680 ( .A(KEYINPUT46), .B(KEYINPUT85), .Z(n589) );
  XNOR2_X1 U681 ( .A(KEYINPUT64), .B(n589), .ZN(n590) );
  NAND2_X1 U682 ( .A1(n593), .A2(KEYINPUT47), .ZN(n595) );
  INV_X1 U683 ( .A(n677), .ZN(n596) );
  NAND2_X1 U684 ( .A1(n596), .A2(KEYINPUT47), .ZN(n597) );
  NAND2_X1 U685 ( .A1(n598), .A2(n597), .ZN(n603) );
  NAND2_X1 U686 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U687 ( .A(n621), .B(KEYINPUT84), .ZN(n602) );
  NOR2_X1 U688 ( .A1(n603), .A2(n602), .ZN(n604) );
  XOR2_X1 U689 ( .A(n604), .B(KEYINPUT82), .Z(n605) );
  NOR2_X1 U690 ( .A1(n607), .A2(n606), .ZN(n608) );
  XOR2_X1 U691 ( .A(n608), .B(KEYINPUT43), .Z(n610) );
  NAND2_X1 U692 ( .A1(n610), .A2(n609), .ZN(n620) );
  NAND2_X1 U693 ( .A1(n611), .A2(n652), .ZN(n657) );
  AND2_X1 U694 ( .A1(n620), .A2(n657), .ZN(n612) );
  AND2_X2 U695 ( .A1(n613), .A2(n612), .ZN(n736) );
  INV_X1 U696 ( .A(KEYINPUT2), .ZN(n693) );
  XNOR2_X1 U697 ( .A(n619), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U698 ( .A(n620), .B(G140), .ZN(G42) );
  XOR2_X1 U699 ( .A(G143), .B(n621), .Z(G45) );
  XNOR2_X1 U700 ( .A(n354), .B(G110), .ZN(G12) );
  NAND2_X1 U701 ( .A1(n712), .A2(G475), .ZN(n626) );
  XNOR2_X1 U702 ( .A(KEYINPUT121), .B(KEYINPUT59), .ZN(n623) );
  XNOR2_X1 U703 ( .A(n624), .B(n623), .ZN(n625) );
  INV_X1 U704 ( .A(KEYINPUT60), .ZN(n627) );
  XNOR2_X1 U705 ( .A(n628), .B(n627), .ZN(G60) );
  NAND2_X1 U706 ( .A1(n712), .A2(G210), .ZN(n634) );
  BUF_X1 U707 ( .A(n629), .Z(n630) );
  XNOR2_X1 U708 ( .A(KEYINPUT89), .B(KEYINPUT54), .ZN(n632) );
  XNOR2_X1 U709 ( .A(KEYINPUT55), .B(KEYINPUT80), .ZN(n631) );
  XNOR2_X1 U710 ( .A(n632), .B(n631), .ZN(n633) );
  INV_X1 U711 ( .A(KEYINPUT56), .ZN(n635) );
  XNOR2_X1 U712 ( .A(n636), .B(n635), .ZN(G51) );
  XNOR2_X1 U713 ( .A(G101), .B(n637), .ZN(G3) );
  NAND2_X1 U714 ( .A1(n639), .A2(n649), .ZN(n638) );
  XNOR2_X1 U715 ( .A(n638), .B(G104), .ZN(G6) );
  XOR2_X1 U716 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n641) );
  NAND2_X1 U717 ( .A1(n639), .A2(n652), .ZN(n640) );
  XNOR2_X1 U718 ( .A(n641), .B(n640), .ZN(n642) );
  XNOR2_X1 U719 ( .A(G107), .B(n642), .ZN(G9) );
  XOR2_X1 U720 ( .A(KEYINPUT29), .B(KEYINPUT113), .Z(n644) );
  NAND2_X1 U721 ( .A1(n646), .A2(n652), .ZN(n643) );
  XNOR2_X1 U722 ( .A(n644), .B(n643), .ZN(n645) );
  XOR2_X1 U723 ( .A(G128), .B(n645), .Z(G30) );
  NAND2_X1 U724 ( .A1(n646), .A2(n649), .ZN(n647) );
  XNOR2_X1 U725 ( .A(n647), .B(KEYINPUT114), .ZN(n648) );
  XNOR2_X1 U726 ( .A(G146), .B(n648), .ZN(G48) );
  XOR2_X1 U727 ( .A(G113), .B(KEYINPUT115), .Z(n651) );
  NAND2_X1 U728 ( .A1(n653), .A2(n649), .ZN(n650) );
  XNOR2_X1 U729 ( .A(n651), .B(n650), .ZN(G15) );
  NAND2_X1 U730 ( .A1(n653), .A2(n652), .ZN(n654) );
  XNOR2_X1 U731 ( .A(n654), .B(G116), .ZN(G18) );
  XNOR2_X1 U732 ( .A(n655), .B(G125), .ZN(n656) );
  XNOR2_X1 U733 ( .A(n656), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U734 ( .A(G134), .B(n657), .ZN(G36) );
  NAND2_X1 U735 ( .A1(n685), .A2(n673), .ZN(n703) );
  NOR2_X1 U736 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U737 ( .A(n660), .B(KEYINPUT49), .ZN(n661) );
  XNOR2_X1 U738 ( .A(n661), .B(KEYINPUT116), .ZN(n668) );
  AND2_X1 U739 ( .A1(n663), .A2(n374), .ZN(n664) );
  XNOR2_X1 U740 ( .A(n664), .B(KEYINPUT50), .ZN(n665) );
  NOR2_X1 U741 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U742 ( .A1(n668), .A2(n667), .ZN(n670) );
  NAND2_X1 U743 ( .A1(n670), .A2(n669), .ZN(n671) );
  XOR2_X1 U744 ( .A(KEYINPUT51), .B(n671), .Z(n672) );
  NAND2_X1 U745 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U746 ( .A(KEYINPUT117), .B(n674), .ZN(n688) );
  INV_X1 U747 ( .A(n675), .ZN(n683) );
  NAND2_X1 U748 ( .A1(n677), .A2(n676), .ZN(n679) );
  NAND2_X1 U749 ( .A1(n679), .A2(n678), .ZN(n681) );
  NAND2_X1 U750 ( .A1(n681), .A2(n680), .ZN(n682) );
  NAND2_X1 U751 ( .A1(n683), .A2(n682), .ZN(n684) );
  NAND2_X1 U752 ( .A1(n685), .A2(n684), .ZN(n686) );
  XOR2_X1 U753 ( .A(n686), .B(KEYINPUT118), .Z(n687) );
  NOR2_X1 U754 ( .A1(n688), .A2(n687), .ZN(n689) );
  XOR2_X1 U755 ( .A(KEYINPUT52), .B(n689), .Z(n690) );
  XNOR2_X1 U756 ( .A(n690), .B(KEYINPUT119), .ZN(n691) );
  NOR2_X1 U757 ( .A1(n692), .A2(n691), .ZN(n701) );
  NAND2_X1 U758 ( .A1(n694), .A2(n693), .ZN(n697) );
  NAND2_X1 U759 ( .A1(n425), .A2(KEYINPUT81), .ZN(n695) );
  NAND2_X1 U760 ( .A1(n695), .A2(KEYINPUT2), .ZN(n696) );
  AND2_X1 U761 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U762 ( .A1(n740), .A2(n699), .ZN(n700) );
  NOR2_X1 U763 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U764 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U765 ( .A1(n713), .A2(G469), .ZN(n706) );
  XOR2_X1 U766 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n705) );
  NOR2_X1 U767 ( .A1(n716), .A2(n708), .ZN(G54) );
  NAND2_X1 U768 ( .A1(n713), .A2(G478), .ZN(n709) );
  NOR2_X1 U769 ( .A1(n711), .A2(n716), .ZN(G63) );
  NAND2_X1 U770 ( .A1(n713), .A2(G217), .ZN(n714) );
  BUF_X1 U771 ( .A(n717), .Z(n718) );
  NAND2_X1 U772 ( .A1(n718), .A2(n740), .ZN(n723) );
  XOR2_X1 U773 ( .A(KEYINPUT61), .B(KEYINPUT123), .Z(n720) );
  NAND2_X1 U774 ( .A1(G224), .A2(G953), .ZN(n719) );
  XNOR2_X1 U775 ( .A(n720), .B(n719), .ZN(n721) );
  NAND2_X1 U776 ( .A1(n721), .A2(G898), .ZN(n722) );
  NAND2_X1 U777 ( .A1(n723), .A2(n722), .ZN(n730) );
  XNOR2_X1 U778 ( .A(G101), .B(KEYINPUT124), .ZN(n725) );
  XNOR2_X1 U779 ( .A(n726), .B(n725), .ZN(n728) );
  NAND2_X1 U780 ( .A1(n728), .A2(n727), .ZN(n729) );
  XOR2_X1 U781 ( .A(n730), .B(n729), .Z(G69) );
  XNOR2_X1 U782 ( .A(n731), .B(KEYINPUT125), .ZN(n733) );
  XNOR2_X1 U783 ( .A(n733), .B(n732), .ZN(n734) );
  XOR2_X1 U784 ( .A(n735), .B(n734), .Z(n738) );
  XOR2_X1 U785 ( .A(n736), .B(n738), .Z(n737) );
  NOR2_X1 U786 ( .A1(G953), .A2(n737), .ZN(n743) );
  XNOR2_X1 U787 ( .A(G227), .B(n738), .ZN(n739) );
  NAND2_X1 U788 ( .A1(n739), .A2(G900), .ZN(n741) );
  NOR2_X1 U789 ( .A1(n741), .A2(n740), .ZN(n742) );
  NOR2_X1 U790 ( .A1(n743), .A2(n742), .ZN(n744) );
  XNOR2_X1 U791 ( .A(KEYINPUT126), .B(n744), .ZN(G72) );
  XOR2_X1 U792 ( .A(G131), .B(n745), .Z(G33) );
  XOR2_X1 U793 ( .A(n746), .B(G122), .Z(G24) );
  XNOR2_X1 U794 ( .A(G119), .B(n747), .ZN(G21) );
  XOR2_X1 U795 ( .A(G137), .B(n748), .Z(G39) );
endmodule

