//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 0 1 1 0 0 1 0 0 1 0 1 0 0 1 0 1 1 1 1 0 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 0 1 1 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:51 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n555, new_n556, new_n557, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n577, new_n578, new_n579, new_n580, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n648, new_n650, new_n651, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT65), .Z(new_n447));
  XNOR2_X1  g022(.A(new_n447), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n452), .A2(new_n456), .B1(new_n457), .B2(new_n453), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT66), .Z(new_n459));
  XOR2_X1   g034(.A(new_n459), .B(KEYINPUT67), .Z(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  AND2_X1   g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  XNOR2_X1  g037(.A(new_n462), .B(KEYINPUT68), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G101), .ZN(new_n464));
  INV_X1    g039(.A(G137), .ZN(new_n465));
  AND2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  OR2_X1    g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(new_n461), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n464), .B1(new_n465), .B2(new_n469), .ZN(new_n470));
  AOI22_X1  g045(.A1(new_n468), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n471), .A2(new_n461), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n470), .A2(new_n472), .ZN(G160));
  OAI21_X1  g048(.A(G2104), .B1(new_n461), .B2(G112), .ZN(new_n474));
  INV_X1    g049(.A(G100), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n474), .B1(new_n475), .B2(new_n461), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n468), .A2(G2105), .ZN(new_n477));
  XNOR2_X1  g052(.A(new_n477), .B(KEYINPUT70), .ZN(new_n478));
  AND2_X1   g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n466), .A2(new_n467), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT69), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n481), .A2(new_n482), .ZN(new_n485));
  OR2_X1    g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AOI211_X1 g061(.A(new_n476), .B(new_n479), .C1(G136), .C2(new_n486), .ZN(G162));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n488));
  INV_X1    g063(.A(G138), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n488), .B1(new_n469), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n481), .A2(KEYINPUT4), .A3(G138), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(G114), .A2(G2104), .ZN(new_n493));
  INV_X1    g068(.A(G126), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n493), .B1(new_n480), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n462), .A2(G102), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n492), .A2(new_n498), .ZN(G164));
  INV_X1    g074(.A(G651), .ZN(new_n500));
  OAI21_X1  g075(.A(KEYINPUT6), .B1(new_n500), .B2(KEYINPUT71), .ZN(new_n501));
  NAND2_X1  g076(.A1(KEYINPUT72), .A2(G651), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT71), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n502), .A2(KEYINPUT71), .A3(KEYINPUT6), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AND2_X1   g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  NOR2_X1   g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G88), .ZN(new_n511));
  INV_X1    g086(.A(G62), .ZN(new_n512));
  OR2_X1    g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G651), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n511), .B1(new_n512), .B2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT71), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G651), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n519), .A2(KEYINPUT6), .B1(KEYINPUT71), .B2(new_n502), .ZN(new_n520));
  AND3_X1   g095(.A1(new_n502), .A2(KEYINPUT71), .A3(KEYINPUT6), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n522), .A2(G50), .B1(G75), .B2(G651), .ZN(new_n523));
  INV_X1    g098(.A(G543), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n517), .A2(new_n525), .ZN(G166));
  OAI21_X1  g101(.A(KEYINPUT73), .B1(new_n520), .B2(new_n521), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT73), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n504), .A2(new_n528), .A3(new_n505), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n524), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G51), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT7), .ZN(new_n533));
  INV_X1    g108(.A(G63), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n533), .B1(new_n516), .B2(new_n534), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n535), .B1(G89), .B2(new_n510), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n531), .A2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(new_n537), .ZN(G168));
  NAND2_X1  g113(.A1(new_n530), .A2(G52), .ZN(new_n539));
  NAND2_X1  g114(.A1(G77), .A2(G543), .ZN(new_n540));
  INV_X1    g115(.A(G64), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n540), .B1(new_n509), .B2(new_n541), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n510), .A2(G90), .B1(G651), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n539), .A2(new_n543), .ZN(G301));
  INV_X1    g119(.A(G301), .ZN(G171));
  NAND2_X1  g120(.A1(new_n530), .A2(G43), .ZN(new_n546));
  NAND2_X1  g121(.A1(G68), .A2(G543), .ZN(new_n547));
  INV_X1    g122(.A(G56), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n509), .B2(new_n548), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n510), .A2(G81), .B1(G651), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n546), .A2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(new_n557));
  XOR2_X1   g132(.A(new_n557), .B(KEYINPUT74), .Z(G188));
  NAND3_X1  g133(.A1(new_n513), .A2(KEYINPUT76), .A3(new_n514), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT76), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n560), .B1(new_n507), .B2(new_n508), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  AND2_X1   g137(.A1(new_n562), .A2(G65), .ZN(new_n563));
  AND2_X1   g138(.A1(G78), .A2(G543), .ZN(new_n564));
  OAI21_X1  g139(.A(G651), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n522), .A2(G91), .A3(new_n515), .ZN(new_n566));
  NAND2_X1  g141(.A1(KEYINPUT75), .A2(KEYINPUT9), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(new_n568));
  NOR2_X1   g143(.A1(KEYINPUT75), .A2(KEYINPUT9), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n527), .A2(new_n529), .ZN(new_n571));
  NAND2_X1  g146(.A1(G53), .A2(G543), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n570), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  AOI211_X1 g149(.A(new_n572), .B(new_n568), .C1(new_n527), .C2(new_n529), .ZN(new_n575));
  OAI211_X1 g150(.A(new_n565), .B(new_n566), .C1(new_n574), .C2(new_n575), .ZN(G299));
  INV_X1    g151(.A(KEYINPUT77), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n531), .A2(new_n536), .A3(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n577), .B1(new_n531), .B2(new_n536), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n579), .A2(new_n580), .ZN(G286));
  INV_X1    g156(.A(G166), .ZN(G303));
  OAI21_X1  g157(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n583));
  OR2_X1    g158(.A1(new_n583), .A2(KEYINPUT78), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(KEYINPUT78), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n584), .A2(new_n585), .B1(G87), .B2(new_n510), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n530), .A2(G49), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(G288));
  INV_X1    g163(.A(G61), .ZN(new_n589));
  OR3_X1    g164(.A1(new_n509), .A2(KEYINPUT79), .A3(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(new_n591));
  OAI21_X1  g166(.A(KEYINPUT79), .B1(new_n509), .B2(new_n589), .ZN(new_n592));
  INV_X1    g167(.A(G73), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n593), .B2(new_n524), .ZN(new_n594));
  OAI21_X1  g169(.A(G651), .B1(new_n591), .B2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT80), .ZN(new_n596));
  OR2_X1    g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n595), .A2(new_n596), .ZN(new_n598));
  NAND4_X1  g173(.A1(new_n522), .A2(KEYINPUT81), .A3(G48), .A4(G543), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT81), .ZN(new_n600));
  NAND2_X1  g175(.A1(G48), .A2(G543), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n506), .B2(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n599), .A2(new_n602), .B1(G86), .B2(new_n510), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n597), .A2(new_n598), .A3(new_n603), .ZN(G305));
  NAND2_X1  g179(.A1(G72), .A2(G543), .ZN(new_n605));
  INV_X1    g180(.A(G60), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n509), .B2(new_n606), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n510), .A2(G85), .B1(G651), .B2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(G47), .ZN(new_n609));
  NOR3_X1   g184(.A1(new_n520), .A2(new_n521), .A3(KEYINPUT73), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n528), .B1(new_n504), .B2(new_n505), .ZN(new_n611));
  OAI21_X1  g186(.A(G543), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n608), .B1(new_n609), .B2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT82), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n613), .B(new_n614), .ZN(G290));
  INV_X1    g190(.A(G868), .ZN(new_n616));
  NOR2_X1   g191(.A1(G301), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n562), .A2(G66), .ZN(new_n618));
  NAND2_X1  g193(.A1(G79), .A2(G543), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND4_X1  g195(.A1(new_n522), .A2(KEYINPUT10), .A3(G92), .A4(new_n515), .ZN(new_n621));
  NAND4_X1  g196(.A1(new_n504), .A2(G92), .A3(new_n515), .A4(new_n505), .ZN(new_n622));
  INV_X1    g197(.A(KEYINPUT10), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AOI22_X1  g199(.A1(G651), .A2(new_n620), .B1(new_n621), .B2(new_n624), .ZN(new_n625));
  INV_X1    g200(.A(KEYINPUT83), .ZN(new_n626));
  OAI21_X1  g201(.A(G54), .B1(new_n530), .B2(new_n626), .ZN(new_n627));
  AOI211_X1 g202(.A(KEYINPUT83), .B(new_n524), .C1(new_n527), .C2(new_n529), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n625), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n629), .A2(KEYINPUT84), .ZN(new_n630));
  INV_X1    g205(.A(new_n630), .ZN(new_n631));
  AND2_X1   g206(.A1(new_n629), .A2(KEYINPUT84), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n617), .B1(new_n634), .B2(new_n616), .ZN(G284));
  AOI21_X1  g210(.A(new_n617), .B1(new_n634), .B2(new_n616), .ZN(G321));
  NOR2_X1   g211(.A1(G286), .A2(new_n616), .ZN(new_n637));
  AOI22_X1  g212(.A1(new_n562), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n566), .B1(new_n638), .B2(new_n500), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n573), .B1(new_n610), .B2(new_n611), .ZN(new_n640));
  INV_X1    g215(.A(new_n570), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n571), .A2(new_n573), .A3(new_n567), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n639), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT85), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n637), .B1(new_n616), .B2(new_n645), .ZN(G297));
  AOI21_X1  g221(.A(new_n637), .B1(new_n616), .B2(new_n645), .ZN(G280));
  INV_X1    g222(.A(G559), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n634), .B1(new_n648), .B2(G860), .ZN(G148));
  NAND2_X1  g224(.A1(new_n551), .A2(new_n616), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n633), .A2(G559), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n650), .B1(new_n651), .B2(new_n616), .ZN(G323));
  XNOR2_X1  g227(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g228(.A1(new_n486), .A2(G135), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n478), .A2(G123), .ZN(new_n655));
  NOR2_X1   g230(.A1(G99), .A2(G2105), .ZN(new_n656));
  OAI21_X1  g231(.A(G2104), .B1(new_n461), .B2(G111), .ZN(new_n657));
  OAI211_X1 g232(.A(new_n654), .B(new_n655), .C1(new_n656), .C2(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT86), .Z(new_n659));
  INV_X1    g234(.A(G2096), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n659), .A2(new_n660), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n463), .A2(new_n468), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT12), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT13), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(G2100), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n661), .A2(new_n662), .A3(new_n666), .ZN(G156));
  XNOR2_X1  g242(.A(G2427), .B(G2438), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(G2430), .ZN(new_n669));
  XNOR2_X1  g244(.A(KEYINPUT15), .B(G2435), .ZN(new_n670));
  OR2_X1    g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n669), .A2(new_n670), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n671), .A2(KEYINPUT14), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT88), .ZN(new_n674));
  XOR2_X1   g249(.A(G1341), .B(G1348), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G2443), .B(G2446), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(G2451), .B(G2454), .Z(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT87), .B(KEYINPUT16), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n682), .A2(G14), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n678), .A2(new_n681), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(G401));
  XOR2_X1   g261(.A(G2072), .B(G2078), .Z(new_n687));
  XOR2_X1   g262(.A(G2084), .B(G2090), .Z(new_n688));
  XNOR2_X1  g263(.A(G2067), .B(G2678), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(KEYINPUT89), .B(KEYINPUT18), .Z(new_n691));
  AOI21_X1  g266(.A(new_n687), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  AND2_X1   g267(.A1(new_n690), .A2(KEYINPUT17), .ZN(new_n693));
  OR2_X1    g268(.A1(new_n688), .A2(new_n689), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n691), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  MUX2_X1   g270(.A(new_n692), .B(new_n687), .S(new_n695), .Z(new_n696));
  XNOR2_X1  g271(.A(G2096), .B(G2100), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(G227));
  XNOR2_X1  g273(.A(G1971), .B(G1976), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT19), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1961), .B(G1966), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT90), .ZN(new_n702));
  XOR2_X1   g277(.A(G1956), .B(G2474), .Z(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  XOR2_X1   g279(.A(KEYINPUT91), .B(KEYINPUT20), .Z(new_n705));
  OR2_X1    g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  OR2_X1    g281(.A1(new_n702), .A2(new_n703), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n700), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n707), .A2(new_n704), .A3(new_n700), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n705), .B1(new_n704), .B2(new_n700), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(G1981), .ZN(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  XOR2_X1   g290(.A(G1991), .B(G1996), .Z(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT92), .B(G1986), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n715), .A2(new_n717), .ZN(new_n720));
  AND3_X1   g295(.A1(new_n718), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n719), .B1(new_n718), .B2(new_n720), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n721), .A2(new_n722), .ZN(G229));
  INV_X1    g298(.A(G16), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G23), .ZN(new_n725));
  INV_X1    g300(.A(G288), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n725), .B1(new_n726), .B2(new_n724), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT94), .ZN(new_n728));
  XOR2_X1   g303(.A(KEYINPUT33), .B(G1976), .Z(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  OR2_X1    g305(.A1(G6), .A2(G16), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G305), .B2(new_n724), .ZN(new_n732));
  XOR2_X1   g307(.A(KEYINPUT32), .B(G1981), .Z(new_n733));
  NAND2_X1  g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  OR2_X1    g309(.A1(new_n732), .A2(new_n733), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n724), .A2(G22), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G166), .B2(new_n724), .ZN(new_n737));
  INV_X1    g312(.A(G1971), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  NAND4_X1  g314(.A1(new_n730), .A2(new_n734), .A3(new_n735), .A4(new_n739), .ZN(new_n740));
  OR2_X1    g315(.A1(new_n740), .A2(KEYINPUT34), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(KEYINPUT34), .ZN(new_n742));
  INV_X1    g317(.A(G290), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n743), .A2(G16), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G16), .B2(G24), .ZN(new_n745));
  INV_X1    g320(.A(G1986), .ZN(new_n746));
  AND2_X1   g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n745), .A2(new_n746), .ZN(new_n748));
  INV_X1    g323(.A(G29), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n749), .A2(G25), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n486), .A2(G131), .ZN(new_n751));
  OR2_X1    g326(.A1(G95), .A2(G2105), .ZN(new_n752));
  OAI211_X1 g327(.A(new_n752), .B(G2104), .C1(G107), .C2(new_n461), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT93), .Z(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(new_n478), .B2(G119), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n751), .A2(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(new_n756), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n750), .B1(new_n757), .B2(new_n749), .ZN(new_n758));
  XOR2_X1   g333(.A(KEYINPUT35), .B(G1991), .Z(new_n759));
  XOR2_X1   g334(.A(new_n758), .B(new_n759), .Z(new_n760));
  NOR3_X1   g335(.A1(new_n747), .A2(new_n748), .A3(new_n760), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n741), .A2(new_n742), .A3(new_n761), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT36), .Z(new_n763));
  NOR2_X1   g338(.A1(G4), .A2(G16), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT95), .Z(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(new_n633), .B2(new_n724), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(G1348), .Z(new_n767));
  NAND2_X1  g342(.A1(new_n724), .A2(G19), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(new_n552), .B2(new_n724), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(G1341), .Z(new_n770));
  NAND2_X1  g345(.A1(new_n724), .A2(G21), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G168), .B2(new_n724), .ZN(new_n772));
  INV_X1    g347(.A(G1966), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n749), .A2(G35), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT101), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G162), .B2(new_n749), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT29), .Z(new_n778));
  INV_X1    g353(.A(G2090), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  OAI211_X1 g355(.A(new_n770), .B(new_n774), .C1(new_n780), .C2(KEYINPUT102), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n749), .B1(KEYINPUT24), .B2(G34), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(KEYINPUT24), .B2(G34), .ZN(new_n783));
  INV_X1    g358(.A(G160), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n783), .B1(new_n784), .B2(G29), .ZN(new_n785));
  INV_X1    g360(.A(G2084), .ZN(new_n786));
  OR2_X1    g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n785), .A2(new_n786), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT31), .B(G11), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT100), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT30), .ZN(new_n791));
  AOI21_X1  g366(.A(G29), .B1(new_n791), .B2(G28), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(new_n791), .B2(G28), .ZN(new_n793));
  NAND4_X1  g368(.A1(new_n787), .A2(new_n788), .A3(new_n790), .A4(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(G164), .A2(new_n749), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(G27), .B2(new_n749), .ZN(new_n796));
  INV_X1    g371(.A(G2078), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n749), .A2(G33), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n800));
  INV_X1    g375(.A(KEYINPUT25), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  AOI22_X1  g377(.A1(new_n468), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n802), .B1(new_n803), .B2(new_n461), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(new_n486), .B2(G139), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n799), .B1(new_n805), .B2(new_n749), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n806), .A2(G2072), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n796), .A2(new_n797), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n806), .A2(G2072), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n798), .A2(new_n807), .A3(new_n808), .A4(new_n809), .ZN(new_n810));
  AOI211_X1 g385(.A(new_n794), .B(new_n810), .C1(G29), .C2(new_n659), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n724), .A2(G5), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(G171), .B2(new_n724), .ZN(new_n813));
  INV_X1    g388(.A(G1961), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n811), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n486), .A2(G141), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n463), .A2(G105), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT97), .ZN(new_n819));
  NAND3_X1  g394(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT26), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n821), .B1(new_n478), .B2(G129), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n817), .A2(new_n819), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n823), .A2(KEYINPUT98), .ZN(new_n824));
  INV_X1    g399(.A(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n823), .A2(KEYINPUT98), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n827), .A2(new_n749), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n828), .B1(new_n749), .B2(G32), .ZN(new_n829));
  XNOR2_X1  g404(.A(KEYINPUT27), .B(G1996), .ZN(new_n830));
  OAI22_X1  g405(.A1(new_n829), .A2(new_n830), .B1(new_n779), .B2(new_n778), .ZN(new_n831));
  NOR3_X1   g406(.A1(new_n781), .A2(new_n816), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n724), .A2(G20), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(KEYINPUT23), .Z(new_n834));
  AOI21_X1  g409(.A(new_n834), .B1(G299), .B2(G16), .ZN(new_n835));
  INV_X1    g410(.A(G1956), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n749), .A2(G26), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(KEYINPUT28), .Z(new_n839));
  NAND2_X1  g414(.A1(new_n486), .A2(G140), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n478), .A2(G128), .ZN(new_n841));
  OR2_X1    g416(.A1(G104), .A2(G2105), .ZN(new_n842));
  OAI211_X1 g417(.A(new_n842), .B(G2104), .C1(G116), .C2(new_n461), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n840), .A2(new_n841), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n839), .B1(new_n844), .B2(G29), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT96), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(G2067), .ZN(new_n847));
  AOI211_X1 g422(.A(new_n837), .B(new_n847), .C1(new_n780), .C2(KEYINPUT102), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n829), .A2(new_n830), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT99), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n832), .A2(new_n848), .A3(new_n850), .ZN(new_n851));
  NOR3_X1   g426(.A1(new_n763), .A2(new_n767), .A3(new_n851), .ZN(G311));
  INV_X1    g427(.A(G311), .ZN(G150));
  NAND2_X1  g428(.A1(G80), .A2(G543), .ZN(new_n854));
  INV_X1    g429(.A(G67), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n854), .B1(new_n509), .B2(new_n855), .ZN(new_n856));
  AOI22_X1  g431(.A1(new_n510), .A2(G93), .B1(G651), .B2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(G55), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n857), .B1(new_n858), .B2(new_n612), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(G860), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT104), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT37), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n633), .A2(new_n648), .ZN(new_n863));
  AND2_X1   g438(.A1(new_n859), .A2(new_n551), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n859), .A2(new_n551), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT38), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n863), .B(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT39), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(KEYINPUT103), .ZN(new_n871));
  INV_X1    g446(.A(G860), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n872), .B1(new_n868), .B2(new_n869), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n862), .B1(new_n871), .B2(new_n873), .ZN(G145));
  INV_X1    g449(.A(new_n805), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT105), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n492), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n490), .A2(KEYINPUT105), .A3(new_n491), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n498), .A2(KEYINPUT106), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT106), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n496), .A2(new_n881), .A3(new_n497), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n879), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(KEYINPUT107), .ZN(new_n885));
  AOI22_X1  g460(.A1(new_n877), .A2(new_n878), .B1(new_n880), .B2(new_n882), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT107), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(new_n844), .ZN(new_n890));
  INV_X1    g465(.A(new_n844), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n885), .A2(new_n891), .A3(new_n888), .ZN(new_n892));
  AND3_X1   g467(.A1(new_n890), .A2(new_n823), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n823), .B1(new_n890), .B2(new_n892), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n875), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT109), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  OAI211_X1 g472(.A(KEYINPUT109), .B(new_n875), .C1(new_n893), .C2(new_n894), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n890), .A2(new_n892), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT108), .ZN(new_n901));
  NOR3_X1   g476(.A1(new_n825), .A2(new_n826), .A3(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n826), .ZN(new_n903));
  AOI21_X1  g478(.A(KEYINPUT108), .B1(new_n903), .B2(new_n824), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n900), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n901), .B1(new_n825), .B2(new_n826), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n903), .A2(KEYINPUT108), .A3(new_n824), .ZN(new_n907));
  NAND4_X1  g482(.A1(new_n906), .A2(new_n907), .A3(new_n890), .A4(new_n892), .ZN(new_n908));
  AND3_X1   g483(.A1(new_n905), .A2(new_n805), .A3(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n899), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT110), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n756), .B(new_n664), .ZN(new_n913));
  OAI21_X1  g488(.A(G2104), .B1(new_n461), .B2(G118), .ZN(new_n914));
  INV_X1    g489(.A(G106), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n914), .B1(new_n915), .B2(new_n461), .ZN(new_n916));
  AND2_X1   g491(.A1(new_n478), .A2(G130), .ZN(new_n917));
  AOI211_X1 g492(.A(new_n916), .B(new_n917), .C1(G142), .C2(new_n486), .ZN(new_n918));
  XOR2_X1   g493(.A(new_n913), .B(new_n918), .Z(new_n919));
  NAND3_X1  g494(.A1(new_n911), .A2(new_n912), .A3(new_n919), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n659), .B(new_n784), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n921), .B(G162), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n909), .B1(new_n897), .B2(new_n898), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n919), .A2(new_n912), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n922), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(G37), .B1(new_n920), .B2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n919), .ZN(new_n927));
  AND2_X1   g502(.A1(new_n923), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n923), .A2(new_n927), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n922), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n926), .A2(new_n930), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n931), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g507(.A1(new_n859), .A2(new_n616), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n859), .B(new_n551), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n651), .B(new_n934), .ZN(new_n935));
  OAI21_X1  g510(.A(KEYINPUT111), .B1(new_n629), .B2(new_n644), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT111), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n612), .A2(KEYINPUT83), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n530), .A2(new_n626), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n938), .A2(new_n939), .A3(G54), .ZN(new_n940));
  NAND4_X1  g515(.A1(G299), .A2(new_n937), .A3(new_n940), .A4(new_n625), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n936), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n629), .A2(new_n644), .ZN(new_n943));
  AOI21_X1  g518(.A(KEYINPUT41), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n936), .A2(KEYINPUT112), .A3(new_n941), .ZN(new_n945));
  AOI21_X1  g520(.A(KEYINPUT112), .B1(new_n936), .B2(new_n941), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n943), .A2(KEYINPUT41), .ZN(new_n947));
  NOR3_X1   g522(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n935), .B1(new_n944), .B2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT112), .ZN(new_n950));
  NOR3_X1   g525(.A1(new_n629), .A2(new_n644), .A3(KEYINPUT111), .ZN(new_n951));
  INV_X1    g526(.A(G66), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n952), .B1(new_n559), .B2(new_n561), .ZN(new_n953));
  INV_X1    g528(.A(new_n619), .ZN(new_n954));
  OAI21_X1  g529(.A(G651), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  AND2_X1   g530(.A1(new_n622), .A2(new_n623), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n622), .A2(new_n623), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n955), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(G54), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n959), .B1(new_n612), .B2(KEYINPUT83), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n958), .B1(new_n960), .B2(new_n939), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n937), .B1(new_n961), .B2(G299), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n950), .B1(new_n951), .B2(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n936), .A2(KEYINPUT112), .A3(new_n941), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n963), .A2(new_n943), .A3(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n949), .B1(new_n966), .B2(new_n935), .ZN(new_n967));
  XNOR2_X1  g542(.A(G290), .B(G166), .ZN(new_n968));
  XNOR2_X1  g543(.A(G305), .B(G288), .ZN(new_n969));
  XNOR2_X1  g544(.A(new_n968), .B(new_n969), .ZN(new_n970));
  XOR2_X1   g545(.A(new_n970), .B(KEYINPUT42), .Z(new_n971));
  XNOR2_X1  g546(.A(new_n967), .B(new_n971), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n933), .B1(new_n972), .B2(new_n616), .ZN(G295));
  OAI21_X1  g548(.A(new_n933), .B1(new_n972), .B2(new_n616), .ZN(G331));
  INV_X1    g549(.A(KEYINPUT114), .ZN(new_n975));
  INV_X1    g550(.A(new_n580), .ZN(new_n976));
  AOI21_X1  g551(.A(G301), .B1(new_n976), .B2(new_n578), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n537), .A2(G301), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n866), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(G171), .B1(new_n579), .B2(new_n580), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n934), .A2(new_n981), .A3(new_n978), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n965), .A2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n947), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n963), .A2(new_n964), .A3(new_n985), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n943), .B1(new_n951), .B2(new_n962), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT41), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n983), .B1(new_n986), .B2(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n984), .B1(new_n990), .B2(KEYINPUT113), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT113), .ZN(new_n992));
  AOI211_X1 g567(.A(new_n992), .B(new_n983), .C1(new_n986), .C2(new_n989), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n975), .B1(new_n991), .B2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(new_n983), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n995), .B1(new_n948), .B2(new_n944), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(new_n992), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n990), .A2(KEYINPUT113), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n997), .A2(KEYINPUT114), .A3(new_n998), .A4(new_n984), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n994), .A2(new_n999), .A3(new_n970), .ZN(new_n1000));
  INV_X1    g575(.A(G37), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n991), .A2(new_n993), .ZN(new_n1002));
  INV_X1    g577(.A(new_n970), .ZN(new_n1003));
  AOI21_X1  g578(.A(KEYINPUT115), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT115), .ZN(new_n1005));
  NOR4_X1   g580(.A1(new_n991), .A2(new_n993), .A3(new_n970), .A4(new_n1005), .ZN(new_n1006));
  OAI211_X1 g581(.A(new_n1000), .B(new_n1001), .C1(new_n1004), .C2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(KEYINPUT43), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT44), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n997), .A2(new_n998), .A3(new_n984), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1005), .B1(new_n1010), .B2(new_n970), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1002), .A2(KEYINPUT115), .A3(new_n1003), .ZN(new_n1012));
  AOI21_X1  g587(.A(KEYINPUT43), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n995), .A2(KEYINPUT41), .A3(new_n987), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n970), .A2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n965), .B1(new_n995), .B2(KEYINPUT41), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1017), .A2(G37), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1013), .A2(new_n1018), .ZN(new_n1019));
  AND3_X1   g594(.A1(new_n1008), .A2(new_n1009), .A3(new_n1019), .ZN(new_n1020));
  AND2_X1   g595(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(new_n1013), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1018), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(KEYINPUT43), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1009), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(KEYINPUT116), .B1(new_n1020), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(KEYINPUT44), .ZN(new_n1028));
  AOI22_X1  g603(.A1(new_n1007), .A2(KEYINPUT43), .B1(new_n1013), .B2(new_n1018), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(new_n1009), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT116), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1028), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1026), .A2(new_n1032), .ZN(G397));
  INV_X1    g608(.A(G1384), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n885), .A2(new_n1034), .A3(new_n888), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT45), .ZN(new_n1036));
  AND2_X1   g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(G160), .A2(G40), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(G1996), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n827), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n823), .A2(G1996), .ZN(new_n1044));
  INV_X1    g619(.A(G2067), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n891), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n844), .A2(G2067), .ZN(new_n1047));
  AND2_X1   g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1043), .A2(new_n1044), .A3(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  XNOR2_X1  g625(.A(new_n756), .B(new_n759), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1050), .B(new_n1051), .C1(new_n746), .C2(new_n743), .ZN(new_n1052));
  NOR2_X1   g627(.A1(G290), .A2(G1986), .ZN(new_n1053));
  XNOR2_X1  g628(.A(new_n1053), .B(KEYINPUT117), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1041), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT118), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n884), .A2(new_n1056), .A3(new_n1034), .ZN(new_n1057));
  OAI21_X1  g632(.A(KEYINPUT118), .B1(new_n886), .B2(G1384), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT50), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NOR2_X1   g636(.A1(G164), .A2(G1384), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1038), .B1(new_n1063), .B2(KEYINPUT50), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1061), .A2(new_n786), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT120), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1064), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1068), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1069), .A2(KEYINPUT120), .A3(new_n786), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1038), .B1(new_n1062), .B2(KEYINPUT45), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1071), .B1(new_n1059), .B2(KEYINPUT45), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(new_n773), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1067), .A2(new_n1070), .A3(G168), .A4(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(G8), .ZN(new_n1075));
  AOI22_X1  g650(.A1(new_n1065), .A2(new_n1066), .B1(new_n1072), .B2(new_n773), .ZN(new_n1076));
  AOI21_X1  g651(.A(G168), .B1(new_n1076), .B2(new_n1070), .ZN(new_n1077));
  OAI21_X1  g652(.A(KEYINPUT51), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT62), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT51), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1074), .A2(new_n1080), .A3(G8), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1078), .A2(new_n1079), .A3(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT126), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n885), .A2(KEYINPUT45), .A3(new_n888), .A4(new_n1034), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1063), .A2(new_n1036), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1084), .A2(new_n1039), .A3(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(new_n738), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1057), .A2(new_n1058), .A3(KEYINPUT50), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1038), .B1(new_n1062), .B2(new_n1060), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1087), .B1(G2090), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(G8), .ZN(new_n1092));
  NAND2_X1  g667(.A1(G303), .A2(G8), .ZN(new_n1093));
  XNOR2_X1  g668(.A(new_n1093), .B(KEYINPUT55), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(G8), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1096), .B1(new_n1059), .B2(new_n1039), .ZN(new_n1097));
  INV_X1    g672(.A(G1976), .ZN(new_n1098));
  NOR2_X1   g673(.A1(G288), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(KEYINPUT52), .B1(G288), .B2(new_n1098), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1097), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  AOI211_X1 g677(.A(new_n1096), .B(new_n1099), .C1(new_n1059), .C2(new_n1039), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT52), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1102), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  OR2_X1    g680(.A1(G305), .A2(G1981), .ZN(new_n1106));
  NAND2_X1  g681(.A1(G305), .A2(G1981), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT49), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1106), .A2(KEYINPUT49), .A3(new_n1107), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1110), .A2(new_n1097), .A3(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(KEYINPUT119), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT119), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1110), .A2(new_n1114), .A3(new_n1097), .A4(new_n1111), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1105), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1069), .A2(new_n779), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1096), .B1(new_n1117), .B2(new_n1087), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1094), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1061), .A2(new_n1064), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1084), .A2(new_n797), .A3(new_n1039), .A4(new_n1085), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT53), .ZN(new_n1123));
  AOI22_X1  g698(.A1(new_n1121), .A2(new_n814), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n797), .A2(KEYINPUT53), .ZN(new_n1125));
  OR2_X1    g700(.A1(new_n1072), .A2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(G301), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1127));
  AND4_X1   g702(.A1(new_n1095), .A2(new_n1116), .A3(new_n1120), .A4(new_n1127), .ZN(new_n1128));
  AND3_X1   g703(.A1(new_n1082), .A2(new_n1083), .A3(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1083), .B1(new_n1082), .B2(new_n1128), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1079), .B1(new_n1078), .B2(new_n1081), .ZN(new_n1131));
  NOR3_X1   g706(.A1(new_n1129), .A2(new_n1130), .A3(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1133));
  XNOR2_X1  g708(.A(G301), .B(KEYINPUT54), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1037), .A2(new_n1125), .ZN(new_n1135));
  AND2_X1   g710(.A1(new_n1084), .A2(new_n1039), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1134), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  AOI22_X1  g712(.A1(new_n1133), .A2(new_n1134), .B1(new_n1137), .B2(new_n1124), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1138), .A2(new_n1095), .A3(new_n1116), .A4(new_n1120), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1139), .B1(new_n1078), .B2(new_n1081), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1059), .A2(new_n1045), .A3(new_n1039), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1141), .B1(new_n1069), .B2(G1348), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT60), .ZN(new_n1143));
  OR3_X1    g718(.A1(new_n1142), .A2(new_n1143), .A3(new_n633), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n633), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1144), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  XNOR2_X1  g722(.A(G299), .B(KEYINPUT123), .ZN(new_n1148));
  AOI21_X1  g723(.A(KEYINPUT122), .B1(new_n642), .B2(new_n643), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1149), .A2(KEYINPUT57), .ZN(new_n1150));
  XNOR2_X1  g725(.A(new_n1148), .B(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1151), .ZN(new_n1152));
  XNOR2_X1  g727(.A(KEYINPUT56), .B(G2072), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1153), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1086), .A2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(G1956), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1152), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1157), .A2(KEYINPUT125), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1136), .A2(new_n1085), .A3(new_n1153), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1156), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1159), .A2(new_n1151), .A3(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT125), .ZN(new_n1162));
  OAI211_X1 g737(.A(new_n1152), .B(new_n1162), .C1(new_n1155), .C2(new_n1156), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1158), .A2(KEYINPUT61), .A3(new_n1161), .A4(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1157), .A2(new_n1161), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT61), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1059), .A2(new_n1039), .ZN(new_n1168));
  XOR2_X1   g743(.A(KEYINPUT58), .B(G1341), .Z(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1084), .A2(new_n1042), .A3(new_n1039), .A4(new_n1085), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n551), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  XOR2_X1   g747(.A(new_n1172), .B(KEYINPUT59), .Z(new_n1173));
  NAND4_X1  g748(.A1(new_n1147), .A2(new_n1164), .A3(new_n1167), .A4(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1142), .A2(new_n634), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1175), .A2(KEYINPUT124), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT124), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1142), .A2(new_n1177), .A3(new_n634), .ZN(new_n1178));
  NAND4_X1  g753(.A1(new_n1176), .A2(new_n1158), .A3(new_n1163), .A4(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1179), .A2(new_n1161), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1174), .A2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1140), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1076), .A2(new_n1070), .ZN(new_n1183));
  NOR2_X1   g758(.A1(G286), .A2(new_n1096), .ZN(new_n1184));
  AND2_X1   g759(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NAND4_X1  g760(.A1(new_n1185), .A2(new_n1095), .A3(new_n1120), .A4(new_n1116), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT63), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT121), .ZN(new_n1189));
  AND2_X1   g764(.A1(new_n1116), .A2(new_n1120), .ZN(new_n1190));
  AOI22_X1  g765(.A1(new_n1069), .A2(new_n779), .B1(new_n1086), .B2(new_n738), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1094), .B1(new_n1191), .B2(new_n1096), .ZN(new_n1192));
  NAND4_X1  g767(.A1(new_n1192), .A2(new_n1183), .A3(KEYINPUT63), .A4(new_n1184), .ZN(new_n1193));
  INV_X1    g768(.A(new_n1193), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n1189), .B1(new_n1190), .B2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1116), .A2(new_n1120), .ZN(new_n1196));
  NOR3_X1   g771(.A1(new_n1196), .A2(new_n1193), .A3(KEYINPUT121), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1188), .B1(new_n1195), .B2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n1199), .A2(new_n1098), .A3(new_n726), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1200), .A2(new_n1106), .ZN(new_n1201));
  INV_X1    g776(.A(new_n1120), .ZN(new_n1202));
  AOI22_X1  g777(.A1(new_n1201), .A2(new_n1097), .B1(new_n1202), .B2(new_n1116), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1182), .A2(new_n1198), .A3(new_n1203), .ZN(new_n1204));
  OAI21_X1  g779(.A(new_n1055), .B1(new_n1132), .B2(new_n1204), .ZN(new_n1205));
  NOR2_X1   g780(.A1(new_n1040), .A2(G1996), .ZN(new_n1206));
  AND2_X1   g781(.A1(new_n1206), .A2(KEYINPUT46), .ZN(new_n1207));
  NOR2_X1   g782(.A1(new_n1206), .A2(KEYINPUT46), .ZN(new_n1208));
  INV_X1    g783(.A(new_n823), .ZN(new_n1209));
  AOI21_X1  g784(.A(new_n1040), .B1(new_n1209), .B2(new_n1048), .ZN(new_n1210));
  NOR3_X1   g785(.A1(new_n1207), .A2(new_n1208), .A3(new_n1210), .ZN(new_n1211));
  AND2_X1   g786(.A1(new_n1211), .A2(KEYINPUT47), .ZN(new_n1212));
  NOR2_X1   g787(.A1(new_n1211), .A2(KEYINPUT47), .ZN(new_n1213));
  AOI21_X1  g788(.A(new_n1040), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1214));
  AND3_X1   g789(.A1(new_n1041), .A2(KEYINPUT48), .A3(new_n1054), .ZN(new_n1215));
  AOI21_X1  g790(.A(KEYINPUT48), .B1(new_n1041), .B2(new_n1054), .ZN(new_n1216));
  NOR3_X1   g791(.A1(new_n1214), .A2(new_n1215), .A3(new_n1216), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n757), .A2(new_n759), .ZN(new_n1218));
  OAI21_X1  g793(.A(new_n1046), .B1(new_n1049), .B2(new_n1218), .ZN(new_n1219));
  AND2_X1   g794(.A1(new_n1219), .A2(new_n1041), .ZN(new_n1220));
  NOR4_X1   g795(.A1(new_n1212), .A2(new_n1213), .A3(new_n1217), .A4(new_n1220), .ZN(new_n1221));
  NAND2_X1  g796(.A1(new_n1205), .A2(new_n1221), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g797(.A1(G227), .A2(new_n459), .ZN(new_n1224));
  OAI211_X1 g798(.A(new_n685), .B(new_n1224), .C1(new_n721), .C2(new_n722), .ZN(new_n1225));
  INV_X1    g799(.A(new_n1225), .ZN(new_n1226));
  NAND2_X1  g800(.A1(new_n923), .A2(new_n924), .ZN(new_n1227));
  INV_X1    g801(.A(new_n922), .ZN(new_n1228));
  NAND2_X1  g802(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  NOR3_X1   g803(.A1(new_n923), .A2(KEYINPUT110), .A3(new_n927), .ZN(new_n1230));
  OAI21_X1  g804(.A(new_n1001), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g805(.A1(new_n911), .A2(new_n919), .ZN(new_n1232));
  NAND2_X1  g806(.A1(new_n923), .A2(new_n927), .ZN(new_n1233));
  AOI21_X1  g807(.A(new_n1228), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  OAI21_X1  g808(.A(new_n1226), .B1(new_n1231), .B2(new_n1234), .ZN(new_n1235));
  OAI21_X1  g809(.A(KEYINPUT127), .B1(new_n1235), .B2(new_n1029), .ZN(new_n1236));
  AOI21_X1  g810(.A(new_n1225), .B1(new_n926), .B2(new_n930), .ZN(new_n1237));
  INV_X1    g811(.A(KEYINPUT127), .ZN(new_n1238));
  INV_X1    g812(.A(new_n1019), .ZN(new_n1239));
  AND2_X1   g813(.A1(new_n1007), .A2(KEYINPUT43), .ZN(new_n1240));
  OAI211_X1 g814(.A(new_n1237), .B(new_n1238), .C1(new_n1239), .C2(new_n1240), .ZN(new_n1241));
  AND2_X1   g815(.A1(new_n1236), .A2(new_n1241), .ZN(G308));
  OAI21_X1  g816(.A(new_n1237), .B1(new_n1240), .B2(new_n1239), .ZN(G225));
endmodule


