

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U564 ( .A1(n622), .A2(n621), .ZN(n1016) );
  XNOR2_X2 U565 ( .A(n688), .B(KEYINPUT32), .ZN(n697) );
  NAND2_X4 U566 ( .A1(n608), .A2(n708), .ZN(n680) );
  NOR2_X2 U567 ( .A1(n617), .A2(n616), .ZN(n619) );
  XOR2_X1 U568 ( .A(KEYINPUT1), .B(n542), .Z(n799) );
  NOR2_X2 U569 ( .A1(n643), .A2(n1009), .ZN(n636) );
  NOR2_X1 U570 ( .A1(G2104), .A2(G2105), .ZN(n535) );
  XNOR2_X1 U571 ( .A(n619), .B(n618), .ZN(n622) );
  NOR2_X2 U572 ( .A1(G2104), .A2(n536), .ZN(n553) );
  NOR2_X1 U573 ( .A1(n1016), .A2(n624), .ZN(n626) );
  INV_X1 U574 ( .A(KEYINPUT29), .ZN(n659) );
  NOR2_X1 U575 ( .A1(n749), .A2(n702), .ZN(n703) );
  INV_X1 U576 ( .A(KEYINPUT13), .ZN(n614) );
  NOR2_X1 U577 ( .A1(n1018), .A2(n704), .ZN(n738) );
  XNOR2_X1 U578 ( .A(n615), .B(n614), .ZN(n616) );
  INV_X1 U579 ( .A(KEYINPUT71), .ZN(n618) );
  NOR2_X1 U580 ( .A1(n591), .A2(n545), .ZN(n803) );
  NOR2_X2 U581 ( .A1(n530), .A2(G2105), .ZN(n891) );
  NOR2_X1 U582 ( .A1(G651), .A2(n591), .ZN(n798) );
  BUF_X1 U583 ( .A(n606), .Z(G160) );
  INV_X1 U584 ( .A(G2104), .ZN(n530) );
  NAND2_X1 U585 ( .A1(G101), .A2(n891), .ZN(n531) );
  XOR2_X1 U586 ( .A(n531), .B(KEYINPUT23), .Z(n534) );
  INV_X1 U587 ( .A(G2105), .ZN(n536) );
  NAND2_X1 U588 ( .A1(G125), .A2(n553), .ZN(n532) );
  XNOR2_X1 U589 ( .A(n532), .B(KEYINPUT64), .ZN(n533) );
  NAND2_X1 U590 ( .A1(n534), .A2(n533), .ZN(n540) );
  XOR2_X2 U591 ( .A(KEYINPUT17), .B(n535), .Z(n892) );
  NAND2_X1 U592 ( .A1(n892), .A2(G137), .ZN(n538) );
  AND2_X1 U593 ( .A1(G2104), .A2(G2105), .ZN(n895) );
  NAND2_X1 U594 ( .A1(n895), .A2(G113), .ZN(n537) );
  NAND2_X1 U595 ( .A1(n538), .A2(n537), .ZN(n539) );
  NOR2_X1 U596 ( .A1(n540), .A2(n539), .ZN(n606) );
  XOR2_X1 U597 ( .A(G543), .B(KEYINPUT0), .Z(n591) );
  NAND2_X1 U598 ( .A1(G48), .A2(n798), .ZN(n541) );
  XNOR2_X1 U599 ( .A(n541), .B(KEYINPUT84), .ZN(n550) );
  NOR2_X1 U600 ( .A1(G543), .A2(G651), .ZN(n802) );
  NAND2_X1 U601 ( .A1(G86), .A2(n802), .ZN(n544) );
  INV_X1 U602 ( .A(G651), .ZN(n545) );
  NOR2_X1 U603 ( .A1(G543), .A2(n545), .ZN(n542) );
  NAND2_X1 U604 ( .A1(G61), .A2(n799), .ZN(n543) );
  NAND2_X1 U605 ( .A1(n544), .A2(n543), .ZN(n548) );
  NAND2_X1 U606 ( .A1(n803), .A2(G73), .ZN(n546) );
  XOR2_X1 U607 ( .A(KEYINPUT2), .B(n546), .Z(n547) );
  NOR2_X1 U608 ( .A1(n548), .A2(n547), .ZN(n549) );
  NAND2_X1 U609 ( .A1(n550), .A2(n549), .ZN(G305) );
  NAND2_X1 U610 ( .A1(G102), .A2(n891), .ZN(n552) );
  NAND2_X1 U611 ( .A1(G138), .A2(n892), .ZN(n551) );
  NAND2_X1 U612 ( .A1(n552), .A2(n551), .ZN(n557) );
  NAND2_X1 U613 ( .A1(G126), .A2(n553), .ZN(n555) );
  NAND2_X1 U614 ( .A1(G114), .A2(n895), .ZN(n554) );
  NAND2_X1 U615 ( .A1(n555), .A2(n554), .ZN(n556) );
  NOR2_X1 U616 ( .A1(n557), .A2(n556), .ZN(G164) );
  NAND2_X1 U617 ( .A1(G53), .A2(n798), .ZN(n559) );
  NAND2_X1 U618 ( .A1(G65), .A2(n799), .ZN(n558) );
  NAND2_X1 U619 ( .A1(n559), .A2(n558), .ZN(n563) );
  NAND2_X1 U620 ( .A1(G91), .A2(n802), .ZN(n561) );
  NAND2_X1 U621 ( .A1(G78), .A2(n803), .ZN(n560) );
  NAND2_X1 U622 ( .A1(n561), .A2(n560), .ZN(n562) );
  NOR2_X1 U623 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U624 ( .A(KEYINPUT68), .B(n564), .Z(G299) );
  NAND2_X1 U625 ( .A1(G90), .A2(n802), .ZN(n566) );
  NAND2_X1 U626 ( .A1(G77), .A2(n803), .ZN(n565) );
  NAND2_X1 U627 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U628 ( .A(n567), .B(KEYINPUT9), .ZN(n569) );
  NAND2_X1 U629 ( .A1(G52), .A2(n798), .ZN(n568) );
  NAND2_X1 U630 ( .A1(n569), .A2(n568), .ZN(n572) );
  NAND2_X1 U631 ( .A1(G64), .A2(n799), .ZN(n570) );
  XNOR2_X1 U632 ( .A(KEYINPUT67), .B(n570), .ZN(n571) );
  NOR2_X1 U633 ( .A1(n572), .A2(n571), .ZN(G171) );
  NAND2_X1 U634 ( .A1(n802), .A2(G89), .ZN(n573) );
  XNOR2_X1 U635 ( .A(n573), .B(KEYINPUT4), .ZN(n575) );
  NAND2_X1 U636 ( .A1(G76), .A2(n803), .ZN(n574) );
  NAND2_X1 U637 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U638 ( .A(KEYINPUT5), .B(n576), .ZN(n583) );
  XNOR2_X1 U639 ( .A(KEYINPUT77), .B(KEYINPUT78), .ZN(n581) );
  NAND2_X1 U640 ( .A1(G51), .A2(n798), .ZN(n578) );
  NAND2_X1 U641 ( .A1(G63), .A2(n799), .ZN(n577) );
  NAND2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U643 ( .A(n579), .B(KEYINPUT6), .ZN(n580) );
  XNOR2_X1 U644 ( .A(n581), .B(n580), .ZN(n582) );
  NAND2_X1 U645 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U646 ( .A(KEYINPUT7), .B(n584), .ZN(G168) );
  XOR2_X1 U647 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U648 ( .A1(G88), .A2(n802), .ZN(n586) );
  NAND2_X1 U649 ( .A1(G75), .A2(n803), .ZN(n585) );
  NAND2_X1 U650 ( .A1(n586), .A2(n585), .ZN(n590) );
  NAND2_X1 U651 ( .A1(G50), .A2(n798), .ZN(n588) );
  NAND2_X1 U652 ( .A1(G62), .A2(n799), .ZN(n587) );
  NAND2_X1 U653 ( .A1(n588), .A2(n587), .ZN(n589) );
  NOR2_X1 U654 ( .A1(n590), .A2(n589), .ZN(G166) );
  INV_X1 U655 ( .A(G166), .ZN(G303) );
  NAND2_X1 U656 ( .A1(G49), .A2(n798), .ZN(n593) );
  NAND2_X1 U657 ( .A1(G87), .A2(n591), .ZN(n592) );
  NAND2_X1 U658 ( .A1(n593), .A2(n592), .ZN(n594) );
  NOR2_X1 U659 ( .A1(n799), .A2(n594), .ZN(n597) );
  NAND2_X1 U660 ( .A1(G74), .A2(G651), .ZN(n595) );
  XOR2_X1 U661 ( .A(KEYINPUT83), .B(n595), .Z(n596) );
  NAND2_X1 U662 ( .A1(n597), .A2(n596), .ZN(G288) );
  NAND2_X1 U663 ( .A1(G60), .A2(n799), .ZN(n598) );
  XNOR2_X1 U664 ( .A(n598), .B(KEYINPUT66), .ZN(n600) );
  NAND2_X1 U665 ( .A1(n803), .A2(G72), .ZN(n599) );
  NAND2_X1 U666 ( .A1(n600), .A2(n599), .ZN(n603) );
  NAND2_X1 U667 ( .A1(G85), .A2(n802), .ZN(n601) );
  XNOR2_X1 U668 ( .A(KEYINPUT65), .B(n601), .ZN(n602) );
  NOR2_X1 U669 ( .A1(n603), .A2(n602), .ZN(n605) );
  NAND2_X1 U670 ( .A1(n798), .A2(G47), .ZN(n604) );
  NAND2_X1 U671 ( .A1(n605), .A2(n604), .ZN(G290) );
  XNOR2_X1 U672 ( .A(G1981), .B(G305), .ZN(n1018) );
  NAND2_X1 U673 ( .A1(G40), .A2(n606), .ZN(n607) );
  XNOR2_X1 U674 ( .A(n607), .B(KEYINPUT88), .ZN(n707) );
  INV_X1 U675 ( .A(n707), .ZN(n608) );
  NOR2_X1 U676 ( .A1(G164), .A2(G1384), .ZN(n708) );
  NAND2_X1 U677 ( .A1(G8), .A2(n680), .ZN(n749) );
  XOR2_X1 U678 ( .A(KEYINPUT70), .B(KEYINPUT14), .Z(n610) );
  NAND2_X1 U679 ( .A1(G56), .A2(n799), .ZN(n609) );
  XNOR2_X1 U680 ( .A(n610), .B(n609), .ZN(n617) );
  NAND2_X1 U681 ( .A1(G68), .A2(n803), .ZN(n613) );
  NAND2_X1 U682 ( .A1(n802), .A2(G81), .ZN(n611) );
  XNOR2_X1 U683 ( .A(n611), .B(KEYINPUT12), .ZN(n612) );
  NAND2_X1 U684 ( .A1(n613), .A2(n612), .ZN(n615) );
  NAND2_X1 U685 ( .A1(n798), .A2(G43), .ZN(n620) );
  XNOR2_X1 U686 ( .A(KEYINPUT72), .B(n620), .ZN(n621) );
  INV_X1 U687 ( .A(G1996), .ZN(n983) );
  NOR2_X1 U688 ( .A1(n680), .A2(n983), .ZN(n623) );
  XNOR2_X1 U689 ( .A(n623), .B(KEYINPUT26), .ZN(n624) );
  NAND2_X1 U690 ( .A1(G1341), .A2(n680), .ZN(n625) );
  NAND2_X1 U691 ( .A1(n626), .A2(n625), .ZN(n643) );
  NAND2_X1 U692 ( .A1(n803), .A2(G79), .ZN(n633) );
  NAND2_X1 U693 ( .A1(G54), .A2(n798), .ZN(n628) );
  NAND2_X1 U694 ( .A1(G66), .A2(n799), .ZN(n627) );
  NAND2_X1 U695 ( .A1(n628), .A2(n627), .ZN(n631) );
  NAND2_X1 U696 ( .A1(G92), .A2(n802), .ZN(n629) );
  XNOR2_X1 U697 ( .A(KEYINPUT75), .B(n629), .ZN(n630) );
  NOR2_X1 U698 ( .A1(n631), .A2(n630), .ZN(n632) );
  NAND2_X1 U699 ( .A1(n633), .A2(n632), .ZN(n634) );
  XOR2_X1 U700 ( .A(KEYINPUT15), .B(n634), .Z(n1009) );
  INV_X1 U701 ( .A(KEYINPUT100), .ZN(n635) );
  XNOR2_X1 U702 ( .A(n636), .B(n635), .ZN(n642) );
  INV_X1 U703 ( .A(G2067), .ZN(n637) );
  NOR2_X1 U704 ( .A1(n680), .A2(n637), .ZN(n638) );
  XNOR2_X1 U705 ( .A(n638), .B(KEYINPUT101), .ZN(n640) );
  NAND2_X1 U706 ( .A1(n680), .A2(G1348), .ZN(n639) );
  NAND2_X1 U707 ( .A1(n640), .A2(n639), .ZN(n641) );
  NAND2_X1 U708 ( .A1(n642), .A2(n641), .ZN(n645) );
  NAND2_X1 U709 ( .A1(n643), .A2(n1009), .ZN(n644) );
  NAND2_X1 U710 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U711 ( .A(KEYINPUT102), .B(n646), .ZN(n653) );
  INV_X1 U712 ( .A(G2072), .ZN(n971) );
  NOR2_X1 U713 ( .A1(n680), .A2(n971), .ZN(n648) );
  XNOR2_X1 U714 ( .A(KEYINPUT27), .B(KEYINPUT98), .ZN(n647) );
  XNOR2_X1 U715 ( .A(n648), .B(n647), .ZN(n650) );
  NAND2_X1 U716 ( .A1(n680), .A2(G1956), .ZN(n649) );
  NAND2_X1 U717 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U718 ( .A(KEYINPUT99), .B(n651), .ZN(n655) );
  INV_X1 U719 ( .A(G299), .ZN(n654) );
  NAND2_X1 U720 ( .A1(n655), .A2(n654), .ZN(n652) );
  NAND2_X1 U721 ( .A1(n653), .A2(n652), .ZN(n658) );
  NOR2_X1 U722 ( .A1(n655), .A2(n654), .ZN(n656) );
  XOR2_X1 U723 ( .A(n656), .B(KEYINPUT28), .Z(n657) );
  NAND2_X1 U724 ( .A1(n658), .A2(n657), .ZN(n660) );
  XNOR2_X1 U725 ( .A(n660), .B(n659), .ZN(n667) );
  XOR2_X1 U726 ( .A(G2078), .B(KEYINPUT25), .Z(n984) );
  NOR2_X1 U727 ( .A1(n984), .A2(n680), .ZN(n661) );
  XOR2_X1 U728 ( .A(KEYINPUT96), .B(n661), .Z(n664) );
  XOR2_X1 U729 ( .A(KEYINPUT94), .B(G1961), .Z(n929) );
  NAND2_X1 U730 ( .A1(n929), .A2(n680), .ZN(n662) );
  XOR2_X1 U731 ( .A(KEYINPUT95), .B(n662), .Z(n663) );
  NAND2_X1 U732 ( .A1(n664), .A2(n663), .ZN(n672) );
  NAND2_X1 U733 ( .A1(G171), .A2(n672), .ZN(n665) );
  XOR2_X1 U734 ( .A(KEYINPUT97), .B(n665), .Z(n666) );
  NAND2_X1 U735 ( .A1(n667), .A2(n666), .ZN(n677) );
  NOR2_X1 U736 ( .A1(G1966), .A2(n749), .ZN(n691) );
  NOR2_X1 U737 ( .A1(G2084), .A2(n680), .ZN(n692) );
  NOR2_X1 U738 ( .A1(n691), .A2(n692), .ZN(n668) );
  NAND2_X1 U739 ( .A1(G8), .A2(n668), .ZN(n669) );
  XNOR2_X1 U740 ( .A(KEYINPUT30), .B(n669), .ZN(n670) );
  XOR2_X1 U741 ( .A(KEYINPUT103), .B(n670), .Z(n671) );
  NOR2_X1 U742 ( .A1(G168), .A2(n671), .ZN(n674) );
  NOR2_X1 U743 ( .A1(G171), .A2(n672), .ZN(n673) );
  NOR2_X1 U744 ( .A1(n674), .A2(n673), .ZN(n675) );
  XOR2_X1 U745 ( .A(KEYINPUT31), .B(n675), .Z(n676) );
  NAND2_X1 U746 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U747 ( .A(n678), .B(KEYINPUT104), .ZN(n689) );
  AND2_X1 U748 ( .A1(G286), .A2(G8), .ZN(n679) );
  NAND2_X1 U749 ( .A1(n689), .A2(n679), .ZN(n687) );
  INV_X1 U750 ( .A(G8), .ZN(n685) );
  NOR2_X1 U751 ( .A1(G1971), .A2(n749), .ZN(n682) );
  NOR2_X1 U752 ( .A1(G2090), .A2(n680), .ZN(n681) );
  NOR2_X1 U753 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U754 ( .A1(n683), .A2(G303), .ZN(n684) );
  OR2_X1 U755 ( .A1(n685), .A2(n684), .ZN(n686) );
  AND2_X1 U756 ( .A1(n687), .A2(n686), .ZN(n688) );
  INV_X1 U757 ( .A(n689), .ZN(n690) );
  NOR2_X1 U758 ( .A1(n691), .A2(n690), .ZN(n695) );
  NAND2_X1 U759 ( .A1(G8), .A2(n692), .ZN(n693) );
  XOR2_X1 U760 ( .A(KEYINPUT93), .B(n693), .Z(n694) );
  NAND2_X1 U761 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U762 ( .A1(n697), .A2(n696), .ZN(n741) );
  NOR2_X1 U763 ( .A1(G1976), .A2(G288), .ZN(n698) );
  XOR2_X1 U764 ( .A(KEYINPUT105), .B(n698), .Z(n1005) );
  NOR2_X1 U765 ( .A1(G1971), .A2(G303), .ZN(n699) );
  NOR2_X1 U766 ( .A1(n1005), .A2(n699), .ZN(n700) );
  NAND2_X1 U767 ( .A1(n741), .A2(n700), .ZN(n701) );
  NAND2_X1 U768 ( .A1(G1976), .A2(G288), .ZN(n1006) );
  NAND2_X1 U769 ( .A1(n701), .A2(n1006), .ZN(n702) );
  NOR2_X1 U770 ( .A1(KEYINPUT33), .A2(n703), .ZN(n704) );
  INV_X1 U771 ( .A(n1005), .ZN(n705) );
  NOR2_X1 U772 ( .A1(n749), .A2(n705), .ZN(n706) );
  NAND2_X1 U773 ( .A1(KEYINPUT33), .A2(n706), .ZN(n736) );
  NOR2_X1 U774 ( .A1(n707), .A2(n708), .ZN(n768) );
  XNOR2_X1 U775 ( .A(KEYINPUT37), .B(G2067), .ZN(n758) );
  NAND2_X1 U776 ( .A1(G104), .A2(n891), .ZN(n710) );
  NAND2_X1 U777 ( .A1(G140), .A2(n892), .ZN(n709) );
  NAND2_X1 U778 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U779 ( .A(KEYINPUT34), .B(n711), .ZN(n716) );
  NAND2_X1 U780 ( .A1(G128), .A2(n553), .ZN(n713) );
  NAND2_X1 U781 ( .A1(G116), .A2(n895), .ZN(n712) );
  NAND2_X1 U782 ( .A1(n713), .A2(n712), .ZN(n714) );
  XOR2_X1 U783 ( .A(KEYINPUT35), .B(n714), .Z(n715) );
  NOR2_X1 U784 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U785 ( .A(KEYINPUT36), .B(n717), .ZN(n888) );
  NOR2_X1 U786 ( .A1(n758), .A2(n888), .ZN(n963) );
  NAND2_X1 U787 ( .A1(n768), .A2(n963), .ZN(n765) );
  NAND2_X1 U788 ( .A1(G131), .A2(n892), .ZN(n724) );
  NAND2_X1 U789 ( .A1(G119), .A2(n553), .ZN(n719) );
  NAND2_X1 U790 ( .A1(G107), .A2(n895), .ZN(n718) );
  NAND2_X1 U791 ( .A1(n719), .A2(n718), .ZN(n722) );
  NAND2_X1 U792 ( .A1(G95), .A2(n891), .ZN(n720) );
  XNOR2_X1 U793 ( .A(KEYINPUT89), .B(n720), .ZN(n721) );
  NOR2_X1 U794 ( .A1(n722), .A2(n721), .ZN(n723) );
  NAND2_X1 U795 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U796 ( .A(n725), .B(KEYINPUT90), .ZN(n871) );
  NAND2_X1 U797 ( .A1(n871), .A2(G1991), .ZN(n734) );
  NAND2_X1 U798 ( .A1(G117), .A2(n895), .ZN(n727) );
  NAND2_X1 U799 ( .A1(G141), .A2(n892), .ZN(n726) );
  NAND2_X1 U800 ( .A1(n727), .A2(n726), .ZN(n730) );
  NAND2_X1 U801 ( .A1(n891), .A2(G105), .ZN(n728) );
  XOR2_X1 U802 ( .A(KEYINPUT38), .B(n728), .Z(n729) );
  NOR2_X1 U803 ( .A1(n730), .A2(n729), .ZN(n732) );
  NAND2_X1 U804 ( .A1(n553), .A2(G129), .ZN(n731) );
  NAND2_X1 U805 ( .A1(n732), .A2(n731), .ZN(n887) );
  NAND2_X1 U806 ( .A1(G1996), .A2(n887), .ZN(n733) );
  NAND2_X1 U807 ( .A1(n734), .A2(n733), .ZN(n964) );
  NAND2_X1 U808 ( .A1(n768), .A2(n964), .ZN(n761) );
  XOR2_X1 U809 ( .A(KEYINPUT91), .B(n761), .Z(n735) );
  AND2_X1 U810 ( .A1(n765), .A2(n735), .ZN(n745) );
  AND2_X1 U811 ( .A1(n736), .A2(n745), .ZN(n737) );
  NAND2_X1 U812 ( .A1(n738), .A2(n737), .ZN(n755) );
  NOR2_X1 U813 ( .A1(G2090), .A2(G303), .ZN(n739) );
  NAND2_X1 U814 ( .A1(G8), .A2(n739), .ZN(n740) );
  NAND2_X1 U815 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U816 ( .A(n742), .B(KEYINPUT106), .ZN(n744) );
  AND2_X1 U817 ( .A1(n749), .A2(n745), .ZN(n743) );
  NAND2_X1 U818 ( .A1(n744), .A2(n743), .ZN(n753) );
  INV_X1 U819 ( .A(n745), .ZN(n751) );
  NOR2_X1 U820 ( .A1(G1981), .A2(G305), .ZN(n746) );
  XOR2_X1 U821 ( .A(n746), .B(KEYINPUT92), .Z(n747) );
  XNOR2_X1 U822 ( .A(KEYINPUT24), .B(n747), .ZN(n748) );
  OR2_X1 U823 ( .A1(n749), .A2(n748), .ZN(n750) );
  OR2_X1 U824 ( .A1(n751), .A2(n750), .ZN(n752) );
  AND2_X1 U825 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U826 ( .A1(n755), .A2(n754), .ZN(n757) );
  XNOR2_X1 U827 ( .A(G1986), .B(G290), .ZN(n1015) );
  NAND2_X1 U828 ( .A1(n1015), .A2(n768), .ZN(n756) );
  NAND2_X1 U829 ( .A1(n757), .A2(n756), .ZN(n771) );
  NAND2_X1 U830 ( .A1(n758), .A2(n888), .ZN(n975) );
  NOR2_X1 U831 ( .A1(G1991), .A2(n871), .ZN(n962) );
  NOR2_X1 U832 ( .A1(G1986), .A2(G290), .ZN(n759) );
  NOR2_X1 U833 ( .A1(n962), .A2(n759), .ZN(n760) );
  XNOR2_X1 U834 ( .A(n760), .B(KEYINPUT107), .ZN(n762) );
  NAND2_X1 U835 ( .A1(n762), .A2(n761), .ZN(n763) );
  OR2_X1 U836 ( .A1(n887), .A2(G1996), .ZN(n957) );
  NAND2_X1 U837 ( .A1(n763), .A2(n957), .ZN(n764) );
  XOR2_X1 U838 ( .A(KEYINPUT39), .B(n764), .Z(n766) );
  NAND2_X1 U839 ( .A1(n766), .A2(n765), .ZN(n767) );
  NAND2_X1 U840 ( .A1(n975), .A2(n767), .ZN(n769) );
  NAND2_X1 U841 ( .A1(n769), .A2(n768), .ZN(n770) );
  NAND2_X1 U842 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U843 ( .A(n772), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U844 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U845 ( .A1(G111), .A2(n895), .ZN(n774) );
  NAND2_X1 U846 ( .A1(G135), .A2(n892), .ZN(n773) );
  NAND2_X1 U847 ( .A1(n774), .A2(n773), .ZN(n778) );
  NAND2_X1 U848 ( .A1(G123), .A2(n553), .ZN(n775) );
  XNOR2_X1 U849 ( .A(n775), .B(KEYINPUT81), .ZN(n776) );
  XNOR2_X1 U850 ( .A(n776), .B(KEYINPUT18), .ZN(n777) );
  NOR2_X1 U851 ( .A1(n778), .A2(n777), .ZN(n780) );
  NAND2_X1 U852 ( .A1(n891), .A2(G99), .ZN(n779) );
  NAND2_X1 U853 ( .A1(n780), .A2(n779), .ZN(n959) );
  XNOR2_X1 U854 ( .A(G2096), .B(n959), .ZN(n781) );
  OR2_X1 U855 ( .A1(G2100), .A2(n781), .ZN(G156) );
  INV_X1 U856 ( .A(G57), .ZN(G237) );
  INV_X1 U857 ( .A(G120), .ZN(G236) );
  NAND2_X1 U858 ( .A1(G7), .A2(G661), .ZN(n782) );
  XNOR2_X1 U859 ( .A(n782), .B(KEYINPUT10), .ZN(G223) );
  XNOR2_X1 U860 ( .A(G223), .B(KEYINPUT69), .ZN(n834) );
  NAND2_X1 U861 ( .A1(n834), .A2(G567), .ZN(n783) );
  XOR2_X1 U862 ( .A(KEYINPUT11), .B(n783), .Z(G234) );
  INV_X1 U863 ( .A(G860), .ZN(n790) );
  OR2_X1 U864 ( .A1(n1016), .A2(n790), .ZN(n784) );
  XOR2_X1 U865 ( .A(KEYINPUT73), .B(n784), .Z(G153) );
  XOR2_X1 U866 ( .A(G171), .B(KEYINPUT74), .Z(G301) );
  INV_X1 U867 ( .A(G868), .ZN(n817) );
  NOR2_X1 U868 ( .A1(G301), .A2(n817), .ZN(n786) );
  NOR2_X1 U869 ( .A1(G868), .A2(n1009), .ZN(n785) );
  NOR2_X1 U870 ( .A1(n786), .A2(n785), .ZN(n787) );
  XNOR2_X1 U871 ( .A(KEYINPUT76), .B(n787), .ZN(G284) );
  NOR2_X1 U872 ( .A1(G286), .A2(n817), .ZN(n789) );
  NOR2_X1 U873 ( .A1(G299), .A2(G868), .ZN(n788) );
  NOR2_X1 U874 ( .A1(n789), .A2(n788), .ZN(G297) );
  NAND2_X1 U875 ( .A1(n790), .A2(G559), .ZN(n791) );
  INV_X1 U876 ( .A(n1009), .ZN(n908) );
  NAND2_X1 U877 ( .A1(n791), .A2(n908), .ZN(n792) );
  XNOR2_X1 U878 ( .A(n792), .B(KEYINPUT16), .ZN(n793) );
  XOR2_X1 U879 ( .A(KEYINPUT79), .B(n793), .Z(G148) );
  NOR2_X1 U880 ( .A1(n1009), .A2(n817), .ZN(n794) );
  XOR2_X1 U881 ( .A(KEYINPUT80), .B(n794), .Z(n795) );
  NOR2_X1 U882 ( .A1(G559), .A2(n795), .ZN(n797) );
  NOR2_X1 U883 ( .A1(G868), .A2(n1016), .ZN(n796) );
  NOR2_X1 U884 ( .A1(n797), .A2(n796), .ZN(G282) );
  NAND2_X1 U885 ( .A1(n908), .A2(G559), .ZN(n838) );
  XNOR2_X1 U886 ( .A(G290), .B(G288), .ZN(n814) );
  XOR2_X1 U887 ( .A(KEYINPUT85), .B(KEYINPUT19), .Z(n810) );
  NAND2_X1 U888 ( .A1(G55), .A2(n798), .ZN(n801) );
  NAND2_X1 U889 ( .A1(G67), .A2(n799), .ZN(n800) );
  NAND2_X1 U890 ( .A1(n801), .A2(n800), .ZN(n807) );
  NAND2_X1 U891 ( .A1(G93), .A2(n802), .ZN(n805) );
  NAND2_X1 U892 ( .A1(G80), .A2(n803), .ZN(n804) );
  NAND2_X1 U893 ( .A1(n805), .A2(n804), .ZN(n806) );
  NOR2_X1 U894 ( .A1(n807), .A2(n806), .ZN(n808) );
  XOR2_X1 U895 ( .A(KEYINPUT82), .B(n808), .Z(n841) );
  XNOR2_X1 U896 ( .A(G166), .B(n841), .ZN(n809) );
  XNOR2_X1 U897 ( .A(n810), .B(n809), .ZN(n811) );
  XNOR2_X1 U898 ( .A(G299), .B(n811), .ZN(n812) );
  XNOR2_X1 U899 ( .A(n812), .B(G305), .ZN(n813) );
  XNOR2_X1 U900 ( .A(n814), .B(n813), .ZN(n815) );
  XNOR2_X1 U901 ( .A(n1016), .B(n815), .ZN(n907) );
  XNOR2_X1 U902 ( .A(n838), .B(n907), .ZN(n816) );
  NAND2_X1 U903 ( .A1(n816), .A2(G868), .ZN(n819) );
  NAND2_X1 U904 ( .A1(n841), .A2(n817), .ZN(n818) );
  NAND2_X1 U905 ( .A1(n819), .A2(n818), .ZN(G295) );
  NAND2_X1 U906 ( .A1(G2078), .A2(G2084), .ZN(n820) );
  XOR2_X1 U907 ( .A(KEYINPUT20), .B(n820), .Z(n821) );
  NAND2_X1 U908 ( .A1(G2090), .A2(n821), .ZN(n822) );
  XNOR2_X1 U909 ( .A(KEYINPUT21), .B(n822), .ZN(n823) );
  NAND2_X1 U910 ( .A1(n823), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U911 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U912 ( .A1(G236), .A2(G237), .ZN(n824) );
  NAND2_X1 U913 ( .A1(G69), .A2(n824), .ZN(n825) );
  XNOR2_X1 U914 ( .A(KEYINPUT87), .B(n825), .ZN(n826) );
  NAND2_X1 U915 ( .A1(n826), .A2(G108), .ZN(n842) );
  NAND2_X1 U916 ( .A1(n842), .A2(G567), .ZN(n832) );
  NAND2_X1 U917 ( .A1(G132), .A2(G82), .ZN(n827) );
  XNOR2_X1 U918 ( .A(n827), .B(KEYINPUT86), .ZN(n828) );
  XNOR2_X1 U919 ( .A(n828), .B(KEYINPUT22), .ZN(n829) );
  NOR2_X1 U920 ( .A1(G218), .A2(n829), .ZN(n830) );
  NAND2_X1 U921 ( .A1(G96), .A2(n830), .ZN(n843) );
  NAND2_X1 U922 ( .A1(n843), .A2(G2106), .ZN(n831) );
  NAND2_X1 U923 ( .A1(n832), .A2(n831), .ZN(n844) );
  NAND2_X1 U924 ( .A1(G483), .A2(G661), .ZN(n833) );
  NOR2_X1 U925 ( .A1(n844), .A2(n833), .ZN(n837) );
  NAND2_X1 U926 ( .A1(n837), .A2(G36), .ZN(G176) );
  NAND2_X1 U927 ( .A1(G2106), .A2(n834), .ZN(G217) );
  AND2_X1 U928 ( .A1(G15), .A2(G2), .ZN(n835) );
  NAND2_X1 U929 ( .A1(G661), .A2(n835), .ZN(G259) );
  NAND2_X1 U930 ( .A1(G3), .A2(G1), .ZN(n836) );
  NAND2_X1 U931 ( .A1(n837), .A2(n836), .ZN(G188) );
  XNOR2_X1 U933 ( .A(n1016), .B(n838), .ZN(n839) );
  NOR2_X1 U934 ( .A1(G860), .A2(n839), .ZN(n840) );
  XOR2_X1 U935 ( .A(n841), .B(n840), .Z(G145) );
  INV_X1 U936 ( .A(G132), .ZN(G219) );
  INV_X1 U937 ( .A(G108), .ZN(G238) );
  INV_X1 U938 ( .A(G82), .ZN(G220) );
  NOR2_X1 U939 ( .A1(n843), .A2(n842), .ZN(G325) );
  INV_X1 U940 ( .A(G325), .ZN(G261) );
  INV_X1 U941 ( .A(n844), .ZN(G319) );
  XOR2_X1 U942 ( .A(KEYINPUT42), .B(G2090), .Z(n846) );
  XNOR2_X1 U943 ( .A(G2072), .B(G2078), .ZN(n845) );
  XNOR2_X1 U944 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U945 ( .A(n847), .B(G2100), .Z(n849) );
  XNOR2_X1 U946 ( .A(G2067), .B(G2084), .ZN(n848) );
  XNOR2_X1 U947 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U948 ( .A(G2096), .B(KEYINPUT43), .Z(n851) );
  XNOR2_X1 U949 ( .A(KEYINPUT109), .B(G2678), .ZN(n850) );
  XNOR2_X1 U950 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U951 ( .A(n853), .B(n852), .Z(G227) );
  XOR2_X1 U952 ( .A(G1976), .B(G1971), .Z(n855) );
  XNOR2_X1 U953 ( .A(G1986), .B(G1966), .ZN(n854) );
  XNOR2_X1 U954 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U955 ( .A(n856), .B(G2474), .Z(n858) );
  XNOR2_X1 U956 ( .A(G1996), .B(G1991), .ZN(n857) );
  XNOR2_X1 U957 ( .A(n858), .B(n857), .ZN(n862) );
  XOR2_X1 U958 ( .A(KEYINPUT41), .B(G1981), .Z(n860) );
  XNOR2_X1 U959 ( .A(G1956), .B(G1961), .ZN(n859) );
  XNOR2_X1 U960 ( .A(n860), .B(n859), .ZN(n861) );
  XNOR2_X1 U961 ( .A(n862), .B(n861), .ZN(G229) );
  NAND2_X1 U962 ( .A1(G112), .A2(n895), .ZN(n863) );
  XNOR2_X1 U963 ( .A(n863), .B(KEYINPUT110), .ZN(n866) );
  NAND2_X1 U964 ( .A1(G124), .A2(n553), .ZN(n864) );
  XNOR2_X1 U965 ( .A(n864), .B(KEYINPUT44), .ZN(n865) );
  NAND2_X1 U966 ( .A1(n866), .A2(n865), .ZN(n870) );
  NAND2_X1 U967 ( .A1(G100), .A2(n891), .ZN(n868) );
  NAND2_X1 U968 ( .A1(G136), .A2(n892), .ZN(n867) );
  NAND2_X1 U969 ( .A1(n868), .A2(n867), .ZN(n869) );
  NOR2_X1 U970 ( .A1(n870), .A2(n869), .ZN(G162) );
  XOR2_X1 U971 ( .A(G160), .B(n871), .Z(n872) );
  XNOR2_X1 U972 ( .A(n959), .B(n872), .ZN(n886) );
  NAND2_X1 U973 ( .A1(n895), .A2(G118), .ZN(n873) );
  XNOR2_X1 U974 ( .A(KEYINPUT112), .B(n873), .ZN(n876) );
  NAND2_X1 U975 ( .A1(n553), .A2(G130), .ZN(n874) );
  XOR2_X1 U976 ( .A(KEYINPUT111), .B(n874), .Z(n875) );
  NAND2_X1 U977 ( .A1(n876), .A2(n875), .ZN(n877) );
  XNOR2_X1 U978 ( .A(n877), .B(KEYINPUT113), .ZN(n883) );
  NAND2_X1 U979 ( .A1(n891), .A2(G106), .ZN(n878) );
  XNOR2_X1 U980 ( .A(n878), .B(KEYINPUT114), .ZN(n880) );
  NAND2_X1 U981 ( .A1(G142), .A2(n892), .ZN(n879) );
  NAND2_X1 U982 ( .A1(n880), .A2(n879), .ZN(n881) );
  XNOR2_X1 U983 ( .A(KEYINPUT45), .B(n881), .ZN(n882) );
  NAND2_X1 U984 ( .A1(n883), .A2(n882), .ZN(n884) );
  XNOR2_X1 U985 ( .A(n884), .B(G162), .ZN(n885) );
  XNOR2_X1 U986 ( .A(n886), .B(n885), .ZN(n890) );
  XOR2_X1 U987 ( .A(n888), .B(n887), .Z(n889) );
  XNOR2_X1 U988 ( .A(n890), .B(n889), .ZN(n905) );
  XOR2_X1 U989 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n902) );
  NAND2_X1 U990 ( .A1(G103), .A2(n891), .ZN(n894) );
  NAND2_X1 U991 ( .A1(G139), .A2(n892), .ZN(n893) );
  NAND2_X1 U992 ( .A1(n894), .A2(n893), .ZN(n900) );
  NAND2_X1 U993 ( .A1(G127), .A2(n553), .ZN(n897) );
  NAND2_X1 U994 ( .A1(G115), .A2(n895), .ZN(n896) );
  NAND2_X1 U995 ( .A1(n897), .A2(n896), .ZN(n898) );
  XOR2_X1 U996 ( .A(KEYINPUT47), .B(n898), .Z(n899) );
  NOR2_X1 U997 ( .A1(n900), .A2(n899), .ZN(n970) );
  XNOR2_X1 U998 ( .A(n970), .B(KEYINPUT115), .ZN(n901) );
  XNOR2_X1 U999 ( .A(n902), .B(n901), .ZN(n903) );
  XNOR2_X1 U1000 ( .A(G164), .B(n903), .ZN(n904) );
  XNOR2_X1 U1001 ( .A(n905), .B(n904), .ZN(n906) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n906), .ZN(G395) );
  XNOR2_X1 U1003 ( .A(n907), .B(KEYINPUT116), .ZN(n910) );
  XNOR2_X1 U1004 ( .A(n908), .B(G286), .ZN(n909) );
  XNOR2_X1 U1005 ( .A(n910), .B(n909), .ZN(n911) );
  XOR2_X1 U1006 ( .A(G171), .B(n911), .Z(n912) );
  NOR2_X1 U1007 ( .A1(G37), .A2(n912), .ZN(G397) );
  XOR2_X1 U1008 ( .A(G2438), .B(KEYINPUT108), .Z(n914) );
  XNOR2_X1 U1009 ( .A(G2443), .B(G2430), .ZN(n913) );
  XNOR2_X1 U1010 ( .A(n914), .B(n913), .ZN(n915) );
  XOR2_X1 U1011 ( .A(n915), .B(G2435), .Z(n917) );
  XNOR2_X1 U1012 ( .A(G1341), .B(G1348), .ZN(n916) );
  XNOR2_X1 U1013 ( .A(n917), .B(n916), .ZN(n921) );
  XOR2_X1 U1014 ( .A(G2451), .B(G2427), .Z(n919) );
  XNOR2_X1 U1015 ( .A(G2454), .B(G2446), .ZN(n918) );
  XNOR2_X1 U1016 ( .A(n919), .B(n918), .ZN(n920) );
  XOR2_X1 U1017 ( .A(n921), .B(n920), .Z(n922) );
  NAND2_X1 U1018 ( .A1(G14), .A2(n922), .ZN(n928) );
  NAND2_X1 U1019 ( .A1(G319), .A2(n928), .ZN(n925) );
  NOR2_X1 U1020 ( .A1(G227), .A2(G229), .ZN(n923) );
  XNOR2_X1 U1021 ( .A(KEYINPUT49), .B(n923), .ZN(n924) );
  NOR2_X1 U1022 ( .A1(n925), .A2(n924), .ZN(n927) );
  NOR2_X1 U1023 ( .A1(G395), .A2(G397), .ZN(n926) );
  NAND2_X1 U1024 ( .A1(n927), .A2(n926), .ZN(G225) );
  INV_X1 U1025 ( .A(G225), .ZN(G308) );
  INV_X1 U1026 ( .A(G96), .ZN(G221) );
  INV_X1 U1027 ( .A(G69), .ZN(G235) );
  INV_X1 U1028 ( .A(n928), .ZN(G401) );
  XNOR2_X1 U1029 ( .A(n929), .B(G5), .ZN(n948) );
  XNOR2_X1 U1030 ( .A(KEYINPUT59), .B(G4), .ZN(n930) );
  XNOR2_X1 U1031 ( .A(n930), .B(KEYINPUT125), .ZN(n931) );
  XNOR2_X1 U1032 ( .A(G1348), .B(n931), .ZN(n933) );
  XNOR2_X1 U1033 ( .A(G1981), .B(G6), .ZN(n932) );
  NOR2_X1 U1034 ( .A1(n933), .A2(n932), .ZN(n937) );
  XNOR2_X1 U1035 ( .A(G1956), .B(G20), .ZN(n935) );
  XNOR2_X1 U1036 ( .A(G19), .B(G1341), .ZN(n934) );
  NOR2_X1 U1037 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1038 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1039 ( .A(n938), .B(KEYINPUT60), .ZN(n946) );
  XNOR2_X1 U1040 ( .A(G1986), .B(G24), .ZN(n940) );
  XNOR2_X1 U1041 ( .A(G1971), .B(G22), .ZN(n939) );
  NOR2_X1 U1042 ( .A1(n940), .A2(n939), .ZN(n943) );
  XOR2_X1 U1043 ( .A(G1976), .B(KEYINPUT126), .Z(n941) );
  XNOR2_X1 U1044 ( .A(G23), .B(n941), .ZN(n942) );
  NAND2_X1 U1045 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1046 ( .A(KEYINPUT58), .B(n944), .ZN(n945) );
  NOR2_X1 U1047 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1048 ( .A1(n948), .A2(n947), .ZN(n950) );
  XNOR2_X1 U1049 ( .A(G21), .B(G1966), .ZN(n949) );
  NOR2_X1 U1050 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1051 ( .A(KEYINPUT61), .B(n951), .ZN(n953) );
  INV_X1 U1052 ( .A(G16), .ZN(n952) );
  NAND2_X1 U1053 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1054 ( .A1(n954), .A2(G11), .ZN(n1035) );
  XNOR2_X1 U1055 ( .A(G2090), .B(G162), .ZN(n955) );
  XNOR2_X1 U1056 ( .A(n955), .B(KEYINPUT118), .ZN(n956) );
  NAND2_X1 U1057 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1058 ( .A(n958), .B(KEYINPUT51), .ZN(n969) );
  XNOR2_X1 U1059 ( .A(G160), .B(G2084), .ZN(n960) );
  NAND2_X1 U1060 ( .A1(n960), .A2(n959), .ZN(n961) );
  NOR2_X1 U1061 ( .A1(n962), .A2(n961), .ZN(n966) );
  NOR2_X1 U1062 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1063 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1064 ( .A(KEYINPUT117), .B(n967), .ZN(n968) );
  NAND2_X1 U1065 ( .A1(n969), .A2(n968), .ZN(n978) );
  XOR2_X1 U1066 ( .A(G164), .B(G2078), .Z(n973) );
  XNOR2_X1 U1067 ( .A(n971), .B(n970), .ZN(n972) );
  NOR2_X1 U1068 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1069 ( .A(n974), .B(KEYINPUT50), .ZN(n976) );
  NAND2_X1 U1070 ( .A1(n976), .A2(n975), .ZN(n977) );
  NOR2_X1 U1071 ( .A1(n978), .A2(n977), .ZN(n979) );
  XOR2_X1 U1072 ( .A(KEYINPUT52), .B(n979), .Z(n980) );
  NOR2_X1 U1073 ( .A1(KEYINPUT55), .A2(n980), .ZN(n981) );
  XNOR2_X1 U1074 ( .A(KEYINPUT119), .B(n981), .ZN(n982) );
  NAND2_X1 U1075 ( .A1(n982), .A2(G29), .ZN(n1033) );
  XNOR2_X1 U1076 ( .A(G32), .B(n983), .ZN(n988) );
  XNOR2_X1 U1077 ( .A(G2067), .B(G26), .ZN(n986) );
  XNOR2_X1 U1078 ( .A(G27), .B(n984), .ZN(n985) );
  NOR2_X1 U1079 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1080 ( .A1(n988), .A2(n987), .ZN(n990) );
  XNOR2_X1 U1081 ( .A(G33), .B(G2072), .ZN(n989) );
  NOR2_X1 U1082 ( .A1(n990), .A2(n989), .ZN(n991) );
  XOR2_X1 U1083 ( .A(KEYINPUT120), .B(n991), .Z(n993) );
  XNOR2_X1 U1084 ( .A(G1991), .B(G25), .ZN(n992) );
  NOR2_X1 U1085 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1086 ( .A1(G28), .A2(n994), .ZN(n995) );
  XNOR2_X1 U1087 ( .A(n995), .B(KEYINPUT53), .ZN(n998) );
  XOR2_X1 U1088 ( .A(G2084), .B(G34), .Z(n996) );
  XNOR2_X1 U1089 ( .A(KEYINPUT54), .B(n996), .ZN(n997) );
  NAND2_X1 U1090 ( .A1(n998), .A2(n997), .ZN(n1000) );
  XNOR2_X1 U1091 ( .A(G35), .B(G2090), .ZN(n999) );
  NOR2_X1 U1092 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XOR2_X1 U1093 ( .A(KEYINPUT55), .B(n1001), .Z(n1002) );
  NOR2_X1 U1094 ( .A1(G29), .A2(n1002), .ZN(n1003) );
  XOR2_X1 U1095 ( .A(KEYINPUT121), .B(n1003), .Z(n1031) );
  XOR2_X1 U1096 ( .A(G16), .B(KEYINPUT56), .Z(n1028) );
  XOR2_X1 U1097 ( .A(G1961), .B(G171), .Z(n1004) );
  NOR2_X1 U1098 ( .A1(n1005), .A2(n1004), .ZN(n1007) );
  NAND2_X1 U1099 ( .A1(n1007), .A2(n1006), .ZN(n1025) );
  XNOR2_X1 U1100 ( .A(G1971), .B(G166), .ZN(n1008) );
  XNOR2_X1 U1101 ( .A(n1008), .B(KEYINPUT122), .ZN(n1013) );
  XNOR2_X1 U1102 ( .A(n1009), .B(G1348), .ZN(n1011) );
  XNOR2_X1 U1103 ( .A(G299), .B(G1956), .ZN(n1010) );
  NOR2_X1 U1104 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1105 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NOR2_X1 U1106 ( .A1(n1015), .A2(n1014), .ZN(n1023) );
  XNOR2_X1 U1107 ( .A(n1016), .B(G1341), .ZN(n1021) );
  XOR2_X1 U1108 ( .A(G1966), .B(G168), .Z(n1017) );
  NOR2_X1 U1109 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1110 ( .A(KEYINPUT57), .B(n1019), .ZN(n1020) );
  NOR2_X1 U1111 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1112 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NOR2_X1 U1113 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XOR2_X1 U1114 ( .A(KEYINPUT123), .B(n1026), .Z(n1027) );
  NOR2_X1 U1115 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XNOR2_X1 U1116 ( .A(KEYINPUT124), .B(n1029), .ZN(n1030) );
  NOR2_X1 U1117 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NAND2_X1 U1118 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NOR2_X1 U1119 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  XOR2_X1 U1120 ( .A(KEYINPUT62), .B(n1036), .Z(n1037) );
  XNOR2_X1 U1121 ( .A(KEYINPUT127), .B(n1037), .ZN(G311) );
  INV_X1 U1122 ( .A(G311), .ZN(G150) );
endmodule

