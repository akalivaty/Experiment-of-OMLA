//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 0 0 0 1 0 0 1 1 0 1 1 1 0 0 1 1 0 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 0 0 0 1 0 0 1 1 1 1 0 1 0 0 0 0 1 0 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:26 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n550, new_n552,
    new_n553, new_n554, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n572, new_n574, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n600, new_n601, new_n604,
    new_n605, new_n607, new_n608, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  XNOR2_X1  g031(.A(G325), .B(KEYINPUT64), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT65), .ZN(G319));
  NAND2_X1  g034(.A1(G101), .A2(G2104), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT66), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  OAI21_X1  g037(.A(new_n461), .B1(new_n462), .B2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n464), .A2(KEYINPUT66), .A3(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G137), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n460), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n464), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n467), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G125), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n473), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G2105), .ZN(new_n478));
  AND2_X1   g053(.A1(new_n472), .A2(new_n478), .ZN(G160));
  AOI22_X1  g054(.A1(new_n463), .A2(new_n465), .B1(KEYINPUT3), .B2(new_n462), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(new_n471), .ZN(new_n481));
  INV_X1    g056(.A(G136), .ZN(new_n482));
  NOR2_X1   g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(new_n471), .B2(G112), .ZN(new_n484));
  OAI22_X1  g059(.A1(new_n481), .A2(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n480), .A2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n485), .B1(G124), .B2(new_n487), .ZN(G162));
  NAND4_X1  g063(.A1(new_n467), .A2(new_n474), .A3(G138), .A4(new_n471), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n462), .A2(G2105), .ZN(new_n491));
  AOI22_X1  g066(.A1(new_n489), .A2(new_n490), .B1(G102), .B2(new_n491), .ZN(new_n492));
  AND2_X1   g067(.A1(KEYINPUT4), .A2(G138), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n466), .A2(new_n471), .A3(new_n467), .A4(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  AND3_X1   g070(.A1(new_n464), .A2(KEYINPUT66), .A3(G2104), .ZN(new_n496));
  AOI21_X1  g071(.A(KEYINPUT66), .B1(new_n464), .B2(G2104), .ZN(new_n497));
  OAI211_X1 g072(.A(G126), .B(new_n467), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  XNOR2_X1  g073(.A(KEYINPUT67), .B(G114), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(G2104), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n471), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n495), .A2(new_n501), .ZN(G164));
  NAND2_X1  g077(.A1(G75), .A2(G543), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT5), .ZN(new_n504));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n504), .B1(new_n505), .B2(KEYINPUT69), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT69), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n507), .A2(KEYINPUT5), .A3(G543), .ZN(new_n508));
  AND2_X1   g083(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G62), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n503), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G651), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT6), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G651), .ZN(new_n514));
  XNOR2_X1  g089(.A(new_n514), .B(KEYINPUT68), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n506), .A2(new_n508), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(KEYINPUT6), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n515), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G88), .ZN(new_n520));
  INV_X1    g095(.A(G50), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n515), .A2(G543), .A3(new_n518), .ZN(new_n522));
  OAI221_X1 g097(.A(new_n512), .B1(new_n519), .B2(new_n520), .C1(new_n521), .C2(new_n522), .ZN(G303));
  INV_X1    g098(.A(G303), .ZN(G166));
  INV_X1    g099(.A(new_n522), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G51), .ZN(new_n526));
  INV_X1    g101(.A(new_n519), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G89), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n516), .A2(G63), .A3(G651), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT7), .ZN(new_n531));
  NAND4_X1  g106(.A1(new_n526), .A2(new_n528), .A3(new_n529), .A4(new_n531), .ZN(G286));
  INV_X1    g107(.A(G286), .ZN(G168));
  NAND2_X1  g108(.A1(G77), .A2(G543), .ZN(new_n534));
  INV_X1    g109(.A(G64), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n534), .B1(new_n509), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G651), .ZN(new_n537));
  INV_X1    g112(.A(G90), .ZN(new_n538));
  INV_X1    g113(.A(G52), .ZN(new_n539));
  OAI221_X1 g114(.A(new_n537), .B1(new_n519), .B2(new_n538), .C1(new_n539), .C2(new_n522), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT70), .ZN(G171));
  INV_X1    g116(.A(G43), .ZN(new_n542));
  INV_X1    g117(.A(G81), .ZN(new_n543));
  OAI22_X1  g118(.A1(new_n542), .A2(new_n522), .B1(new_n519), .B2(new_n543), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT71), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n516), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n546), .A2(new_n517), .ZN(new_n547));
  AND2_X1   g122(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  AND3_X1   g124(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G36), .ZN(G176));
  XOR2_X1   g126(.A(KEYINPUT72), .B(KEYINPUT8), .Z(new_n552));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n552), .B(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n550), .A2(new_n554), .ZN(G188));
  XNOR2_X1  g130(.A(new_n516), .B(KEYINPUT74), .ZN(new_n556));
  INV_X1    g131(.A(G65), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  AND2_X1   g133(.A1(G78), .A2(G543), .ZN(new_n559));
  OAI21_X1  g134(.A(G651), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT75), .ZN(new_n561));
  OR2_X1    g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n560), .A2(new_n561), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n562), .A2(new_n563), .B1(G91), .B2(new_n527), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n525), .A2(KEYINPUT9), .A3(G53), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT9), .ZN(new_n566));
  INV_X1    g141(.A(G53), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n566), .B1(new_n522), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  XOR2_X1   g144(.A(new_n569), .B(KEYINPUT73), .Z(new_n570));
  NAND2_X1  g145(.A1(new_n564), .A2(new_n570), .ZN(G299));
  INV_X1    g146(.A(KEYINPUT70), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n540), .B(new_n572), .ZN(G301));
  NAND4_X1  g148(.A1(new_n515), .A2(G49), .A3(G543), .A4(new_n518), .ZN(new_n574));
  OAI21_X1  g149(.A(G651), .B1(new_n516), .B2(G74), .ZN(new_n575));
  INV_X1    g150(.A(G87), .ZN(new_n576));
  OAI211_X1 g151(.A(new_n574), .B(new_n575), .C1(new_n519), .C2(new_n576), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n577), .B(KEYINPUT76), .ZN(G288));
  NAND2_X1  g153(.A1(new_n525), .A2(G48), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n527), .A2(G86), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n516), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n581));
  OR2_X1    g156(.A1(new_n581), .A2(new_n517), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n579), .A2(new_n580), .A3(new_n582), .ZN(G305));
  NAND2_X1  g158(.A1(new_n527), .A2(G85), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n525), .A2(G47), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n516), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n586));
  OAI211_X1 g161(.A(new_n584), .B(new_n585), .C1(new_n517), .C2(new_n586), .ZN(G290));
  NAND2_X1  g162(.A1(G301), .A2(G868), .ZN(new_n588));
  INV_X1    g163(.A(G66), .ZN(new_n589));
  OR2_X1    g164(.A1(new_n556), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(G79), .A2(G543), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n517), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n592), .B1(G54), .B2(new_n525), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n527), .A2(G92), .ZN(new_n594));
  XOR2_X1   g169(.A(new_n594), .B(KEYINPUT10), .Z(new_n595));
  NAND2_X1  g170(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n588), .B1(new_n597), .B2(G868), .ZN(G284));
  OAI21_X1  g173(.A(new_n588), .B1(new_n597), .B2(G868), .ZN(G321));
  NAND2_X1  g174(.A1(G286), .A2(G868), .ZN(new_n600));
  INV_X1    g175(.A(G299), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n601), .B2(G868), .ZN(G297));
  OAI21_X1  g177(.A(new_n600), .B1(new_n601), .B2(G868), .ZN(G280));
  INV_X1    g178(.A(G559), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n597), .B1(new_n604), .B2(G860), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n605), .B(KEYINPUT77), .ZN(G148));
  NAND2_X1  g181(.A1(new_n597), .A2(new_n604), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n607), .A2(G868), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(G868), .B2(new_n548), .ZN(G323));
  XNOR2_X1  g184(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g185(.A1(new_n487), .A2(G123), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n468), .A2(G2105), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(G135), .ZN(new_n613));
  NOR2_X1   g188(.A1(G99), .A2(G2105), .ZN(new_n614));
  OAI21_X1  g189(.A(G2104), .B1(new_n471), .B2(G111), .ZN(new_n615));
  OAI211_X1 g190(.A(new_n611), .B(new_n613), .C1(new_n614), .C2(new_n615), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(G2096), .Z(new_n617));
  NAND3_X1  g192(.A1(new_n471), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(KEYINPUT12), .Z(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT13), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(G2100), .Z(new_n621));
  NAND2_X1  g196(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(KEYINPUT78), .Z(G156));
  XNOR2_X1  g198(.A(KEYINPUT15), .B(G2430), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2435), .ZN(new_n625));
  XOR2_X1   g200(.A(G2427), .B(G2438), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(KEYINPUT14), .ZN(new_n628));
  XOR2_X1   g203(.A(G2451), .B(G2454), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT16), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n628), .B(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(G1341), .B(G1348), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2443), .B(G2446), .ZN(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n633), .B(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(G14), .ZN(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(G401));
  XNOR2_X1  g213(.A(G2072), .B(G2078), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT17), .Z(new_n640));
  XOR2_X1   g215(.A(G2084), .B(G2090), .Z(new_n641));
  XNOR2_X1  g216(.A(G2067), .B(G2678), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n640), .A2(new_n641), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT79), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n640), .A2(new_n643), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n646), .A2(new_n641), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n647), .B1(new_n639), .B2(new_n642), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n641), .A2(new_n639), .A3(new_n642), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(KEYINPUT18), .Z(new_n650));
  NAND3_X1  g225(.A1(new_n645), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2096), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2100), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(G227));
  XOR2_X1   g229(.A(G1956), .B(G2474), .Z(new_n655));
  XOR2_X1   g230(.A(G1961), .B(G1966), .Z(new_n656));
  NOR2_X1   g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1971), .B(G1976), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT19), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n655), .A2(new_n656), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(KEYINPUT20), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n661), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n658), .A2(new_n660), .A3(new_n662), .ZN(new_n666));
  OAI211_X1 g241(.A(new_n665), .B(new_n666), .C1(new_n664), .C2(new_n663), .ZN(new_n667));
  XOR2_X1   g242(.A(KEYINPUT21), .B(G1986), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(G1991), .B(G1996), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT22), .B(G1981), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n671), .B(new_n672), .Z(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(G229));
  XNOR2_X1  g249(.A(KEYINPUT89), .B(KEYINPUT24), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(G34), .ZN(new_n676));
  MUX2_X1   g251(.A(new_n676), .B(G160), .S(G29), .Z(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(KEYINPUT90), .Z(new_n678));
  INV_X1    g253(.A(G2084), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n680), .B(KEYINPUT92), .Z(new_n681));
  INV_X1    g256(.A(G16), .ZN(new_n682));
  NOR2_X1   g257(.A1(G171), .A2(new_n682), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n683), .B1(G5), .B2(new_n682), .ZN(new_n684));
  INV_X1    g259(.A(G1961), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n678), .A2(new_n679), .ZN(new_n687));
  INV_X1    g262(.A(KEYINPUT30), .ZN(new_n688));
  AND2_X1   g263(.A1(new_n688), .A2(G28), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n688), .A2(G28), .ZN(new_n690));
  NOR3_X1   g265(.A1(new_n689), .A2(new_n690), .A3(G29), .ZN(new_n691));
  INV_X1    g266(.A(G29), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n616), .A2(new_n692), .ZN(new_n693));
  NOR4_X1   g268(.A1(new_n686), .A2(new_n687), .A3(new_n691), .A4(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n684), .A2(new_n685), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n681), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  NOR2_X1   g271(.A1(G29), .A2(G33), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n612), .A2(G139), .ZN(new_n698));
  NAND2_X1  g273(.A1(G115), .A2(G2104), .ZN(new_n699));
  INV_X1    g274(.A(G127), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n699), .B1(new_n475), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G2105), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n491), .A2(G103), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT25), .Z(new_n704));
  NAND3_X1  g279(.A1(new_n698), .A2(new_n702), .A3(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n697), .B1(new_n706), .B2(G29), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(G2072), .ZN(new_n708));
  XOR2_X1   g283(.A(KEYINPUT31), .B(G11), .Z(new_n709));
  NAND2_X1  g284(.A1(new_n692), .A2(G27), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(G164), .B2(new_n692), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(G2078), .ZN(new_n712));
  NOR4_X1   g287(.A1(new_n696), .A2(new_n708), .A3(new_n709), .A4(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n682), .A2(G4), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(new_n597), .B2(new_n682), .ZN(new_n715));
  INV_X1    g290(.A(G1348), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n682), .A2(G19), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(new_n548), .B2(new_n682), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(G1341), .Z(new_n720));
  NOR2_X1   g295(.A1(G104), .A2(G2105), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT86), .ZN(new_n722));
  OAI211_X1 g297(.A(new_n722), .B(G2104), .C1(G116), .C2(new_n471), .ZN(new_n723));
  INV_X1    g298(.A(G128), .ZN(new_n724));
  INV_X1    g299(.A(G140), .ZN(new_n725));
  OAI221_X1 g300(.A(new_n723), .B1(new_n486), .B2(new_n724), .C1(new_n725), .C2(new_n481), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(G29), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT87), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n692), .A2(G26), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT28), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(G2067), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n717), .A2(new_n720), .A3(new_n733), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT88), .Z(new_n735));
  NAND3_X1  g310(.A1(new_n682), .A2(KEYINPUT23), .A3(G20), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT23), .ZN(new_n737));
  INV_X1    g312(.A(G20), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n737), .B1(new_n738), .B2(G16), .ZN(new_n739));
  OAI211_X1 g314(.A(new_n736), .B(new_n739), .C1(new_n601), .C2(new_n682), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT93), .ZN(new_n741));
  INV_X1    g316(.A(G1956), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n713), .A2(new_n735), .A3(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT84), .ZN(new_n745));
  MUX2_X1   g320(.A(G24), .B(G290), .S(G16), .Z(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(G1986), .Z(new_n747));
  NOR2_X1   g322(.A1(G16), .A2(G23), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT81), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n577), .B(new_n749), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n748), .B1(new_n750), .B2(G16), .ZN(new_n751));
  XNOR2_X1  g326(.A(KEYINPUT33), .B(G1976), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  MUX2_X1   g328(.A(G6), .B(G305), .S(G16), .Z(new_n754));
  XOR2_X1   g329(.A(KEYINPUT32), .B(G1981), .Z(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(G22), .ZN(new_n757));
  OAI21_X1  g332(.A(KEYINPUT82), .B1(new_n757), .B2(G16), .ZN(new_n758));
  OR3_X1    g333(.A1(new_n757), .A2(KEYINPUT82), .A3(G16), .ZN(new_n759));
  OAI211_X1 g334(.A(new_n758), .B(new_n759), .C1(G166), .C2(new_n682), .ZN(new_n760));
  INV_X1    g335(.A(G1971), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n753), .A2(new_n756), .A3(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n763), .A2(KEYINPUT34), .ZN(new_n764));
  INV_X1    g339(.A(new_n764), .ZN(new_n765));
  AND2_X1   g340(.A1(new_n763), .A2(KEYINPUT34), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n766), .A2(KEYINPUT83), .ZN(new_n767));
  INV_X1    g342(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n766), .A2(KEYINPUT83), .ZN(new_n769));
  OAI211_X1 g344(.A(new_n747), .B(new_n765), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n692), .A2(G25), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n487), .A2(G119), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n612), .A2(KEYINPUT80), .A3(G131), .ZN(new_n773));
  OR2_X1    g348(.A1(G95), .A2(G2105), .ZN(new_n774));
  OAI211_X1 g349(.A(new_n774), .B(G2104), .C1(G107), .C2(new_n471), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT80), .ZN(new_n776));
  INV_X1    g351(.A(G131), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n776), .B1(new_n481), .B2(new_n777), .ZN(new_n778));
  AND4_X1   g353(.A1(new_n772), .A2(new_n773), .A3(new_n775), .A4(new_n778), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n771), .B1(new_n779), .B2(new_n692), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT35), .B(G1991), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n745), .B1(new_n770), .B2(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(new_n769), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n764), .B1(new_n784), .B2(new_n767), .ZN(new_n785));
  INV_X1    g360(.A(new_n782), .ZN(new_n786));
  NAND4_X1  g361(.A1(new_n785), .A2(KEYINPUT84), .A3(new_n747), .A4(new_n786), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n783), .A2(new_n787), .A3(KEYINPUT36), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n785), .A2(new_n747), .A3(new_n786), .ZN(new_n789));
  OAI21_X1  g364(.A(KEYINPUT85), .B1(new_n789), .B2(KEYINPUT36), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  NAND4_X1  g366(.A1(new_n783), .A2(new_n787), .A3(KEYINPUT85), .A4(KEYINPUT36), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n744), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n487), .A2(G129), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n612), .A2(G141), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n491), .A2(G105), .ZN(new_n796));
  NAND3_X1  g371(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT26), .Z(new_n798));
  NAND4_X1  g373(.A1(new_n794), .A2(new_n795), .A3(new_n796), .A4(new_n798), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n799), .A2(new_n692), .ZN(new_n800));
  INV_X1    g375(.A(KEYINPUT91), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  OAI21_X1  g377(.A(KEYINPUT91), .B1(G29), .B2(G32), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n802), .B1(new_n800), .B2(new_n803), .ZN(new_n804));
  XNOR2_X1  g379(.A(KEYINPUT27), .B(G1996), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n682), .A2(G21), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G168), .B2(new_n682), .ZN(new_n808));
  INV_X1    g383(.A(G1966), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NOR2_X1   g385(.A1(G29), .A2(G35), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n811), .B1(G162), .B2(G29), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT29), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(G2090), .Z(new_n814));
  NAND4_X1  g389(.A1(new_n793), .A2(new_n806), .A3(new_n810), .A4(new_n814), .ZN(G150));
  INV_X1    g390(.A(G150), .ZN(G311));
  NAND2_X1  g391(.A1(new_n527), .A2(G93), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n525), .A2(G55), .ZN(new_n818));
  AOI22_X1  g393(.A1(new_n516), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n819));
  OAI211_X1 g394(.A(new_n817), .B(new_n818), .C1(new_n517), .C2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n820), .A2(G860), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(KEYINPUT37), .Z(new_n822));
  NOR2_X1   g397(.A1(new_n596), .A2(new_n604), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT39), .ZN(new_n824));
  XNOR2_X1  g399(.A(KEYINPUT94), .B(KEYINPUT38), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n545), .A2(new_n547), .A3(new_n820), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n820), .B1(new_n545), .B2(new_n547), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n826), .B(new_n830), .Z(new_n831));
  OAI21_X1  g406(.A(new_n822), .B1(new_n831), .B2(G860), .ZN(G145));
  XOR2_X1   g407(.A(G160), .B(new_n616), .Z(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(G162), .Z(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  OR2_X1    g410(.A1(new_n726), .A2(G164), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n726), .A2(G164), .ZN(new_n837));
  AND3_X1   g412(.A1(new_n836), .A2(new_n799), .A3(new_n837), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n799), .B1(new_n836), .B2(new_n837), .ZN(new_n839));
  OR3_X1    g414(.A1(new_n838), .A2(new_n839), .A3(new_n705), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n705), .B1(new_n838), .B2(new_n839), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n487), .A2(G130), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n612), .A2(G142), .ZN(new_n844));
  OR2_X1    g419(.A1(G106), .A2(G2105), .ZN(new_n845));
  OAI211_X1 g420(.A(new_n845), .B(G2104), .C1(G118), .C2(new_n471), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n843), .A2(new_n844), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n779), .A2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n847), .ZN(new_n849));
  NAND4_X1  g424(.A1(new_n773), .A2(new_n772), .A3(new_n778), .A4(new_n775), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n848), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n852), .A2(KEYINPUT95), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT95), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n848), .A2(new_n854), .A3(new_n851), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n853), .A2(new_n619), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n853), .A2(new_n855), .ZN(new_n857));
  INV_X1    g432(.A(new_n619), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n842), .A2(new_n856), .A3(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT96), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n859), .A2(new_n856), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(new_n842), .ZN(new_n864));
  OAI211_X1 g439(.A(new_n835), .B(new_n862), .C1(new_n864), .C2(new_n861), .ZN(new_n865));
  OR2_X1    g440(.A1(new_n864), .A2(new_n835), .ZN(new_n866));
  INV_X1    g441(.A(G37), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT97), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND4_X1  g445(.A1(new_n865), .A2(new_n866), .A3(KEYINPUT97), .A4(new_n867), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  OR2_X1    g447(.A1(new_n872), .A2(KEYINPUT98), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(KEYINPUT98), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g451(.A1(new_n820), .A2(G868), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n750), .B(G290), .ZN(new_n878));
  XNOR2_X1  g453(.A(G166), .B(G305), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n878), .B(new_n879), .ZN(new_n880));
  XOR2_X1   g455(.A(new_n880), .B(KEYINPUT42), .Z(new_n881));
  XNOR2_X1  g456(.A(new_n607), .B(new_n830), .ZN(new_n882));
  NAND2_X1  g457(.A1(G299), .A2(new_n596), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n597), .A2(new_n564), .A3(new_n570), .ZN(new_n884));
  AND3_X1   g459(.A1(new_n883), .A2(new_n884), .A3(KEYINPUT99), .ZN(new_n885));
  AOI21_X1  g460(.A(KEYINPUT99), .B1(new_n883), .B2(new_n884), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n882), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n883), .A2(new_n884), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT41), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n883), .A2(new_n884), .A3(KEYINPUT41), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n887), .B1(new_n892), .B2(new_n882), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n881), .B1(new_n893), .B2(KEYINPUT100), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n893), .A2(KEYINPUT100), .ZN(new_n895));
  MUX2_X1   g470(.A(new_n894), .B(new_n881), .S(new_n895), .Z(new_n896));
  AOI21_X1  g471(.A(new_n877), .B1(new_n896), .B2(G868), .ZN(G295));
  AOI21_X1  g472(.A(new_n877), .B1(new_n896), .B2(G868), .ZN(G331));
  OR2_X1    g473(.A1(G286), .A2(KEYINPUT101), .ZN(new_n899));
  NAND2_X1  g474(.A1(G286), .A2(KEYINPUT101), .ZN(new_n900));
  NAND3_X1  g475(.A1(G171), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(G301), .A2(KEYINPUT101), .A3(G286), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(new_n830), .ZN(new_n904));
  OAI211_X1 g479(.A(new_n901), .B(new_n902), .C1(new_n828), .C2(new_n829), .ZN(new_n905));
  AOI21_X1  g480(.A(KEYINPUT102), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AND2_X1   g481(.A1(new_n905), .A2(KEYINPUT102), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n888), .ZN(new_n909));
  AND3_X1   g484(.A1(new_n883), .A2(new_n884), .A3(KEYINPUT41), .ZN(new_n910));
  AOI21_X1  g485(.A(KEYINPUT41), .B1(new_n883), .B2(new_n884), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n904), .A2(new_n905), .ZN(new_n913));
  AOI22_X1  g488(.A1(new_n908), .A2(new_n909), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(G37), .B1(new_n914), .B2(new_n880), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT43), .ZN(new_n916));
  OAI211_X1 g491(.A(new_n890), .B(new_n891), .C1(new_n906), .C2(new_n907), .ZN(new_n917));
  INV_X1    g492(.A(new_n913), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n918), .B1(new_n886), .B2(new_n885), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n880), .ZN(new_n921));
  AOI21_X1  g496(.A(KEYINPUT103), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT103), .ZN(new_n923));
  AOI211_X1 g498(.A(new_n923), .B(new_n880), .C1(new_n917), .C2(new_n919), .ZN(new_n924));
  OAI211_X1 g499(.A(new_n915), .B(new_n916), .C1(new_n922), .C2(new_n924), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n892), .A2(new_n918), .ZN(new_n926));
  NOR3_X1   g501(.A1(new_n906), .A2(new_n907), .A3(new_n888), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n921), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n927), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n912), .A2(new_n913), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n929), .A2(new_n880), .A3(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n928), .A2(new_n931), .A3(new_n867), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(KEYINPUT43), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n925), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n932), .A2(new_n916), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n915), .B1(new_n922), .B2(new_n924), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n935), .B1(new_n936), .B2(new_n916), .ZN(new_n937));
  MUX2_X1   g512(.A(new_n934), .B(new_n937), .S(KEYINPUT44), .Z(G397));
  INV_X1    g513(.A(G1384), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n939), .B1(new_n495), .B2(new_n501), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  OR2_X1    g516(.A1(new_n941), .A2(KEYINPUT45), .ZN(new_n942));
  AND3_X1   g517(.A1(new_n472), .A2(G40), .A3(new_n478), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(G1996), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n947), .A2(new_n799), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n945), .B(KEYINPUT104), .ZN(new_n949));
  INV_X1    g524(.A(new_n949), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n726), .B(G2067), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n951), .B(KEYINPUT105), .ZN(new_n952));
  INV_X1    g527(.A(new_n799), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n952), .B1(new_n946), .B2(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n948), .B1(new_n950), .B2(new_n954), .ZN(new_n955));
  XOR2_X1   g530(.A(new_n850), .B(new_n781), .Z(new_n956));
  OAI21_X1  g531(.A(new_n955), .B1(new_n956), .B2(new_n949), .ZN(new_n957));
  XNOR2_X1  g532(.A(G290), .B(G1986), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n957), .B1(new_n945), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(G286), .A2(G8), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  OR2_X1    g536(.A1(new_n961), .A2(KEYINPUT51), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n944), .B1(KEYINPUT50), .B2(new_n940), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT106), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n940), .A2(new_n964), .ZN(new_n965));
  OAI211_X1 g540(.A(KEYINPUT106), .B(new_n939), .C1(new_n495), .C2(new_n501), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n963), .B1(new_n968), .B2(KEYINPUT50), .ZN(new_n969));
  XNOR2_X1  g544(.A(KEYINPUT113), .B(G2084), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  AOI22_X1  g548(.A1(new_n480), .A2(G126), .B1(G2104), .B2(new_n499), .ZN(new_n974));
  OAI211_X1 g549(.A(new_n494), .B(new_n492), .C1(new_n974), .C2(new_n471), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT106), .B1(new_n975), .B2(new_n939), .ZN(new_n976));
  INV_X1    g551(.A(new_n966), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n943), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n943), .A2(KEYINPUT45), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n978), .A2(KEYINPUT111), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n941), .A2(KEYINPUT45), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT111), .ZN(new_n982));
  OAI211_X1 g557(.A(new_n982), .B(new_n943), .C1(new_n967), .C2(KEYINPUT45), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n980), .A2(new_n981), .A3(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT112), .ZN(new_n985));
  AND3_X1   g560(.A1(new_n984), .A2(new_n985), .A3(new_n809), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n985), .B1(new_n984), .B2(new_n809), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n973), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n962), .B1(new_n988), .B2(G8), .ZN(new_n989));
  XOR2_X1   g564(.A(new_n960), .B(KEYINPUT118), .Z(new_n990));
  NAND2_X1  g565(.A1(new_n984), .A2(new_n809), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(KEYINPUT112), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n984), .A2(new_n985), .A3(new_n809), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n972), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(G8), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n990), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  XNOR2_X1  g571(.A(KEYINPUT117), .B(KEYINPUT51), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n989), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n994), .A2(new_n960), .ZN(new_n1000));
  OAI21_X1  g575(.A(KEYINPUT119), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT62), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT119), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1000), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n988), .A2(G8), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n997), .B1(new_n1005), .B2(new_n990), .ZN(new_n1006));
  OAI211_X1 g581(.A(new_n1003), .B(new_n1004), .C1(new_n1006), .C2(new_n989), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1001), .A2(new_n1002), .A3(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n942), .A2(new_n943), .A3(new_n981), .ZN(new_n1009));
  OR2_X1    g584(.A1(new_n1009), .A2(G2078), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT53), .ZN(new_n1011));
  AOI22_X1  g586(.A1(new_n1010), .A2(new_n1011), .B1(new_n969), .B2(new_n685), .ZN(new_n1012));
  OR2_X1    g587(.A1(new_n1011), .A2(G2078), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1012), .B1(new_n984), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(G171), .ZN(new_n1015));
  OR2_X1    g590(.A1(G305), .A2(G1981), .ZN(new_n1016));
  NAND2_X1  g591(.A1(G305), .A2(G1981), .ZN(new_n1017));
  AOI21_X1  g592(.A(KEYINPUT49), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT109), .ZN(new_n1019));
  XNOR2_X1  g594(.A(new_n1018), .B(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT49), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(new_n978), .ZN(new_n1024));
  NOR3_X1   g599(.A1(new_n1023), .A2(new_n995), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n750), .A2(G1976), .ZN(new_n1026));
  OR2_X1    g601(.A1(new_n1026), .A2(KEYINPUT108), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(KEYINPUT108), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1024), .A2(new_n995), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1027), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  AOI22_X1  g605(.A1(new_n1020), .A2(new_n1025), .B1(new_n1030), .B2(KEYINPUT52), .ZN(new_n1031));
  INV_X1    g606(.A(G1976), .ZN(new_n1032));
  AOI21_X1  g607(.A(KEYINPUT52), .B1(G288), .B2(new_n1032), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n1027), .A2(new_n1028), .A3(new_n1029), .A4(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1031), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT107), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1009), .A2(new_n761), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1038), .B1(new_n969), .B2(G2090), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(G8), .ZN(new_n1040));
  NAND2_X1  g615(.A1(G303), .A2(G8), .ZN(new_n1041));
  XOR2_X1   g616(.A(new_n1041), .B(KEYINPUT55), .Z(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1037), .B1(new_n1040), .B2(new_n1043), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1039), .A2(KEYINPUT107), .A3(G8), .A4(new_n1042), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n968), .A2(KEYINPUT50), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1047), .B(new_n943), .C1(KEYINPUT50), .C2(new_n940), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1038), .B1(new_n1048), .B2(G2090), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT110), .ZN(new_n1050));
  AND2_X1   g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(G8), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1043), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1036), .A2(new_n1046), .A3(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT121), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1036), .A2(new_n1053), .A3(KEYINPUT121), .A4(new_n1046), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1015), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  AND3_X1   g633(.A1(new_n1008), .A2(KEYINPUT122), .A3(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT122), .B1(new_n1008), .B2(new_n1058), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1002), .B1(new_n1001), .B2(new_n1007), .ZN(new_n1061));
  NOR3_X1   g636(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT114), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1040), .A2(new_n1043), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1063), .B1(new_n1035), .B2(new_n1065), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1031), .A2(new_n1064), .A3(KEYINPUT114), .A4(new_n1034), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(KEYINPUT63), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1005), .A2(G286), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(new_n1046), .ZN(new_n1071));
  OAI21_X1  g646(.A(KEYINPUT115), .B1(new_n1069), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT63), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1070), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1073), .B1(new_n1054), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1071), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT115), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1076), .A2(new_n1077), .A3(KEYINPUT63), .A4(new_n1068), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1072), .A2(new_n1075), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1046), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1020), .A2(new_n1025), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(new_n1032), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1016), .B1(new_n1082), .B2(G288), .ZN(new_n1083));
  AOI22_X1  g658(.A1(new_n1080), .A2(new_n1036), .B1(new_n1083), .B2(new_n1029), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1001), .A2(new_n1007), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n969), .A2(new_n716), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1024), .A2(new_n732), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n596), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n569), .A2(KEYINPUT57), .ZN(new_n1090));
  AOI22_X1  g665(.A1(G299), .A2(KEYINPUT57), .B1(new_n564), .B2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1048), .A2(new_n742), .ZN(new_n1093));
  XOR2_X1   g668(.A(KEYINPUT56), .B(G2072), .Z(new_n1094));
  OR2_X1    g669(.A1(new_n1009), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1089), .B1(new_n1092), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1092), .A2(new_n1096), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1096), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(new_n1091), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1098), .A2(KEYINPUT61), .A3(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT61), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1099), .A2(new_n1102), .A3(new_n1091), .ZN(new_n1103));
  XOR2_X1   g678(.A(KEYINPUT116), .B(G1341), .Z(new_n1104));
  XNOR2_X1  g679(.A(new_n1104), .B(KEYINPUT58), .ZN(new_n1105));
  OAI22_X1  g680(.A1(new_n1009), .A2(G1996), .B1(new_n1024), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(new_n548), .ZN(new_n1107));
  XNOR2_X1  g682(.A(new_n1107), .B(KEYINPUT59), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1109), .A2(new_n597), .ZN(new_n1110));
  OAI21_X1  g685(.A(KEYINPUT60), .B1(new_n1110), .B2(new_n1089), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1101), .A2(new_n1103), .A3(new_n1108), .A4(new_n1111), .ZN(new_n1112));
  NOR3_X1   g687(.A1(new_n1109), .A2(KEYINPUT60), .A3(new_n596), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1097), .B(new_n1098), .C1(new_n1112), .C2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1012), .B1(new_n1011), .B2(new_n1010), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(G171), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n1116), .B(KEYINPUT54), .C1(G171), .C2(new_n1014), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1085), .A2(new_n1086), .A3(new_n1114), .A4(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1015), .B1(G171), .B2(new_n1115), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT54), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  XNOR2_X1  g696(.A(new_n1121), .B(KEYINPUT120), .ZN(new_n1122));
  OAI211_X1 g697(.A(new_n1079), .B(new_n1084), .C1(new_n1118), .C2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n959), .B1(new_n1062), .B2(new_n1123), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n726), .A2(G2067), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n850), .A2(new_n781), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1125), .B1(new_n955), .B2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1127), .A2(new_n949), .ZN(new_n1128));
  XOR2_X1   g703(.A(new_n1128), .B(KEYINPUT123), .Z(new_n1129));
  AOI21_X1  g704(.A(new_n949), .B1(new_n952), .B2(new_n953), .ZN(new_n1130));
  XOR2_X1   g705(.A(new_n947), .B(KEYINPUT46), .Z(new_n1131));
  NOR2_X1   g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  XNOR2_X1  g707(.A(new_n1132), .B(KEYINPUT47), .ZN(new_n1133));
  NOR2_X1   g708(.A1(G290), .A2(G1986), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n945), .A2(new_n1134), .ZN(new_n1135));
  XNOR2_X1  g710(.A(new_n1135), .B(KEYINPUT124), .ZN(new_n1136));
  XOR2_X1   g711(.A(new_n1136), .B(KEYINPUT48), .Z(new_n1137));
  NOR2_X1   g712(.A1(new_n1137), .A2(new_n957), .ZN(new_n1138));
  NOR3_X1   g713(.A1(new_n1129), .A2(new_n1133), .A3(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1124), .A2(new_n1139), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g715(.A(KEYINPUT127), .ZN(new_n1142));
  AOI21_X1  g716(.A(G229), .B1(new_n925), .B2(new_n933), .ZN(new_n1143));
  NAND3_X1  g717(.A1(new_n637), .A2(new_n458), .A3(new_n653), .ZN(new_n1144));
  XNOR2_X1  g718(.A(new_n1144), .B(KEYINPUT125), .ZN(new_n1145));
  AOI21_X1  g719(.A(new_n1145), .B1(new_n870), .B2(new_n871), .ZN(new_n1146));
  INV_X1    g720(.A(KEYINPUT126), .ZN(new_n1147));
  AND3_X1   g721(.A1(new_n1143), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  AOI21_X1  g722(.A(new_n1147), .B1(new_n1143), .B2(new_n1146), .ZN(new_n1149));
  OAI21_X1  g723(.A(new_n1142), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g724(.A1(new_n1143), .A2(new_n1146), .ZN(new_n1151));
  NAND2_X1  g725(.A1(new_n1151), .A2(KEYINPUT126), .ZN(new_n1152));
  NAND3_X1  g726(.A1(new_n1143), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1153));
  NAND3_X1  g727(.A1(new_n1152), .A2(KEYINPUT127), .A3(new_n1153), .ZN(new_n1154));
  NAND2_X1  g728(.A1(new_n1150), .A2(new_n1154), .ZN(G308));
  NAND2_X1  g729(.A1(new_n1152), .A2(new_n1153), .ZN(G225));
endmodule


