

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765;

  BUF_X1 U380 ( .A(n582), .Z(n599) );
  INV_X1 U381 ( .A(G953), .ZN(n759) );
  NOR2_X1 U382 ( .A1(n586), .A2(n687), .ZN(n568) );
  NOR2_X2 U383 ( .A1(n619), .A2(n567), .ZN(n753) );
  XNOR2_X2 U384 ( .A(n379), .B(KEYINPUT48), .ZN(n619) );
  XNOR2_X2 U385 ( .A(n412), .B(n509), .ZN(n459) );
  XNOR2_X2 U386 ( .A(n477), .B(n498), .ZN(n412) );
  XNOR2_X1 U387 ( .A(n578), .B(KEYINPUT35), .ZN(n765) );
  OR2_X1 U388 ( .A1(n554), .A2(n553), .ZN(n555) );
  NOR2_X1 U389 ( .A1(n577), .A2(n576), .ZN(n578) );
  NAND2_X1 U390 ( .A1(n396), .A2(n395), .ZN(n560) );
  AND2_X1 U391 ( .A1(n393), .A2(n398), .ZN(n396) );
  NOR2_X1 U392 ( .A1(n690), .A2(n688), .ZN(n594) );
  AND2_X1 U393 ( .A1(n528), .A2(n517), .ZN(n519) );
  XNOR2_X1 U394 ( .A(n530), .B(n529), .ZN(n585) );
  OR2_X1 U395 ( .A1(n739), .A2(G902), .ZN(n404) );
  NOR2_X1 U396 ( .A1(G953), .A2(G237), .ZN(n497) );
  XNOR2_X1 U397 ( .A(n383), .B(n527), .ZN(n382) );
  NAND2_X1 U398 ( .A1(n650), .A2(n636), .ZN(n383) );
  NOR2_X1 U399 ( .A1(n726), .A2(n718), .ZN(n723) );
  XNOR2_X2 U400 ( .A(n755), .B(n417), .ZN(n729) );
  NOR2_X1 U401 ( .A1(n619), .A2(n392), .ZN(n391) );
  OR2_X1 U402 ( .A1(n567), .A2(n610), .ZN(n392) );
  INV_X1 U403 ( .A(n491), .ZN(n401) );
  XNOR2_X1 U404 ( .A(G119), .B(G113), .ZN(n455) );
  XNOR2_X1 U405 ( .A(G146), .B(G125), .ZN(n475) );
  NAND2_X1 U406 ( .A1(n382), .A2(n380), .ZN(n379) );
  XNOR2_X1 U407 ( .A(n381), .B(KEYINPUT73), .ZN(n380) );
  OR2_X1 U408 ( .A1(n678), .A2(n400), .ZN(n399) );
  INV_X1 U409 ( .A(n538), .ZN(n683) );
  XNOR2_X1 U410 ( .A(n413), .B(G137), .ZN(n421) );
  INV_X1 U411 ( .A(G140), .ZN(n413) );
  XNOR2_X1 U412 ( .A(G119), .B(G128), .ZN(n422) );
  XNOR2_X1 U413 ( .A(G110), .B(KEYINPUT95), .ZN(n423) );
  XOR2_X1 U414 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n424) );
  XNOR2_X1 U415 ( .A(n407), .B(n406), .ZN(n405) );
  XNOR2_X1 U416 ( .A(G107), .B(KEYINPUT81), .ZN(n406) );
  XNOR2_X1 U417 ( .A(n408), .B(G146), .ZN(n407) );
  INV_X1 U418 ( .A(G101), .ZN(n408) );
  NAND2_X1 U419 ( .A1(n371), .A2(n368), .ZN(n710) );
  AND2_X1 U420 ( .A1(n373), .A2(n372), .ZN(n371) );
  NAND2_X1 U421 ( .A1(n370), .A2(n369), .ZN(n368) );
  NAND2_X1 U422 ( .A1(n585), .A2(KEYINPUT33), .ZN(n372) );
  INV_X1 U423 ( .A(n364), .ZN(n537) );
  XNOR2_X1 U424 ( .A(n430), .B(n358), .ZN(n403) );
  XOR2_X1 U425 ( .A(G104), .B(G122), .Z(n493) );
  XNOR2_X1 U426 ( .A(G113), .B(G143), .ZN(n492) );
  XOR2_X1 U427 ( .A(KEYINPUT64), .B(KEYINPUT46), .Z(n527) );
  XNOR2_X1 U428 ( .A(KEYINPUT15), .B(G902), .ZN(n610) );
  XNOR2_X1 U429 ( .A(G137), .B(G146), .ZN(n451) );
  XOR2_X1 U430 ( .A(G116), .B(KEYINPUT5), .Z(n449) );
  XNOR2_X1 U431 ( .A(n608), .B(n390), .ZN(n389) );
  INV_X1 U432 ( .A(KEYINPUT88), .ZN(n390) );
  XNOR2_X1 U433 ( .A(G143), .B(G128), .ZN(n470) );
  NAND2_X1 U434 ( .A1(G234), .A2(G237), .ZN(n437) );
  NOR2_X1 U435 ( .A1(n687), .A2(n516), .ZN(n528) );
  INV_X1 U436 ( .A(n597), .ZN(n370) );
  NOR2_X1 U437 ( .A1(n585), .A2(KEYINPUT33), .ZN(n369) );
  NAND2_X1 U438 ( .A1(n597), .A2(KEYINPUT33), .ZN(n373) );
  NAND2_X1 U439 ( .A1(n569), .A2(n568), .ZN(n597) );
  XNOR2_X1 U440 ( .A(n539), .B(KEYINPUT19), .ZN(n540) );
  NAND2_X1 U441 ( .A1(n364), .A2(n683), .ZN(n539) );
  XNOR2_X1 U442 ( .A(n461), .B(n641), .ZN(n530) );
  XNOR2_X1 U443 ( .A(G101), .B(KEYINPUT74), .ZN(n454) );
  XNOR2_X1 U444 ( .A(G122), .B(G116), .ZN(n480) );
  XNOR2_X1 U445 ( .A(KEYINPUT18), .B(KEYINPUT82), .ZN(n474) );
  NAND2_X1 U446 ( .A1(n623), .A2(n672), .ZN(n726) );
  XNOR2_X1 U447 ( .A(n384), .B(KEYINPUT66), .ZN(n623) );
  NAND2_X1 U448 ( .A1(n385), .A2(n363), .ZN(n384) );
  NAND2_X1 U449 ( .A1(n394), .A2(n401), .ZN(n395) );
  BUF_X1 U450 ( .A(n530), .Z(n693) );
  INV_X1 U451 ( .A(KEYINPUT98), .ZN(n434) );
  XNOR2_X1 U452 ( .A(n427), .B(n426), .ZN(n739) );
  XNOR2_X1 U453 ( .A(n405), .B(n415), .ZN(n416) );
  AND2_X1 U454 ( .A1(n630), .A2(G953), .ZN(n741) );
  BUF_X1 U455 ( .A(n759), .Z(n375) );
  XNOR2_X1 U456 ( .A(n526), .B(KEYINPUT42), .ZN(n636) );
  AND2_X1 U457 ( .A1(n536), .A2(n690), .ZN(n669) );
  NOR2_X1 U458 ( .A1(n563), .A2(n537), .ZN(n535) );
  XNOR2_X1 U459 ( .A(n374), .B(KEYINPUT34), .ZN(n577) );
  NAND2_X1 U460 ( .A1(n710), .A2(n599), .ZN(n374) );
  XOR2_X1 U461 ( .A(n428), .B(KEYINPUT25), .Z(n358) );
  XOR2_X1 U462 ( .A(n424), .B(n423), .Z(n359) );
  NOR2_X1 U463 ( .A1(n678), .A2(n397), .ZN(n360) );
  AND2_X1 U464 ( .A1(n402), .A2(n467), .ZN(n361) );
  NAND2_X1 U465 ( .A1(n573), .A2(n572), .ZN(n362) );
  XOR2_X1 U466 ( .A(n612), .B(KEYINPUT69), .Z(n363) );
  XNOR2_X2 U467 ( .A(n488), .B(n365), .ZN(n364) );
  XOR2_X1 U468 ( .A(n487), .B(KEYINPUT92), .Z(n365) );
  NAND2_X1 U469 ( .A1(n366), .A2(n568), .ZN(n435) );
  XNOR2_X1 U470 ( .A(n366), .B(KEYINPUT1), .ZN(n569) );
  AND2_X1 U471 ( .A1(n520), .A2(n366), .ZN(n541) );
  XNOR2_X2 U472 ( .A(n418), .B(G469), .ZN(n366) );
  XNOR2_X2 U473 ( .A(n514), .B(KEYINPUT40), .ZN(n650) );
  OR2_X2 U474 ( .A1(n483), .A2(n743), .ZN(n484) );
  NAND2_X1 U475 ( .A1(n753), .A2(n367), .ZN(n673) );
  NAND2_X1 U476 ( .A1(n391), .A2(n367), .ZN(n385) );
  NAND2_X1 U477 ( .A1(n367), .A2(n618), .ZN(n620) );
  NAND2_X1 U478 ( .A1(n367), .A2(n375), .ZN(n746) );
  XNOR2_X2 U479 ( .A(n376), .B(KEYINPUT45), .ZN(n367) );
  XNOR2_X1 U480 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X2 U481 ( .A(n522), .B(n521), .ZN(n677) );
  NAND2_X1 U482 ( .A1(n721), .A2(n610), .ZN(n488) );
  NAND2_X1 U483 ( .A1(n484), .A2(n485), .ZN(n721) );
  NAND2_X1 U484 ( .A1(n377), .A2(n388), .ZN(n376) );
  XNOR2_X1 U485 ( .A(n378), .B(KEYINPUT87), .ZN(n377) );
  NAND2_X1 U486 ( .A1(n387), .A2(n386), .ZN(n378) );
  NAND2_X1 U487 ( .A1(n559), .A2(n638), .ZN(n381) );
  XNOR2_X1 U488 ( .A(n605), .B(KEYINPUT104), .ZN(n386) );
  NAND2_X1 U489 ( .A1(n592), .A2(KEYINPUT44), .ZN(n387) );
  NAND2_X1 U490 ( .A1(n609), .A2(n389), .ZN(n388) );
  NAND2_X1 U491 ( .A1(n540), .A2(n362), .ZN(n575) );
  NAND2_X1 U492 ( .A1(n402), .A2(n360), .ZN(n393) );
  XNOR2_X2 U493 ( .A(n447), .B(n446), .ZN(n402) );
  INV_X1 U494 ( .A(n402), .ZN(n394) );
  NAND2_X1 U495 ( .A1(n467), .A2(n491), .ZN(n397) );
  NAND2_X1 U496 ( .A1(n399), .A2(n401), .ZN(n398) );
  INV_X1 U497 ( .A(n467), .ZN(n400) );
  XNOR2_X2 U498 ( .A(n404), .B(n403), .ZN(n586) );
  XNOR2_X2 U499 ( .A(KEYINPUT91), .B(KEYINPUT17), .ZN(n468) );
  XNOR2_X2 U500 ( .A(n410), .B(KEYINPUT4), .ZN(n477) );
  XNOR2_X1 U501 ( .A(n498), .B(n409), .ZN(n499) );
  AND2_X1 U502 ( .A1(G214), .A2(n497), .ZN(n409) );
  INV_X1 U503 ( .A(KEYINPUT79), .ZN(n450) );
  XNOR2_X1 U504 ( .A(n451), .B(n450), .ZN(n452) );
  NOR2_X1 U505 ( .A1(n531), .A2(n585), .ZN(n532) );
  XNOR2_X1 U506 ( .A(n453), .B(n452), .ZN(n458) );
  INV_X1 U507 ( .A(KEYINPUT80), .ZN(n446) );
  INV_X1 U508 ( .A(n421), .ZN(n414) );
  XNOR2_X1 U509 ( .A(n420), .B(n754), .ZN(n427) );
  BUF_X1 U510 ( .A(n569), .Z(n690) );
  XNOR2_X1 U511 ( .A(n584), .B(n583), .ZN(n591) );
  INV_X1 U512 ( .A(KEYINPUT60), .ZN(n633) );
  XNOR2_X2 U513 ( .A(KEYINPUT65), .B(KEYINPUT70), .ZN(n410) );
  XNOR2_X2 U514 ( .A(KEYINPUT71), .B(KEYINPUT72), .ZN(n411) );
  XNOR2_X2 U515 ( .A(n411), .B(G131), .ZN(n498) );
  XNOR2_X1 U516 ( .A(n470), .B(G134), .ZN(n509) );
  XNOR2_X2 U517 ( .A(n459), .B(n414), .ZN(n755) );
  XNOR2_X1 U518 ( .A(G110), .B(G104), .ZN(n742) );
  XNOR2_X1 U519 ( .A(n742), .B(KEYINPUT75), .ZN(n472) );
  NAND2_X1 U520 ( .A1(G227), .A2(n375), .ZN(n415) );
  XNOR2_X1 U521 ( .A(n472), .B(n416), .ZN(n417) );
  OR2_X2 U522 ( .A1(n729), .A2(G902), .ZN(n418) );
  NAND2_X1 U523 ( .A1(G234), .A2(n759), .ZN(n419) );
  XOR2_X1 U524 ( .A(KEYINPUT8), .B(n419), .Z(n505) );
  NAND2_X1 U525 ( .A1(G221), .A2(n505), .ZN(n420) );
  XNOR2_X1 U526 ( .A(n475), .B(KEYINPUT10), .ZN(n754) );
  XNOR2_X1 U527 ( .A(n422), .B(n421), .ZN(n425) );
  XNOR2_X1 U528 ( .A(n425), .B(n359), .ZN(n426) );
  INV_X1 U529 ( .A(KEYINPUT96), .ZN(n428) );
  NAND2_X1 U530 ( .A1(n610), .A2(G234), .ZN(n429) );
  XNOR2_X1 U531 ( .A(n429), .B(KEYINPUT20), .ZN(n431) );
  NAND2_X1 U532 ( .A1(G217), .A2(n431), .ZN(n430) );
  NAND2_X1 U533 ( .A1(n431), .A2(G221), .ZN(n433) );
  XOR2_X1 U534 ( .A(KEYINPUT21), .B(KEYINPUT97), .Z(n432) );
  XNOR2_X1 U535 ( .A(n433), .B(n432), .ZN(n687) );
  XNOR2_X2 U536 ( .A(n435), .B(n434), .ZN(n600) );
  INV_X1 U537 ( .A(KEYINPUT107), .ZN(n436) );
  XNOR2_X1 U538 ( .A(n600), .B(n436), .ZN(n445) );
  XNOR2_X1 U539 ( .A(KEYINPUT14), .B(n437), .ZN(n440) );
  NAND2_X1 U540 ( .A1(G952), .A2(n440), .ZN(n708) );
  NOR2_X1 U541 ( .A1(G953), .A2(n708), .ZN(n439) );
  INV_X1 U542 ( .A(KEYINPUT94), .ZN(n438) );
  XNOR2_X1 U543 ( .A(n439), .B(n438), .ZN(n573) );
  NAND2_X1 U544 ( .A1(G902), .A2(n440), .ZN(n570) );
  NOR2_X1 U545 ( .A1(G900), .A2(n570), .ZN(n441) );
  NAND2_X1 U546 ( .A1(G953), .A2(n441), .ZN(n443) );
  INV_X1 U547 ( .A(KEYINPUT105), .ZN(n442) );
  XNOR2_X1 U548 ( .A(n443), .B(n442), .ZN(n444) );
  NAND2_X1 U549 ( .A1(n573), .A2(n444), .ZN(n515) );
  NAND2_X1 U550 ( .A1(n445), .A2(n515), .ZN(n447) );
  NAND2_X1 U551 ( .A1(n497), .A2(G210), .ZN(n448) );
  XNOR2_X1 U552 ( .A(n449), .B(n448), .ZN(n453) );
  XNOR2_X1 U553 ( .A(n455), .B(n454), .ZN(n457) );
  XNOR2_X1 U554 ( .A(KEYINPUT90), .B(KEYINPUT3), .ZN(n456) );
  XNOR2_X1 U555 ( .A(n457), .B(n456), .ZN(n482) );
  XNOR2_X1 U556 ( .A(n458), .B(n482), .ZN(n460) );
  XNOR2_X1 U557 ( .A(n459), .B(n460), .ZN(n643) );
  INV_X1 U558 ( .A(G902), .ZN(n512) );
  NAND2_X1 U559 ( .A1(n643), .A2(n512), .ZN(n461) );
  INV_X1 U560 ( .A(G472), .ZN(n641) );
  NOR2_X1 U561 ( .A1(G237), .A2(G902), .ZN(n462) );
  XNOR2_X1 U562 ( .A(n462), .B(KEYINPUT78), .ZN(n486) );
  INV_X1 U563 ( .A(G214), .ZN(n463) );
  OR2_X1 U564 ( .A1(n486), .A2(n463), .ZN(n464) );
  XNOR2_X1 U565 ( .A(n464), .B(KEYINPUT93), .ZN(n538) );
  NOR2_X1 U566 ( .A1(n693), .A2(n538), .ZN(n466) );
  XNOR2_X1 U567 ( .A(KEYINPUT108), .B(KEYINPUT30), .ZN(n465) );
  XNOR2_X1 U568 ( .A(n466), .B(n465), .ZN(n467) );
  NAND2_X1 U569 ( .A1(n759), .A2(G224), .ZN(n469) );
  XNOR2_X1 U570 ( .A(n469), .B(n468), .ZN(n471) );
  XNOR2_X1 U571 ( .A(n471), .B(n470), .ZN(n473) );
  XNOR2_X1 U572 ( .A(n473), .B(n472), .ZN(n479) );
  XNOR2_X1 U573 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U574 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U575 ( .A(n479), .B(n478), .ZN(n483) );
  XNOR2_X1 U576 ( .A(n480), .B(G107), .ZN(n508) );
  XNOR2_X1 U577 ( .A(n508), .B(KEYINPUT16), .ZN(n481) );
  XNOR2_X1 U578 ( .A(n482), .B(n481), .ZN(n743) );
  NAND2_X1 U579 ( .A1(n483), .A2(n743), .ZN(n485) );
  INV_X1 U580 ( .A(G210), .ZN(n718) );
  OR2_X1 U581 ( .A1(n486), .A2(n718), .ZN(n487) );
  XNOR2_X1 U582 ( .A(KEYINPUT77), .B(KEYINPUT38), .ZN(n489) );
  XNOR2_X1 U583 ( .A(n537), .B(n489), .ZN(n678) );
  XOR2_X1 U584 ( .A(KEYINPUT86), .B(KEYINPUT39), .Z(n490) );
  XNOR2_X1 U585 ( .A(n490), .B(KEYINPUT76), .ZN(n491) );
  XNOR2_X1 U586 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U587 ( .A(n754), .B(n494), .ZN(n502) );
  XOR2_X1 U588 ( .A(G140), .B(KEYINPUT12), .Z(n496) );
  XNOR2_X1 U589 ( .A(KEYINPUT11), .B(KEYINPUT99), .ZN(n495) );
  XNOR2_X1 U590 ( .A(n496), .B(n495), .ZN(n500) );
  XNOR2_X1 U591 ( .A(n502), .B(n501), .ZN(n625) );
  NOR2_X1 U592 ( .A1(G902), .A2(n625), .ZN(n504) );
  XNOR2_X1 U593 ( .A(KEYINPUT13), .B(G475), .ZN(n503) );
  XNOR2_X1 U594 ( .A(n504), .B(n503), .ZN(n557) );
  XOR2_X1 U595 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n507) );
  NAND2_X1 U596 ( .A1(G217), .A2(n505), .ZN(n506) );
  XNOR2_X1 U597 ( .A(n507), .B(n506), .ZN(n511) );
  XNOR2_X1 U598 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U599 ( .A(n511), .B(n510), .ZN(n733) );
  NAND2_X1 U600 ( .A1(n733), .A2(n512), .ZN(n513) );
  XNOR2_X1 U601 ( .A(n513), .B(G478), .ZN(n556) );
  INV_X1 U602 ( .A(n556), .ZN(n542) );
  NAND2_X1 U603 ( .A1(n557), .A2(n542), .ZN(n543) );
  INV_X1 U604 ( .A(n543), .ZN(n663) );
  NAND2_X1 U605 ( .A1(n560), .A2(n663), .ZN(n514) );
  NAND2_X1 U606 ( .A1(n515), .A2(n586), .ZN(n516) );
  INV_X1 U607 ( .A(n693), .ZN(n517) );
  XOR2_X1 U608 ( .A(KEYINPUT109), .B(KEYINPUT28), .Z(n518) );
  XNOR2_X1 U609 ( .A(n519), .B(n518), .ZN(n520) );
  OR2_X1 U610 ( .A1(n557), .A2(n556), .ZN(n522) );
  INV_X1 U611 ( .A(KEYINPUT100), .ZN(n521) );
  INV_X1 U612 ( .A(n678), .ZN(n523) );
  AND2_X1 U613 ( .A1(n677), .A2(n523), .ZN(n684) );
  NAND2_X1 U614 ( .A1(n684), .A2(n683), .ZN(n525) );
  XNOR2_X1 U615 ( .A(KEYINPUT110), .B(KEYINPUT41), .ZN(n524) );
  XNOR2_X1 U616 ( .A(n525), .B(n524), .ZN(n709) );
  NAND2_X1 U617 ( .A1(n541), .A2(n709), .ZN(n526) );
  INV_X1 U618 ( .A(n528), .ZN(n531) );
  INV_X1 U619 ( .A(KEYINPUT6), .ZN(n529) );
  XOR2_X1 U620 ( .A(KEYINPUT106), .B(n532), .Z(n533) );
  NOR2_X1 U621 ( .A1(n543), .A2(n533), .ZN(n534) );
  NAND2_X1 U622 ( .A1(n534), .A2(n683), .ZN(n563) );
  XNOR2_X1 U623 ( .A(n535), .B(KEYINPUT36), .ZN(n536) );
  NAND2_X1 U624 ( .A1(n541), .A2(n540), .ZN(n550) );
  OR2_X1 U625 ( .A1(n542), .A2(n557), .ZN(n561) );
  NAND2_X1 U626 ( .A1(n543), .A2(n561), .ZN(n547) );
  INV_X1 U627 ( .A(n547), .ZN(n679) );
  NOR2_X1 U628 ( .A1(n550), .A2(n679), .ZN(n544) );
  NOR2_X1 U629 ( .A1(KEYINPUT85), .A2(n544), .ZN(n545) );
  NOR2_X1 U630 ( .A1(KEYINPUT47), .A2(n545), .ZN(n554) );
  INV_X1 U631 ( .A(KEYINPUT85), .ZN(n546) );
  NAND2_X1 U632 ( .A1(n550), .A2(n546), .ZN(n548) );
  NAND2_X1 U633 ( .A1(n548), .A2(n547), .ZN(n549) );
  NAND2_X1 U634 ( .A1(n549), .A2(KEYINPUT47), .ZN(n552) );
  INV_X1 U635 ( .A(n550), .ZN(n660) );
  NAND2_X1 U636 ( .A1(n660), .A2(KEYINPUT85), .ZN(n551) );
  NAND2_X1 U637 ( .A1(n552), .A2(n551), .ZN(n553) );
  NOR2_X1 U638 ( .A1(n669), .A2(n555), .ZN(n559) );
  NAND2_X1 U639 ( .A1(n557), .A2(n556), .ZN(n576) );
  NOR2_X1 U640 ( .A1(n576), .A2(n537), .ZN(n558) );
  NAND2_X1 U641 ( .A1(n361), .A2(n558), .ZN(n638) );
  INV_X1 U642 ( .A(n561), .ZN(n665) );
  NAND2_X1 U643 ( .A1(n560), .A2(n665), .ZN(n562) );
  XNOR2_X1 U644 ( .A(n562), .B(KEYINPUT111), .ZN(n764) );
  INV_X1 U645 ( .A(n764), .ZN(n566) );
  OR2_X1 U646 ( .A1(n563), .A2(n690), .ZN(n564) );
  XNOR2_X1 U647 ( .A(n564), .B(KEYINPUT43), .ZN(n565) );
  NAND2_X1 U648 ( .A1(n565), .A2(n537), .ZN(n649) );
  NAND2_X1 U649 ( .A1(n566), .A2(n649), .ZN(n567) );
  INV_X1 U650 ( .A(n570), .ZN(n571) );
  NOR2_X1 U651 ( .A1(G898), .A2(n375), .ZN(n744) );
  NAND2_X1 U652 ( .A1(n571), .A2(n744), .ZN(n572) );
  INV_X1 U653 ( .A(KEYINPUT0), .ZN(n574) );
  XNOR2_X2 U654 ( .A(n575), .B(n574), .ZN(n582) );
  INV_X1 U655 ( .A(n687), .ZN(n579) );
  NAND2_X1 U656 ( .A1(n677), .A2(n579), .ZN(n580) );
  XNOR2_X1 U657 ( .A(n580), .B(KEYINPUT101), .ZN(n581) );
  NAND2_X1 U658 ( .A1(n582), .A2(n581), .ZN(n584) );
  XNOR2_X1 U659 ( .A(KEYINPUT67), .B(KEYINPUT22), .ZN(n583) );
  NAND2_X1 U660 ( .A1(n591), .A2(n585), .ZN(n593) );
  XNOR2_X1 U661 ( .A(n586), .B(KEYINPUT102), .ZN(n688) );
  NAND2_X1 U662 ( .A1(n690), .A2(n688), .ZN(n587) );
  NOR2_X1 U663 ( .A1(n593), .A2(n587), .ZN(n588) );
  XNOR2_X1 U664 ( .A(n588), .B(KEYINPUT32), .ZN(n640) );
  NAND2_X1 U665 ( .A1(n693), .A2(n586), .ZN(n589) );
  NOR2_X1 U666 ( .A1(n690), .A2(n589), .ZN(n590) );
  AND2_X1 U667 ( .A1(n591), .A2(n590), .ZN(n635) );
  NOR2_X1 U668 ( .A1(n640), .A2(n635), .ZN(n607) );
  NAND2_X1 U669 ( .A1(n765), .A2(n607), .ZN(n592) );
  INV_X1 U670 ( .A(n593), .ZN(n595) );
  NAND2_X1 U671 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X2 U672 ( .A(n596), .B(KEYINPUT103), .ZN(n639) );
  NOR2_X1 U673 ( .A1(n597), .A2(n693), .ZN(n697) );
  NAND2_X1 U674 ( .A1(n697), .A2(n599), .ZN(n598) );
  XNOR2_X1 U675 ( .A(n598), .B(KEYINPUT31), .ZN(n666) );
  INV_X1 U676 ( .A(n599), .ZN(n602) );
  NAND2_X1 U677 ( .A1(n600), .A2(n693), .ZN(n601) );
  NOR2_X1 U678 ( .A1(n602), .A2(n601), .ZN(n653) );
  NOR2_X1 U679 ( .A1(n666), .A2(n653), .ZN(n603) );
  NOR2_X1 U680 ( .A1(n603), .A2(n679), .ZN(n604) );
  NOR2_X2 U681 ( .A1(n639), .A2(n604), .ZN(n605) );
  INV_X1 U682 ( .A(n765), .ZN(n606) );
  NOR2_X1 U683 ( .A1(n606), .A2(KEYINPUT44), .ZN(n609) );
  INV_X1 U684 ( .A(n607), .ZN(n608) );
  INV_X1 U685 ( .A(n610), .ZN(n611) );
  NAND2_X1 U686 ( .A1(n611), .A2(KEYINPUT2), .ZN(n612) );
  INV_X1 U687 ( .A(KEYINPUT83), .ZN(n613) );
  NAND2_X1 U688 ( .A1(n613), .A2(KEYINPUT2), .ZN(n614) );
  NOR2_X1 U689 ( .A1(n673), .A2(n614), .ZN(n622) );
  INV_X1 U690 ( .A(KEYINPUT2), .ZN(n615) );
  NOR2_X1 U691 ( .A1(n764), .A2(n615), .ZN(n617) );
  NAND2_X1 U692 ( .A1(n649), .A2(KEYINPUT83), .ZN(n616) );
  NOR2_X1 U693 ( .A1(n617), .A2(n616), .ZN(n618) );
  NOR2_X1 U694 ( .A1(n620), .A2(n619), .ZN(n621) );
  NOR2_X1 U695 ( .A1(n622), .A2(n621), .ZN(n672) );
  INV_X1 U696 ( .A(n726), .ZN(n624) );
  NAND2_X1 U697 ( .A1(n624), .A2(G475), .ZN(n629) );
  XOR2_X1 U698 ( .A(KEYINPUT89), .B(KEYINPUT68), .Z(n627) );
  XNOR2_X1 U699 ( .A(n625), .B(KEYINPUT59), .ZN(n626) );
  XNOR2_X1 U700 ( .A(n627), .B(n626), .ZN(n628) );
  XNOR2_X1 U701 ( .A(n629), .B(n628), .ZN(n632) );
  INV_X1 U702 ( .A(G952), .ZN(n630) );
  INV_X1 U703 ( .A(n741), .ZN(n631) );
  NAND2_X1 U704 ( .A1(n632), .A2(n631), .ZN(n634) );
  XNOR2_X1 U705 ( .A(n634), .B(n633), .ZN(G60) );
  XOR2_X1 U706 ( .A(G110), .B(n635), .Z(G12) );
  XNOR2_X1 U707 ( .A(G137), .B(KEYINPUT127), .ZN(n637) );
  XOR2_X1 U708 ( .A(n637), .B(n636), .Z(G39) );
  XNOR2_X1 U709 ( .A(n638), .B(G143), .ZN(G45) );
  XOR2_X1 U710 ( .A(n639), .B(G101), .Z(G3) );
  XOR2_X1 U711 ( .A(n640), .B(G119), .Z(G21) );
  NOR2_X1 U712 ( .A1(n726), .A2(n641), .ZN(n645) );
  XNOR2_X1 U713 ( .A(KEYINPUT112), .B(KEYINPUT62), .ZN(n642) );
  XNOR2_X1 U714 ( .A(n643), .B(n642), .ZN(n644) );
  XNOR2_X1 U715 ( .A(n645), .B(n644), .ZN(n646) );
  NOR2_X1 U716 ( .A1(n646), .A2(n741), .ZN(n648) );
  XNOR2_X1 U717 ( .A(KEYINPUT113), .B(KEYINPUT63), .ZN(n647) );
  XNOR2_X1 U718 ( .A(n648), .B(n647), .ZN(G57) );
  XNOR2_X1 U719 ( .A(n649), .B(G140), .ZN(G42) );
  XNOR2_X1 U720 ( .A(n650), .B(G131), .ZN(G33) );
  NAND2_X1 U721 ( .A1(n653), .A2(n663), .ZN(n651) );
  XNOR2_X1 U722 ( .A(n651), .B(KEYINPUT114), .ZN(n652) );
  XNOR2_X1 U723 ( .A(G104), .B(n652), .ZN(G6) );
  XOR2_X1 U724 ( .A(KEYINPUT26), .B(KEYINPUT115), .Z(n655) );
  NAND2_X1 U725 ( .A1(n653), .A2(n665), .ZN(n654) );
  XNOR2_X1 U726 ( .A(n655), .B(n654), .ZN(n657) );
  XOR2_X1 U727 ( .A(G107), .B(KEYINPUT27), .Z(n656) );
  XNOR2_X1 U728 ( .A(n657), .B(n656), .ZN(G9) );
  XOR2_X1 U729 ( .A(G128), .B(KEYINPUT29), .Z(n659) );
  NAND2_X1 U730 ( .A1(n660), .A2(n665), .ZN(n658) );
  XNOR2_X1 U731 ( .A(n659), .B(n658), .ZN(G30) );
  NAND2_X1 U732 ( .A1(n660), .A2(n663), .ZN(n661) );
  XNOR2_X1 U733 ( .A(n661), .B(KEYINPUT116), .ZN(n662) );
  XNOR2_X1 U734 ( .A(G146), .B(n662), .ZN(G48) );
  NAND2_X1 U735 ( .A1(n666), .A2(n663), .ZN(n664) );
  XNOR2_X1 U736 ( .A(n664), .B(G113), .ZN(G15) );
  XOR2_X1 U737 ( .A(G116), .B(KEYINPUT117), .Z(n668) );
  NAND2_X1 U738 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U739 ( .A(n668), .B(n667), .ZN(G18) );
  XNOR2_X1 U740 ( .A(n669), .B(KEYINPUT37), .ZN(n670) );
  XNOR2_X1 U741 ( .A(n670), .B(KEYINPUT118), .ZN(n671) );
  XNOR2_X1 U742 ( .A(G125), .B(n671), .ZN(G27) );
  INV_X1 U743 ( .A(n672), .ZN(n676) );
  INV_X1 U744 ( .A(n673), .ZN(n674) );
  NOR2_X1 U745 ( .A1(n674), .A2(KEYINPUT2), .ZN(n675) );
  NOR2_X1 U746 ( .A1(n676), .A2(n675), .ZN(n716) );
  XOR2_X1 U747 ( .A(KEYINPUT121), .B(KEYINPUT52), .Z(n706) );
  INV_X1 U748 ( .A(n677), .ZN(n681) );
  OR2_X1 U749 ( .A1(n679), .A2(n678), .ZN(n680) );
  NAND2_X1 U750 ( .A1(n681), .A2(n680), .ZN(n682) );
  NAND2_X1 U751 ( .A1(n710), .A2(n682), .ZN(n686) );
  NOR2_X1 U752 ( .A1(n684), .A2(n683), .ZN(n685) );
  OR2_X1 U753 ( .A1(n686), .A2(n685), .ZN(n704) );
  NAND2_X1 U754 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U755 ( .A(n689), .B(KEYINPUT49), .ZN(n695) );
  NOR2_X1 U756 ( .A1(n690), .A2(n568), .ZN(n691) );
  XOR2_X1 U757 ( .A(KEYINPUT50), .B(n691), .Z(n692) );
  NAND2_X1 U758 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U759 ( .A1(n695), .A2(n694), .ZN(n696) );
  NOR2_X1 U760 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U761 ( .A(n698), .B(KEYINPUT119), .ZN(n699) );
  XNOR2_X1 U762 ( .A(KEYINPUT51), .B(n699), .ZN(n701) );
  INV_X1 U763 ( .A(n709), .ZN(n700) );
  NOR2_X1 U764 ( .A1(n701), .A2(n700), .ZN(n702) );
  XOR2_X1 U765 ( .A(KEYINPUT120), .B(n702), .Z(n703) );
  NAND2_X1 U766 ( .A1(n704), .A2(n703), .ZN(n705) );
  XOR2_X1 U767 ( .A(n706), .B(n705), .Z(n707) );
  NOR2_X1 U768 ( .A1(n708), .A2(n707), .ZN(n712) );
  AND2_X1 U769 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U770 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U771 ( .A(n713), .B(KEYINPUT122), .ZN(n714) );
  NAND2_X1 U772 ( .A1(n714), .A2(n375), .ZN(n715) );
  NOR2_X1 U773 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U774 ( .A(KEYINPUT53), .B(n717), .ZN(G75) );
  XNOR2_X1 U775 ( .A(KEYINPUT55), .B(KEYINPUT54), .ZN(n719) );
  XOR2_X1 U776 ( .A(n719), .B(KEYINPUT84), .Z(n720) );
  XNOR2_X1 U777 ( .A(n721), .B(n720), .ZN(n722) );
  XNOR2_X1 U778 ( .A(n723), .B(n722), .ZN(n724) );
  NOR2_X1 U779 ( .A1(n741), .A2(n724), .ZN(n725) );
  XNOR2_X1 U780 ( .A(KEYINPUT56), .B(n725), .ZN(G51) );
  INV_X1 U781 ( .A(n726), .ZN(n737) );
  NAND2_X1 U782 ( .A1(n737), .A2(G469), .ZN(n731) );
  XOR2_X1 U783 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n727) );
  XOR2_X1 U784 ( .A(n727), .B(KEYINPUT123), .Z(n728) );
  XNOR2_X1 U785 ( .A(n729), .B(n728), .ZN(n730) );
  XNOR2_X1 U786 ( .A(n731), .B(n730), .ZN(n732) );
  NOR2_X1 U787 ( .A1(n741), .A2(n732), .ZN(G54) );
  NAND2_X1 U788 ( .A1(n737), .A2(G478), .ZN(n735) );
  XOR2_X1 U789 ( .A(KEYINPUT124), .B(n733), .Z(n734) );
  XNOR2_X1 U790 ( .A(n735), .B(n734), .ZN(n736) );
  NOR2_X1 U791 ( .A1(n741), .A2(n736), .ZN(G63) );
  NAND2_X1 U792 ( .A1(n737), .A2(G217), .ZN(n738) );
  XNOR2_X1 U793 ( .A(n739), .B(n738), .ZN(n740) );
  NOR2_X1 U794 ( .A1(n741), .A2(n740), .ZN(G66) );
  XNOR2_X1 U795 ( .A(n743), .B(n742), .ZN(n745) );
  NOR2_X1 U796 ( .A1(n745), .A2(n744), .ZN(n752) );
  XOR2_X1 U797 ( .A(KEYINPUT125), .B(n746), .Z(n750) );
  NAND2_X1 U798 ( .A1(G953), .A2(G224), .ZN(n747) );
  XNOR2_X1 U799 ( .A(KEYINPUT61), .B(n747), .ZN(n748) );
  NAND2_X1 U800 ( .A1(n748), .A2(G898), .ZN(n749) );
  NAND2_X1 U801 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U802 ( .A(n752), .B(n751), .ZN(G69) );
  XNOR2_X1 U803 ( .A(n755), .B(n754), .ZN(n757) );
  XNOR2_X1 U804 ( .A(n753), .B(n757), .ZN(n756) );
  NOR2_X1 U805 ( .A1(n756), .A2(G953), .ZN(n762) );
  XOR2_X1 U806 ( .A(G227), .B(n757), .Z(n758) );
  NAND2_X1 U807 ( .A1(n758), .A2(G900), .ZN(n760) );
  NOR2_X1 U808 ( .A1(n760), .A2(n375), .ZN(n761) );
  NOR2_X1 U809 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U810 ( .A(KEYINPUT126), .B(n763), .ZN(G72) );
  XOR2_X1 U811 ( .A(G134), .B(n764), .Z(G36) );
  XNOR2_X1 U812 ( .A(n765), .B(G122), .ZN(G24) );
endmodule

