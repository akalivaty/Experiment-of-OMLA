//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 0 0 1 0 1 1 0 0 1 0 1 1 0 0 0 0 1 0 0 0 0 0 0 0 0 1 1 0 0 0 0 1 1 1 1 0 0 0 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n708, new_n709, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n727, new_n728, new_n730,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n810, new_n811, new_n813, new_n814,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n878, new_n879, new_n881, new_n882,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n895, new_n896, new_n897, new_n899,
    new_n900, new_n901, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n919, new_n921, new_n922, new_n923, new_n924,
    new_n926, new_n927;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT0), .ZN(new_n203));
  XNOR2_X1  g002(.A(G57gat), .B(G85gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  XNOR2_X1  g004(.A(G127gat), .B(G134gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(KEYINPUT70), .B(KEYINPUT1), .ZN(new_n207));
  INV_X1    g006(.A(G113gat), .ZN(new_n208));
  INV_X1    g007(.A(G120gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n206), .A2(new_n207), .A3(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n208), .A2(KEYINPUT69), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT69), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(G113gat), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n209), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  OAI21_X1  g014(.A(KEYINPUT71), .B1(new_n211), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n212), .A2(new_n214), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(G120gat), .ZN(new_n218));
  OR2_X1    g017(.A1(KEYINPUT70), .A2(KEYINPUT1), .ZN(new_n219));
  NAND2_X1  g018(.A1(KEYINPUT70), .A2(KEYINPUT1), .ZN(new_n220));
  AOI22_X1  g019(.A1(new_n219), .A2(new_n220), .B1(new_n208), .B2(new_n209), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT71), .ZN(new_n222));
  NAND4_X1  g021(.A1(new_n218), .A2(new_n221), .A3(new_n222), .A4(new_n206), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n216), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT1), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n225), .B1(G113gat), .B2(G120gat), .ZN(new_n226));
  AND2_X1   g025(.A1(G113gat), .A2(G120gat), .ZN(new_n227));
  OAI22_X1  g026(.A1(new_n226), .A2(new_n227), .B1(G127gat), .B2(G134gat), .ZN(new_n228));
  INV_X1    g027(.A(G127gat), .ZN(new_n229));
  OR2_X1    g028(.A1(KEYINPUT68), .A2(G134gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(KEYINPUT68), .A2(G134gat), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n229), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n228), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n224), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(KEYINPUT72), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT79), .ZN(new_n237));
  NAND2_X1  g036(.A1(G141gat), .A2(G148gat), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  NOR2_X1   g038(.A1(G141gat), .A2(G148gat), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n237), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(G141gat), .ZN(new_n242));
  INV_X1    g041(.A(G148gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n244), .A2(KEYINPUT79), .A3(new_n238), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT2), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n241), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  XOR2_X1   g046(.A(G155gat), .B(G162gat), .Z(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT80), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n247), .A2(KEYINPUT80), .A3(new_n248), .ZN(new_n252));
  INV_X1    g051(.A(G155gat), .ZN(new_n253));
  INV_X1    g052(.A(G162gat), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NOR3_X1   g054(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n256));
  OAI211_X1 g055(.A(new_n244), .B(new_n238), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  AND3_X1   g056(.A1(new_n251), .A2(new_n252), .A3(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n233), .B1(new_n216), .B2(new_n223), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT72), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n236), .A2(new_n258), .A3(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n258), .A2(KEYINPUT4), .A3(new_n259), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n251), .A2(new_n252), .A3(new_n257), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(KEYINPUT3), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT3), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n251), .A2(new_n269), .A3(new_n252), .A4(new_n257), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n268), .A2(new_n270), .A3(new_n235), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT5), .ZN(new_n272));
  NAND2_X1  g071(.A1(G225gat), .A2(G233gat), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n271), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n266), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n271), .A2(new_n273), .ZN(new_n277));
  NOR3_X1   g076(.A1(new_n267), .A2(new_n235), .A3(KEYINPUT4), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n262), .A2(KEYINPUT4), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n278), .B1(new_n279), .B2(KEYINPUT81), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT81), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n262), .A2(new_n281), .A3(KEYINPUT4), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n277), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n267), .B(new_n259), .ZN(new_n284));
  OAI21_X1  g083(.A(KEYINPUT5), .B1(new_n284), .B2(new_n273), .ZN(new_n285));
  OAI211_X1 g084(.A(new_n205), .B(new_n276), .C1(new_n283), .C2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(KEYINPUT82), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n276), .B1(new_n283), .B2(new_n285), .ZN(new_n288));
  INV_X1    g087(.A(new_n205), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(KEYINPUT6), .B1(new_n287), .B2(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n260), .B1(new_n224), .B2(new_n234), .ZN(new_n292));
  AOI211_X1 g091(.A(KEYINPUT72), .B(new_n233), .C1(new_n216), .C2(new_n223), .ZN(new_n293));
  NOR3_X1   g092(.A1(new_n292), .A2(new_n293), .A3(new_n267), .ZN(new_n294));
  OAI21_X1  g093(.A(KEYINPUT81), .B1(new_n294), .B2(new_n263), .ZN(new_n295));
  INV_X1    g094(.A(new_n278), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n295), .A2(new_n282), .A3(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n277), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n285), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT82), .ZN(new_n302));
  NAND4_X1  g101(.A1(new_n301), .A2(new_n302), .A3(new_n205), .A4(new_n276), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT6), .ZN(new_n304));
  AOI22_X1  g103(.A1(new_n303), .A2(new_n304), .B1(new_n289), .B2(new_n288), .ZN(new_n305));
  XNOR2_X1  g104(.A(KEYINPUT27), .B(G183gat), .ZN(new_n306));
  INV_X1    g105(.A(G190gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n308), .B(KEYINPUT28), .ZN(new_n309));
  NAND2_X1  g108(.A1(G183gat), .A2(G190gat), .ZN(new_n310));
  NOR2_X1   g109(.A1(G169gat), .A2(G176gat), .ZN(new_n311));
  XOR2_X1   g110(.A(new_n311), .B(KEYINPUT26), .Z(new_n312));
  NAND2_X1  g111(.A1(G169gat), .A2(G176gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(KEYINPUT65), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT65), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n315), .A2(G169gat), .A3(G176gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n310), .B1(new_n312), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n310), .A2(KEYINPUT24), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT24), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n321), .A2(G183gat), .A3(G190gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT66), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n324), .B1(G183gat), .B2(G190gat), .ZN(new_n325));
  INV_X1    g124(.A(G183gat), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n326), .A2(new_n307), .A3(KEYINPUT66), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n323), .A2(new_n325), .A3(new_n327), .ZN(new_n328));
  OAI21_X1  g127(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT23), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n311), .A2(new_n330), .ZN(new_n331));
  AOI22_X1  g130(.A1(new_n329), .A2(new_n331), .B1(new_n314), .B2(new_n316), .ZN(new_n332));
  AND3_X1   g131(.A1(new_n328), .A2(KEYINPUT25), .A3(new_n332), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n323), .B1(G183gat), .B2(G190gat), .ZN(new_n334));
  AOI21_X1  g133(.A(KEYINPUT25), .B1(new_n334), .B2(new_n332), .ZN(new_n335));
  OAI22_X1  g134(.A1(new_n309), .A2(new_n319), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(G226gat), .ZN(new_n337));
  INV_X1    g136(.A(G233gat), .ZN(new_n338));
  OR3_X1    g137(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(G197gat), .B(G204gat), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT22), .ZN(new_n341));
  INV_X1    g140(.A(G211gat), .ZN(new_n342));
  INV_X1    g141(.A(G218gat), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n341), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n340), .A2(new_n344), .ZN(new_n345));
  XNOR2_X1  g144(.A(G211gat), .B(G218gat), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n346), .A2(new_n340), .A3(new_n344), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n348), .A2(KEYINPUT76), .A3(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT76), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n345), .A2(new_n351), .A3(new_n347), .ZN(new_n352));
  AND2_X1   g151(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n337), .A2(new_n338), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n355), .A2(KEYINPUT29), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n309), .A2(new_n319), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n334), .A2(new_n332), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT25), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n326), .A2(KEYINPUT24), .ZN(new_n362));
  AOI22_X1  g161(.A1(new_n362), .A2(G190gat), .B1(KEYINPUT24), .B2(new_n310), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n327), .A2(new_n325), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n332), .B(KEYINPUT25), .C1(new_n363), .C2(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n361), .A2(new_n365), .A3(KEYINPUT67), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT67), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n367), .B1(new_n333), .B2(new_n335), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n358), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  OAI211_X1 g168(.A(new_n339), .B(new_n354), .C1(new_n357), .C2(new_n369), .ZN(new_n370));
  XOR2_X1   g169(.A(G8gat), .B(G36gat), .Z(new_n371));
  XNOR2_X1  g170(.A(new_n371), .B(KEYINPUT77), .ZN(new_n372));
  XNOR2_X1  g171(.A(G64gat), .B(G92gat), .ZN(new_n373));
  XOR2_X1   g172(.A(new_n372), .B(new_n373), .Z(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  AOI22_X1  g174(.A1(new_n369), .A2(new_n355), .B1(new_n336), .B2(new_n356), .ZN(new_n376));
  OAI211_X1 g175(.A(new_n370), .B(new_n375), .C1(new_n354), .C2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(KEYINPUT78), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(KEYINPUT30), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT30), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n377), .A2(KEYINPUT78), .A3(new_n380), .ZN(new_n381));
  OR2_X1    g180(.A1(new_n376), .A2(new_n354), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(new_n370), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(new_n374), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n379), .A2(new_n381), .A3(new_n384), .ZN(new_n385));
  NOR3_X1   g184(.A1(new_n291), .A2(new_n305), .A3(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT85), .ZN(new_n387));
  NAND2_X1  g186(.A1(G227gat), .A2(G233gat), .ZN(new_n388));
  XOR2_X1   g187(.A(new_n388), .B(KEYINPUT64), .Z(new_n389));
  NOR3_X1   g188(.A1(new_n333), .A2(new_n335), .A3(new_n367), .ZN(new_n390));
  AOI21_X1  g189(.A(KEYINPUT67), .B1(new_n361), .B2(new_n365), .ZN(new_n391));
  OAI22_X1  g190(.A1(new_n390), .A2(new_n391), .B1(new_n309), .B2(new_n319), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT73), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n236), .A2(new_n393), .A3(new_n261), .ZN(new_n394));
  OAI21_X1  g193(.A(KEYINPUT73), .B1(new_n292), .B2(new_n293), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n392), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NOR3_X1   g195(.A1(new_n292), .A2(new_n293), .A3(KEYINPUT73), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n397), .A2(new_n369), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n389), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT33), .ZN(new_n400));
  XOR2_X1   g199(.A(G15gat), .B(G43gat), .Z(new_n401));
  XNOR2_X1  g200(.A(G71gat), .B(G99gat), .ZN(new_n402));
  XNOR2_X1  g201(.A(new_n401), .B(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n399), .B(KEYINPUT32), .C1(new_n400), .C2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n399), .A2(KEYINPUT32), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n399), .A2(new_n400), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n406), .A2(new_n407), .A3(new_n403), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n393), .B1(new_n236), .B2(new_n261), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n369), .B1(new_n409), .B2(new_n397), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n392), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n389), .A2(KEYINPUT34), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n388), .ZN(new_n414));
  NOR3_X1   g213(.A1(new_n396), .A2(new_n398), .A3(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT34), .ZN(new_n416));
  OAI211_X1 g215(.A(KEYINPUT74), .B(new_n413), .C1(new_n415), .C2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n410), .A2(new_n388), .A3(new_n411), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(KEYINPUT34), .ZN(new_n420));
  AOI21_X1  g219(.A(KEYINPUT74), .B1(new_n420), .B2(new_n413), .ZN(new_n421));
  OAI211_X1 g220(.A(new_n405), .B(new_n408), .C1(new_n418), .C2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n408), .A2(new_n405), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(new_n417), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT29), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n270), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(new_n354), .ZN(new_n427));
  AOI21_X1  g226(.A(KEYINPUT29), .B1(new_n348), .B2(new_n349), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n267), .B1(KEYINPUT3), .B2(new_n428), .ZN(new_n429));
  AOI22_X1  g228(.A1(new_n427), .A2(new_n429), .B1(G228gat), .B2(G233gat), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  XOR2_X1   g230(.A(KEYINPUT31), .B(G50gat), .Z(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n353), .B1(new_n426), .B2(KEYINPUT83), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT83), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n270), .A2(new_n435), .A3(new_n425), .ZN(new_n436));
  AND2_X1   g235(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(KEYINPUT3), .B1(new_n353), .B2(new_n425), .ZN(new_n438));
  OAI211_X1 g237(.A(G228gat), .B(G233gat), .C1(new_n438), .C2(new_n258), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n431), .B(new_n433), .C1(new_n437), .C2(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n439), .B1(new_n436), .B2(new_n434), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n432), .B1(new_n441), .B2(new_n430), .ZN(new_n442));
  XNOR2_X1  g241(.A(G78gat), .B(G106gat), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n443), .B(G22gat), .ZN(new_n444));
  AND3_X1   g243(.A1(new_n440), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n444), .B1(new_n440), .B2(new_n442), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n422), .A2(new_n424), .A3(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n386), .A2(new_n387), .A3(new_n449), .A4(KEYINPUT35), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n448), .A2(KEYINPUT35), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT35), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n275), .B1(new_n299), .B2(new_n300), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n302), .B1(new_n453), .B2(new_n205), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n453), .A2(new_n205), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n304), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n304), .B1(new_n286), .B2(KEYINPUT82), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(new_n290), .ZN(new_n458));
  INV_X1    g257(.A(new_n385), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n456), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n422), .A2(new_n424), .A3(new_n447), .A4(new_n387), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n451), .B(new_n452), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n422), .A2(new_n424), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT75), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT36), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  NOR2_X1   g266(.A1(KEYINPUT75), .A2(KEYINPUT36), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n463), .A2(new_n467), .A3(new_n469), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n422), .A2(new_n424), .A3(new_n464), .A4(new_n465), .ZN(new_n471));
  XOR2_X1   g270(.A(KEYINPUT84), .B(KEYINPUT37), .Z(new_n472));
  NAND3_X1  g271(.A1(new_n382), .A2(new_n370), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(new_n374), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT37), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n475), .B1(new_n382), .B2(new_n370), .ZN(new_n476));
  OAI21_X1  g275(.A(KEYINPUT38), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT38), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n339), .B(new_n353), .C1(new_n357), .C2(new_n369), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n479), .B(KEYINPUT37), .C1(new_n353), .C2(new_n376), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n473), .A2(new_n478), .A3(new_n480), .A4(new_n374), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n477), .A2(new_n377), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n482), .B1(new_n456), .B2(new_n458), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT39), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n484), .B1(new_n284), .B2(new_n273), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n264), .A2(new_n271), .A3(new_n265), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n485), .B1(new_n487), .B2(new_n273), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n486), .A2(new_n484), .A3(G225gat), .A4(G233gat), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n488), .A2(new_n205), .A3(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT40), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n488), .A2(KEYINPUT40), .A3(new_n205), .A4(new_n489), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n385), .A2(new_n492), .A3(new_n290), .A4(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(new_n447), .ZN(new_n495));
  OAI211_X1 g294(.A(new_n470), .B(new_n471), .C1(new_n483), .C2(new_n495), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n386), .A2(new_n447), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n450), .B(new_n462), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  XOR2_X1   g297(.A(G15gat), .B(G22gat), .Z(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(G1gat), .ZN(new_n500));
  INV_X1    g299(.A(G1gat), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(KEYINPUT16), .ZN(new_n502));
  OAI221_X1 g301(.A(new_n500), .B1(KEYINPUT92), .B2(G8gat), .C1(new_n499), .C2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(KEYINPUT92), .A2(G8gat), .ZN(new_n504));
  XOR2_X1   g303(.A(new_n503), .B(new_n504), .Z(new_n505));
  XOR2_X1   g304(.A(new_n505), .B(KEYINPUT93), .Z(new_n506));
  XNOR2_X1  g305(.A(G43gat), .B(G50gat), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT87), .ZN(new_n508));
  OR2_X1    g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n507), .A2(new_n508), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n509), .A2(KEYINPUT15), .A3(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(G29gat), .ZN(new_n512));
  INV_X1    g311(.A(G36gat), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  OAI21_X1  g313(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT14), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n517), .A2(new_n512), .A3(new_n513), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n516), .B1(new_n518), .B2(KEYINPUT88), .ZN(new_n519));
  OR2_X1    g318(.A1(new_n518), .A2(KEYINPUT88), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n514), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n511), .A2(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n522), .B(KEYINPUT89), .ZN(new_n523));
  XNOR2_X1  g322(.A(KEYINPUT90), .B(G43gat), .ZN(new_n524));
  INV_X1    g323(.A(G50gat), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  OR2_X1    g325(.A1(new_n525), .A2(G43gat), .ZN(new_n527));
  AOI21_X1  g326(.A(KEYINPUT15), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n528), .B(KEYINPUT91), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n514), .B1(new_n518), .B2(new_n515), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n529), .A2(new_n511), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n523), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n506), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(G229gat), .A2(G233gat), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT17), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n523), .A2(KEYINPUT17), .A3(new_n531), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n536), .A2(new_n505), .A3(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n533), .A2(new_n534), .A3(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT18), .ZN(new_n540));
  OR2_X1    g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n506), .B(new_n532), .ZN(new_n542));
  XOR2_X1   g341(.A(new_n534), .B(KEYINPUT13), .Z(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n539), .A2(new_n540), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n541), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(G113gat), .B(G141gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(G197gat), .ZN(new_n548));
  XOR2_X1   g347(.A(KEYINPUT11), .B(G169gat), .Z(new_n549));
  XNOR2_X1  g348(.A(new_n548), .B(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(KEYINPUT86), .B(KEYINPUT12), .ZN(new_n551));
  XOR2_X1   g350(.A(new_n550), .B(new_n551), .Z(new_n552));
  NAND2_X1  g351(.A1(new_n546), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n552), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n541), .A2(new_n554), .A3(new_n544), .A4(new_n545), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  AND2_X1   g355(.A1(new_n498), .A2(new_n556), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n291), .A2(new_n305), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(KEYINPUT97), .B(KEYINPUT7), .ZN(new_n560));
  AND2_X1   g359(.A1(G85gat), .A2(G92gat), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n560), .B(new_n561), .ZN(new_n562));
  XOR2_X1   g361(.A(KEYINPUT98), .B(G85gat), .Z(new_n563));
  INV_X1    g362(.A(G92gat), .ZN(new_n564));
  NAND2_X1  g363(.A1(G99gat), .A2(G106gat), .ZN(new_n565));
  AOI22_X1  g364(.A1(new_n563), .A2(new_n564), .B1(KEYINPUT8), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n562), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT100), .ZN(new_n568));
  XNOR2_X1  g367(.A(G99gat), .B(G106gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n569), .B(KEYINPUT99), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n567), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n568), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n536), .A2(new_n537), .A3(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n573), .ZN(new_n575));
  AND2_X1   g374(.A1(G232gat), .A2(G233gat), .ZN(new_n576));
  AOI22_X1  g375(.A1(new_n575), .A2(new_n532), .B1(KEYINPUT41), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(G190gat), .B(G218gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n576), .A2(KEYINPUT41), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(KEYINPUT96), .ZN(new_n582));
  XNOR2_X1  g381(.A(G134gat), .B(G162gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n580), .B(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(G64gat), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(G57gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(KEYINPUT95), .B(G57gat), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n588), .B1(new_n590), .B2(new_n587), .ZN(new_n591));
  NOR2_X1   g390(.A1(G71gat), .A2(G78gat), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(KEYINPUT9), .ZN(new_n593));
  NAND2_X1  g392(.A1(G71gat), .A2(G78gat), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g395(.A1(KEYINPUT94), .A2(KEYINPUT9), .ZN(new_n597));
  OR2_X1    g396(.A1(new_n587), .A2(G57gat), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n597), .B1(new_n598), .B2(new_n588), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n592), .B1(KEYINPUT94), .B2(new_n594), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n600), .B1(KEYINPUT94), .B2(new_n594), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n596), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n506), .B1(KEYINPUT21), .B2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT21), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(G231gat), .A2(G233gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(G127gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n604), .B(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(G155gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(G183gat), .B(G211gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n610), .B(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n586), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n573), .A2(new_n602), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT101), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n573), .A2(KEYINPUT101), .A3(new_n602), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n567), .A2(KEYINPUT102), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n570), .B1(new_n621), .B2(KEYINPUT103), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n570), .A2(KEYINPUT103), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n567), .B1(new_n623), .B2(KEYINPUT102), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  AOI22_X1  g424(.A1(new_n619), .A2(new_n620), .B1(new_n603), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(G230gat), .A2(G233gat), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(G120gat), .B(G148gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(G176gat), .B(G204gat), .ZN(new_n631));
  XOR2_X1   g430(.A(new_n630), .B(new_n631), .Z(new_n632));
  INV_X1    g431(.A(KEYINPUT10), .ZN(new_n633));
  NOR3_X1   g432(.A1(new_n573), .A2(new_n633), .A3(new_n602), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n634), .B1(new_n626), .B2(new_n633), .ZN(new_n635));
  INV_X1    g434(.A(new_n627), .ZN(new_n636));
  OAI211_X1 g435(.A(new_n629), .B(new_n632), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n632), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n619), .A2(new_n620), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n625), .A2(new_n603), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n639), .A2(new_n633), .A3(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n634), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n636), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n638), .B1(new_n643), .B2(new_n628), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n637), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n616), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n557), .A2(new_n559), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(G1gat), .ZN(G1324gat));
  INV_X1    g447(.A(KEYINPUT42), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n557), .A2(new_n646), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n650), .A2(new_n459), .ZN(new_n651));
  XOR2_X1   g450(.A(KEYINPUT16), .B(G8gat), .Z(new_n652));
  AOI21_X1  g451(.A(new_n649), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g452(.A(G8gat), .B1(new_n650), .B2(new_n459), .ZN(new_n654));
  NOR2_X1   g453(.A1(KEYINPUT104), .A2(KEYINPUT42), .ZN(new_n655));
  MUX2_X1   g454(.A(KEYINPUT104), .B(new_n655), .S(new_n652), .Z(new_n656));
  AOI22_X1  g455(.A1(new_n653), .A2(new_n654), .B1(new_n651), .B2(new_n656), .ZN(G1325gat));
  INV_X1    g456(.A(new_n650), .ZN(new_n658));
  INV_X1    g457(.A(new_n463), .ZN(new_n659));
  AOI21_X1  g458(.A(G15gat), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  AOI211_X1 g459(.A(new_n466), .B(new_n468), .C1(new_n422), .C2(new_n424), .ZN(new_n661));
  AND4_X1   g460(.A1(new_n464), .A2(new_n422), .A3(new_n424), .A4(new_n465), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(G15gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(KEYINPUT105), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n660), .B1(new_n658), .B2(new_n666), .ZN(G1326gat));
  NOR2_X1   g466(.A1(new_n650), .A2(new_n447), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(KEYINPUT106), .ZN(new_n669));
  XNOR2_X1  g468(.A(KEYINPUT43), .B(G22gat), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(G1327gat));
  INV_X1    g470(.A(new_n615), .ZN(new_n672));
  INV_X1    g471(.A(new_n645), .ZN(new_n673));
  AND4_X1   g472(.A1(new_n557), .A2(new_n672), .A3(new_n585), .A4(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n674), .A2(new_n512), .A3(new_n559), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(KEYINPUT45), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT44), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n677), .B1(new_n498), .B2(new_n585), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n585), .A2(new_n677), .ZN(new_n679));
  AND2_X1   g478(.A1(new_n462), .A2(new_n450), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT108), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n681), .B1(new_n386), .B2(new_n447), .ZN(new_n682));
  OAI211_X1 g481(.A(new_n447), .B(new_n494), .C1(new_n558), .C2(new_n482), .ZN(new_n683));
  INV_X1    g482(.A(new_n447), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n460), .A2(KEYINPUT108), .A3(new_n684), .ZN(new_n685));
  NAND4_X1  g484(.A1(new_n682), .A2(new_n663), .A3(new_n683), .A4(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n679), .B1(new_n680), .B2(new_n686), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n678), .A2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n556), .ZN(new_n689));
  XOR2_X1   g488(.A(new_n645), .B(KEYINPUT107), .Z(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  NOR4_X1   g490(.A1(new_n688), .A2(new_n689), .A3(new_n615), .A4(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(new_n559), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n676), .B1(new_n694), .B2(new_n512), .ZN(G1328gat));
  NAND3_X1  g494(.A1(new_n674), .A2(new_n513), .A3(new_n385), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(KEYINPUT46), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n513), .B1(new_n692), .B2(new_n385), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(KEYINPUT109), .ZN(G1329gat));
  AOI21_X1  g499(.A(new_n524), .B1(new_n674), .B2(new_n659), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n701), .B1(KEYINPUT110), .B2(KEYINPUT47), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n692), .A2(new_n664), .A3(new_n524), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g503(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n705));
  XOR2_X1   g504(.A(new_n704), .B(new_n705), .Z(G1330gat));
  AOI21_X1  g505(.A(new_n525), .B1(new_n692), .B2(new_n684), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n447), .A2(G50gat), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n707), .B1(new_n674), .B2(new_n708), .ZN(new_n709));
  XOR2_X1   g508(.A(KEYINPUT111), .B(KEYINPUT48), .Z(new_n710));
  XNOR2_X1  g509(.A(new_n709), .B(new_n710), .ZN(G1331gat));
  NAND2_X1  g510(.A1(new_n680), .A2(new_n686), .ZN(new_n712));
  NOR3_X1   g511(.A1(new_n690), .A2(new_n616), .A3(new_n556), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(new_n559), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT112), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(new_n589), .ZN(G1332gat));
  XOR2_X1   g517(.A(new_n385), .B(KEYINPUT113), .Z(new_n719));
  NOR2_X1   g518(.A1(new_n714), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g519(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n721));
  AND2_X1   g520(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n720), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n723), .B1(new_n720), .B2(new_n721), .ZN(G1333gat));
  NOR3_X1   g523(.A1(new_n714), .A2(G71gat), .A3(new_n463), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n715), .A2(new_n664), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n725), .B1(G71gat), .B2(new_n726), .ZN(new_n727));
  XNOR2_X1  g526(.A(KEYINPUT114), .B(KEYINPUT50), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n727), .B(new_n728), .ZN(G1334gat));
  NAND2_X1  g528(.A1(new_n715), .A2(new_n684), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g530(.A1(new_n556), .A2(new_n586), .A3(new_n615), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n712), .A2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT51), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n712), .A2(KEYINPUT51), .A3(new_n732), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n737), .A2(new_n559), .A3(new_n563), .A4(new_n645), .ZN(new_n738));
  NOR3_X1   g537(.A1(new_n556), .A2(new_n615), .A3(new_n673), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n739), .B1(new_n678), .B2(new_n687), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(KEYINPUT115), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT115), .ZN(new_n742));
  OAI211_X1 g541(.A(new_n742), .B(new_n739), .C1(new_n678), .C2(new_n687), .ZN(new_n743));
  AND2_X1   g542(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  AND2_X1   g543(.A1(new_n744), .A2(new_n559), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n738), .B1(new_n745), .B2(new_n563), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(KEYINPUT116), .ZN(G1336gat));
  INV_X1    g546(.A(new_n719), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n737), .A2(new_n564), .A3(new_n691), .A4(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT52), .ZN(new_n750));
  OAI21_X1  g549(.A(G92gat), .B1(new_n740), .B2(new_n719), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n749), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(new_n749), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n744), .A2(new_n385), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n753), .B1(new_n754), .B2(G92gat), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n752), .B1(new_n755), .B2(new_n750), .ZN(G1337gat));
  AND2_X1   g555(.A1(new_n744), .A2(new_n664), .ZN(new_n757));
  INV_X1    g556(.A(G99gat), .ZN(new_n758));
  INV_X1    g557(.A(new_n737), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n659), .A2(new_n758), .A3(new_n645), .ZN(new_n760));
  OAI22_X1  g559(.A1(new_n757), .A2(new_n758), .B1(new_n759), .B2(new_n760), .ZN(G1338gat));
  NOR3_X1   g560(.A1(new_n690), .A2(G106gat), .A3(new_n447), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n763), .B1(new_n735), .B2(new_n736), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT53), .ZN(new_n766));
  OAI21_X1  g565(.A(G106gat), .B1(new_n740), .B2(new_n447), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n765), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n741), .A2(new_n684), .A3(new_n743), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(G106gat), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(new_n765), .ZN(new_n771));
  AOI21_X1  g570(.A(KEYINPUT117), .B1(new_n771), .B2(KEYINPUT53), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n764), .B1(new_n769), .B2(G106gat), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT117), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n773), .A2(new_n774), .A3(new_n766), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n768), .B1(new_n772), .B2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT118), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  OAI211_X1 g577(.A(KEYINPUT118), .B(new_n768), .C1(new_n772), .C2(new_n775), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(G1339gat));
  AOI21_X1  g579(.A(new_n534), .B1(new_n533), .B2(new_n538), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT119), .ZN(new_n782));
  OAI22_X1  g581(.A1(new_n542), .A2(new_n543), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  AND2_X1   g582(.A1(new_n781), .A2(new_n782), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n550), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n785), .A2(new_n555), .ZN(new_n786));
  AND2_X1   g585(.A1(new_n786), .A2(new_n585), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n641), .A2(new_n642), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(new_n627), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n641), .A2(new_n636), .A3(new_n642), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n789), .A2(KEYINPUT54), .A3(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT54), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n632), .B1(new_n643), .B2(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n791), .A2(KEYINPUT55), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(new_n637), .ZN(new_n795));
  AOI21_X1  g594(.A(KEYINPUT55), .B1(new_n791), .B2(new_n793), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n787), .A2(new_n797), .ZN(new_n798));
  AOI22_X1  g597(.A1(new_n797), .A2(new_n556), .B1(new_n645), .B2(new_n786), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n798), .B1(new_n799), .B2(new_n585), .ZN(new_n800));
  AOI22_X1  g599(.A1(new_n800), .A2(new_n672), .B1(new_n689), .B2(new_n646), .ZN(new_n801));
  NOR3_X1   g600(.A1(new_n801), .A2(new_n558), .A3(new_n448), .ZN(new_n802));
  AND2_X1   g601(.A1(new_n802), .A2(new_n719), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n803), .A2(new_n212), .A3(new_n214), .A4(new_n556), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n801), .A2(new_n684), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n748), .A2(new_n558), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n805), .A2(new_n659), .A3(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(G113gat), .B1(new_n807), .B2(new_n689), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n804), .A2(new_n808), .ZN(G1340gat));
  NOR3_X1   g608(.A1(new_n807), .A2(new_n209), .A3(new_n690), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n803), .A2(new_n645), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n810), .B1(new_n811), .B2(new_n209), .ZN(G1341gat));
  NAND3_X1  g611(.A1(new_n803), .A2(new_n229), .A3(new_n615), .ZN(new_n813));
  OAI21_X1  g612(.A(G127gat), .B1(new_n807), .B2(new_n672), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(G1342gat));
  NOR2_X1   g614(.A1(new_n586), .A2(new_n385), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n802), .A2(new_n230), .A3(new_n231), .A4(new_n816), .ZN(new_n817));
  OR2_X1    g616(.A1(new_n817), .A2(KEYINPUT56), .ZN(new_n818));
  OAI21_X1  g617(.A(G134gat), .B1(new_n807), .B2(new_n586), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n817), .A2(KEYINPUT56), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n818), .A2(new_n819), .A3(new_n820), .ZN(G1343gat));
  NAND2_X1  g620(.A1(new_n806), .A2(new_n663), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT57), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n447), .A2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT121), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n825), .B1(new_n795), .B2(new_n796), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n791), .A2(new_n793), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT55), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n829), .A2(KEYINPUT121), .A3(new_n637), .A4(new_n794), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n826), .A2(new_n830), .A3(new_n556), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n785), .A2(new_n645), .A3(new_n555), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(KEYINPUT120), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT120), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n785), .A2(new_n645), .A3(new_n834), .A4(new_n555), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n585), .B1(new_n831), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n798), .B1(new_n837), .B2(KEYINPUT122), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT122), .ZN(new_n839));
  AOI211_X1 g638(.A(new_n839), .B(new_n585), .C1(new_n831), .C2(new_n836), .ZN(new_n840));
  OAI211_X1 g639(.A(KEYINPUT123), .B(new_n672), .C1(new_n838), .C2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n646), .A2(new_n689), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n833), .A2(new_n835), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n829), .A2(new_n637), .A3(new_n794), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n689), .B1(new_n845), .B2(new_n825), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n844), .B1(new_n846), .B2(new_n830), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n839), .B1(new_n847), .B2(new_n585), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n837), .A2(KEYINPUT122), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n848), .A2(new_n798), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(KEYINPUT123), .B1(new_n850), .B2(new_n672), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n824), .B1(new_n843), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n823), .B1(new_n801), .B2(new_n447), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n822), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n242), .B1(new_n854), .B2(new_n556), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n801), .A2(new_n558), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n664), .A2(new_n447), .ZN(new_n857));
  AND3_X1   g656(.A1(new_n856), .A2(new_n719), .A3(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n858), .A2(new_n242), .A3(new_n556), .ZN(new_n859));
  INV_X1    g658(.A(new_n859), .ZN(new_n860));
  OAI21_X1  g659(.A(KEYINPUT58), .B1(new_n855), .B2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT58), .ZN(new_n862));
  AOI211_X1 g661(.A(new_n689), .B(new_n822), .C1(new_n852), .C2(new_n853), .ZN(new_n863));
  OAI211_X1 g662(.A(new_n862), .B(new_n859), .C1(new_n863), .C2(new_n242), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n861), .A2(new_n864), .ZN(G1344gat));
  NAND3_X1  g664(.A1(new_n858), .A2(new_n243), .A3(new_n645), .ZN(new_n866));
  XNOR2_X1  g665(.A(new_n866), .B(KEYINPUT124), .ZN(new_n867));
  AOI211_X1 g666(.A(KEYINPUT59), .B(new_n243), .C1(new_n854), .C2(new_n645), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT59), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n837), .B1(new_n797), .B2(new_n787), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n842), .B1(new_n870), .B2(new_n615), .ZN(new_n871));
  AOI21_X1  g670(.A(KEYINPUT57), .B1(new_n871), .B2(new_n684), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n801), .A2(new_n823), .A3(new_n447), .ZN(new_n873));
  OR2_X1    g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n874), .A2(new_n663), .A3(new_n645), .A4(new_n806), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n869), .B1(new_n875), .B2(G148gat), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n867), .B1(new_n868), .B2(new_n876), .ZN(G1345gat));
  NAND3_X1  g676(.A1(new_n858), .A2(new_n253), .A3(new_n615), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n854), .A2(new_n615), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n878), .B1(new_n879), .B2(new_n253), .ZN(G1346gat));
  NAND4_X1  g679(.A1(new_n856), .A2(new_n254), .A3(new_n816), .A4(new_n857), .ZN(new_n881));
  AND2_X1   g680(.A1(new_n854), .A2(new_n585), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n881), .B1(new_n882), .B2(new_n254), .ZN(G1347gat));
  NOR2_X1   g682(.A1(new_n801), .A2(new_n559), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n719), .A2(new_n448), .ZN(new_n885));
  XNOR2_X1  g684(.A(new_n885), .B(KEYINPUT125), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(G169gat), .B1(new_n888), .B2(new_n556), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n559), .A2(new_n459), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  NOR4_X1   g690(.A1(new_n801), .A2(new_n684), .A3(new_n463), .A4(new_n891), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n556), .A2(G169gat), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n889), .B1(new_n892), .B2(new_n893), .ZN(G1348gat));
  INV_X1    g693(.A(G176gat), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n888), .A2(new_n895), .A3(new_n645), .ZN(new_n896));
  AND2_X1   g695(.A1(new_n892), .A2(new_n691), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n896), .B1(new_n895), .B2(new_n897), .ZN(G1349gat));
  NAND3_X1  g697(.A1(new_n888), .A2(new_n306), .A3(new_n615), .ZN(new_n899));
  AND2_X1   g698(.A1(new_n892), .A2(new_n615), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n899), .B1(new_n900), .B2(new_n326), .ZN(new_n901));
  XNOR2_X1  g700(.A(new_n901), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g701(.A1(new_n888), .A2(new_n307), .A3(new_n585), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n892), .A2(new_n585), .ZN(new_n904));
  XNOR2_X1  g703(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n905));
  AND3_X1   g704(.A1(new_n904), .A2(G190gat), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n905), .B1(new_n904), .B2(G190gat), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n903), .B1(new_n906), .B2(new_n907), .ZN(G1351gat));
  AND3_X1   g707(.A1(new_n884), .A2(new_n748), .A3(new_n857), .ZN(new_n909));
  AOI21_X1  g708(.A(G197gat), .B1(new_n909), .B2(new_n556), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n891), .A2(new_n664), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n874), .A2(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(new_n912), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n556), .A2(G197gat), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n910), .B1(new_n913), .B2(new_n914), .ZN(G1352gat));
  INV_X1    g714(.A(G204gat), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n909), .A2(new_n916), .A3(new_n645), .ZN(new_n917));
  XOR2_X1   g716(.A(new_n917), .B(KEYINPUT62), .Z(new_n918));
  OAI21_X1  g717(.A(G204gat), .B1(new_n912), .B2(new_n690), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(G1353gat));
  NAND3_X1  g719(.A1(new_n909), .A2(new_n342), .A3(new_n615), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n874), .A2(new_n615), .A3(new_n911), .ZN(new_n922));
  AND3_X1   g721(.A1(new_n922), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n923));
  AOI21_X1  g722(.A(KEYINPUT63), .B1(new_n922), .B2(G211gat), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n921), .B1(new_n923), .B2(new_n924), .ZN(G1354gat));
  OAI21_X1  g724(.A(G218gat), .B1(new_n912), .B2(new_n586), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n909), .A2(new_n343), .A3(new_n585), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(G1355gat));
endmodule


