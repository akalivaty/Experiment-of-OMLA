

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590;

  XNOR2_X1 U320 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U321 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U322 ( .A(n372), .B(n371), .ZN(n397) );
  XNOR2_X1 U323 ( .A(n385), .B(n307), .ZN(n308) );
  XNOR2_X1 U324 ( .A(n309), .B(n308), .ZN(n311) );
  XNOR2_X1 U325 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U326 ( .A(n318), .B(n317), .ZN(n319) );
  INV_X1 U327 ( .A(KEYINPUT64), .ZN(n443) );
  XNOR2_X1 U328 ( .A(n320), .B(n319), .ZN(n324) );
  XNOR2_X1 U329 ( .A(n444), .B(n443), .ZN(n573) );
  AND2_X1 U330 ( .A1(n541), .A2(n461), .ZN(n462) );
  XNOR2_X1 U331 ( .A(n462), .B(KEYINPUT120), .ZN(n570) );
  XNOR2_X1 U332 ( .A(n469), .B(G190GAT), .ZN(n470) );
  XNOR2_X1 U333 ( .A(n471), .B(n470), .ZN(G1351GAT) );
  XOR2_X1 U334 ( .A(G43GAT), .B(G134GAT), .Z(n380) );
  XNOR2_X1 U335 ( .A(G99GAT), .B(G71GAT), .ZN(n288) );
  XNOR2_X1 U336 ( .A(n288), .B(G120GAT), .ZN(n322) );
  XOR2_X1 U337 ( .A(n380), .B(n322), .Z(n290) );
  NAND2_X1 U338 ( .A1(G227GAT), .A2(G233GAT), .ZN(n289) );
  XNOR2_X1 U339 ( .A(n290), .B(n289), .ZN(n301) );
  XOR2_X1 U340 ( .A(G176GAT), .B(KEYINPUT83), .Z(n292) );
  XNOR2_X1 U341 ( .A(KEYINPUT85), .B(KEYINPUT87), .ZN(n291) );
  XNOR2_X1 U342 ( .A(n292), .B(n291), .ZN(n293) );
  XOR2_X1 U343 ( .A(n293), .B(KEYINPUT88), .Z(n295) );
  XOR2_X1 U344 ( .A(G15GAT), .B(G127GAT), .Z(n365) );
  XNOR2_X1 U345 ( .A(n365), .B(KEYINPUT84), .ZN(n294) );
  XNOR2_X1 U346 ( .A(n295), .B(n294), .ZN(n297) );
  XNOR2_X1 U347 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n296) );
  XNOR2_X1 U348 ( .A(n296), .B(KEYINPUT82), .ZN(n439) );
  XOR2_X1 U349 ( .A(n297), .B(n439), .Z(n299) );
  XNOR2_X1 U350 ( .A(KEYINPUT86), .B(KEYINPUT20), .ZN(n298) );
  XNOR2_X1 U351 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U352 ( .A(n301), .B(n300), .ZN(n306) );
  XOR2_X1 U353 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n303) );
  XNOR2_X1 U354 ( .A(G169GAT), .B(G183GAT), .ZN(n302) );
  XNOR2_X1 U355 ( .A(n303), .B(n302), .ZN(n305) );
  XOR2_X1 U356 ( .A(G190GAT), .B(KEYINPUT19), .Z(n304) );
  XNOR2_X1 U357 ( .A(n305), .B(n304), .ZN(n419) );
  XOR2_X1 U358 ( .A(n306), .B(n419), .Z(n479) );
  INV_X1 U359 ( .A(n479), .ZN(n541) );
  XOR2_X1 U360 ( .A(KEYINPUT13), .B(KEYINPUT71), .Z(n352) );
  XNOR2_X1 U361 ( .A(G57GAT), .B(KEYINPUT72), .ZN(n351) );
  XNOR2_X1 U362 ( .A(n352), .B(n351), .ZN(n309) );
  XOR2_X1 U363 ( .A(G85GAT), .B(G92GAT), .Z(n385) );
  AND2_X1 U364 ( .A1(G230GAT), .A2(G233GAT), .ZN(n307) );
  INV_X1 U365 ( .A(KEYINPUT32), .ZN(n310) );
  NAND2_X1 U366 ( .A1(n311), .A2(n310), .ZN(n314) );
  INV_X1 U367 ( .A(n311), .ZN(n312) );
  NAND2_X1 U368 ( .A1(n312), .A2(KEYINPUT32), .ZN(n313) );
  NAND2_X1 U369 ( .A1(n314), .A2(n313), .ZN(n320) );
  XOR2_X1 U370 ( .A(G176GAT), .B(G64GAT), .Z(n404) );
  XNOR2_X1 U371 ( .A(G204GAT), .B(n404), .ZN(n318) );
  XOR2_X1 U372 ( .A(KEYINPUT73), .B(KEYINPUT31), .Z(n316) );
  XNOR2_X1 U373 ( .A(KEYINPUT74), .B(KEYINPUT33), .ZN(n315) );
  XNOR2_X1 U374 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U375 ( .A(G106GAT), .B(G78GAT), .ZN(n321) );
  XNOR2_X1 U376 ( .A(n321), .B(G148GAT), .ZN(n450) );
  XOR2_X1 U377 ( .A(n322), .B(n450), .Z(n323) );
  XNOR2_X1 U378 ( .A(n324), .B(n323), .ZN(n578) );
  XNOR2_X1 U379 ( .A(n578), .B(KEYINPUT41), .ZN(n559) );
  INV_X1 U380 ( .A(G36GAT), .ZN(n325) );
  NAND2_X1 U381 ( .A1(G29GAT), .A2(n325), .ZN(n328) );
  INV_X1 U382 ( .A(G29GAT), .ZN(n326) );
  NAND2_X1 U383 ( .A1(n326), .A2(G36GAT), .ZN(n327) );
  NAND2_X1 U384 ( .A1(n328), .A2(n327), .ZN(n330) );
  XNOR2_X1 U385 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n329) );
  XNOR2_X1 U386 ( .A(n330), .B(n329), .ZN(n381) );
  XOR2_X1 U387 ( .A(n381), .B(KEYINPUT29), .Z(n332) );
  NAND2_X1 U388 ( .A1(G229GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U389 ( .A(n332), .B(n331), .ZN(n347) );
  XOR2_X1 U390 ( .A(G50GAT), .B(G43GAT), .Z(n334) );
  XNOR2_X1 U391 ( .A(G197GAT), .B(G141GAT), .ZN(n333) );
  XNOR2_X1 U392 ( .A(n334), .B(n333), .ZN(n337) );
  XOR2_X1 U393 ( .A(KEYINPUT68), .B(KEYINPUT69), .Z(n336) );
  XNOR2_X1 U394 ( .A(G22GAT), .B(G1GAT), .ZN(n335) );
  XNOR2_X1 U395 ( .A(n336), .B(n335), .ZN(n366) );
  XOR2_X1 U396 ( .A(n337), .B(n366), .Z(n345) );
  XOR2_X1 U397 ( .A(G8GAT), .B(G113GAT), .Z(n339) );
  XNOR2_X1 U398 ( .A(G169GAT), .B(G15GAT), .ZN(n338) );
  XNOR2_X1 U399 ( .A(n339), .B(n338), .ZN(n343) );
  XOR2_X1 U400 ( .A(KEYINPUT70), .B(KEYINPUT30), .Z(n341) );
  XNOR2_X1 U401 ( .A(KEYINPUT67), .B(KEYINPUT66), .ZN(n340) );
  XNOR2_X1 U402 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U403 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U404 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U405 ( .A(n347), .B(n346), .Z(n543) );
  INV_X1 U406 ( .A(n543), .ZN(n574) );
  NAND2_X1 U407 ( .A1(n559), .A2(n574), .ZN(n349) );
  XNOR2_X1 U408 ( .A(KEYINPUT46), .B(KEYINPUT114), .ZN(n348) );
  XNOR2_X1 U409 ( .A(n349), .B(n348), .ZN(n394) );
  XOR2_X1 U410 ( .A(G8GAT), .B(KEYINPUT76), .Z(n407) );
  INV_X1 U411 ( .A(KEYINPUT12), .ZN(n350) );
  XNOR2_X1 U412 ( .A(n351), .B(n350), .ZN(n353) );
  XNOR2_X1 U413 ( .A(n353), .B(n352), .ZN(n355) );
  NAND2_X1 U414 ( .A1(G231GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U415 ( .A(n355), .B(n354), .ZN(n363) );
  XOR2_X1 U416 ( .A(G155GAT), .B(G78GAT), .Z(n357) );
  XNOR2_X1 U417 ( .A(G183GAT), .B(G211GAT), .ZN(n356) );
  XNOR2_X1 U418 ( .A(n357), .B(n356), .ZN(n361) );
  XOR2_X1 U419 ( .A(KEYINPUT79), .B(KEYINPUT80), .Z(n359) );
  XNOR2_X1 U420 ( .A(G71GAT), .B(G64GAT), .ZN(n358) );
  XNOR2_X1 U421 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U422 ( .A(n407), .B(n364), .Z(n372) );
  XNOR2_X1 U423 ( .A(n366), .B(n365), .ZN(n370) );
  XOR2_X1 U424 ( .A(KEYINPUT78), .B(KEYINPUT77), .Z(n368) );
  XNOR2_X1 U425 ( .A(KEYINPUT15), .B(KEYINPUT14), .ZN(n367) );
  XOR2_X1 U426 ( .A(n368), .B(n367), .Z(n369) );
  INV_X1 U427 ( .A(n397), .ZN(n582) );
  XOR2_X1 U428 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n374) );
  XNOR2_X1 U429 ( .A(G99GAT), .B(KEYINPUT9), .ZN(n373) );
  XNOR2_X1 U430 ( .A(n374), .B(n373), .ZN(n376) );
  XOR2_X1 U431 ( .A(G50GAT), .B(G162GAT), .Z(n445) );
  INV_X1 U432 ( .A(n445), .ZN(n375) );
  NAND2_X1 U433 ( .A1(n376), .A2(n375), .ZN(n379) );
  INV_X1 U434 ( .A(n376), .ZN(n377) );
  NAND2_X1 U435 ( .A1(n377), .A2(n445), .ZN(n378) );
  NAND2_X1 U436 ( .A1(n379), .A2(n378), .ZN(n383) );
  XNOR2_X1 U437 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U438 ( .A(n383), .B(n382), .ZN(n384) );
  XOR2_X1 U439 ( .A(n384), .B(KEYINPUT65), .Z(n387) );
  XNOR2_X1 U440 ( .A(G218GAT), .B(n385), .ZN(n386) );
  XNOR2_X1 U441 ( .A(n387), .B(n386), .ZN(n392) );
  XOR2_X1 U442 ( .A(G106GAT), .B(KEYINPUT75), .Z(n389) );
  NAND2_X1 U443 ( .A1(G232GAT), .A2(G233GAT), .ZN(n388) );
  XNOR2_X1 U444 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U445 ( .A(G190GAT), .B(n390), .Z(n391) );
  XOR2_X1 U446 ( .A(n392), .B(n391), .Z(n566) );
  INV_X1 U447 ( .A(n566), .ZN(n551) );
  NOR2_X1 U448 ( .A1(n582), .A2(n566), .ZN(n393) );
  NAND2_X1 U449 ( .A1(n394), .A2(n393), .ZN(n395) );
  XNOR2_X1 U450 ( .A(n395), .B(KEYINPUT47), .ZN(n402) );
  XNOR2_X1 U451 ( .A(KEYINPUT36), .B(KEYINPUT103), .ZN(n396) );
  XOR2_X1 U452 ( .A(n551), .B(n396), .Z(n587) );
  NOR2_X1 U453 ( .A1(n587), .A2(n397), .ZN(n398) );
  XNOR2_X1 U454 ( .A(n398), .B(KEYINPUT45), .ZN(n400) );
  AND2_X1 U455 ( .A1(n578), .A2(n543), .ZN(n399) );
  AND2_X1 U456 ( .A1(n400), .A2(n399), .ZN(n401) );
  NOR2_X1 U457 ( .A1(n402), .A2(n401), .ZN(n403) );
  XNOR2_X1 U458 ( .A(n403), .B(KEYINPUT48), .ZN(n539) );
  XOR2_X1 U459 ( .A(KEYINPUT98), .B(n404), .Z(n406) );
  NAND2_X1 U460 ( .A1(G226GAT), .A2(G233GAT), .ZN(n405) );
  XNOR2_X1 U461 ( .A(n406), .B(n405), .ZN(n408) );
  XOR2_X1 U462 ( .A(n408), .B(n407), .Z(n418) );
  XOR2_X1 U463 ( .A(KEYINPUT21), .B(KEYINPUT93), .Z(n410) );
  XNOR2_X1 U464 ( .A(G218GAT), .B(KEYINPUT92), .ZN(n409) );
  XNOR2_X1 U465 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U466 ( .A(n411), .B(G211GAT), .Z(n413) );
  XNOR2_X1 U467 ( .A(G197GAT), .B(G204GAT), .ZN(n412) );
  XNOR2_X1 U468 ( .A(n413), .B(n412), .ZN(n456) );
  XOR2_X1 U469 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n415) );
  XNOR2_X1 U470 ( .A(G36GAT), .B(G92GAT), .ZN(n414) );
  XNOR2_X1 U471 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U472 ( .A(n456), .B(n416), .ZN(n417) );
  XNOR2_X1 U473 ( .A(n418), .B(n417), .ZN(n420) );
  XOR2_X1 U474 ( .A(n420), .B(n419), .Z(n528) );
  INV_X1 U475 ( .A(n528), .ZN(n474) );
  NOR2_X1 U476 ( .A1(n539), .A2(n474), .ZN(n421) );
  XOR2_X1 U477 ( .A(KEYINPUT54), .B(n421), .Z(n442) );
  XOR2_X1 U478 ( .A(G85GAT), .B(G162GAT), .Z(n423) );
  XNOR2_X1 U479 ( .A(G29GAT), .B(G134GAT), .ZN(n422) );
  XNOR2_X1 U480 ( .A(n423), .B(n422), .ZN(n427) );
  XOR2_X1 U481 ( .A(KEYINPUT4), .B(G148GAT), .Z(n425) );
  XNOR2_X1 U482 ( .A(G120GAT), .B(G127GAT), .ZN(n424) );
  XNOR2_X1 U483 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U484 ( .A(n427), .B(n426), .Z(n432) );
  XOR2_X1 U485 ( .A(KEYINPUT1), .B(G57GAT), .Z(n429) );
  NAND2_X1 U486 ( .A1(G225GAT), .A2(G233GAT), .ZN(n428) );
  XNOR2_X1 U487 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U488 ( .A(KEYINPUT6), .B(n430), .ZN(n431) );
  XNOR2_X1 U489 ( .A(n432), .B(n431), .ZN(n436) );
  XOR2_X1 U490 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n434) );
  XNOR2_X1 U491 ( .A(G1GAT), .B(KEYINPUT5), .ZN(n433) );
  XNOR2_X1 U492 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U493 ( .A(n436), .B(n435), .Z(n441) );
  XOR2_X1 U494 ( .A(G155GAT), .B(KEYINPUT2), .Z(n438) );
  XNOR2_X1 U495 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n437) );
  XNOR2_X1 U496 ( .A(n438), .B(n437), .ZN(n446) );
  XNOR2_X1 U497 ( .A(n439), .B(n446), .ZN(n440) );
  XNOR2_X1 U498 ( .A(n441), .B(n440), .ZN(n555) );
  NOR2_X1 U499 ( .A1(n442), .A2(n555), .ZN(n444) );
  XOR2_X1 U500 ( .A(n446), .B(n445), .Z(n448) );
  NAND2_X1 U501 ( .A1(G228GAT), .A2(G233GAT), .ZN(n447) );
  XNOR2_X1 U502 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U503 ( .A(n449), .B(KEYINPUT90), .Z(n452) );
  XNOR2_X1 U504 ( .A(n450), .B(KEYINPUT24), .ZN(n451) );
  XNOR2_X1 U505 ( .A(n452), .B(n451), .ZN(n458) );
  XOR2_X1 U506 ( .A(KEYINPUT91), .B(KEYINPUT22), .Z(n454) );
  XNOR2_X1 U507 ( .A(G22GAT), .B(KEYINPUT23), .ZN(n453) );
  XNOR2_X1 U508 ( .A(n454), .B(n453), .ZN(n455) );
  XOR2_X1 U509 ( .A(n456), .B(n455), .Z(n457) );
  XNOR2_X1 U510 ( .A(n458), .B(n457), .ZN(n478) );
  NOR2_X1 U511 ( .A1(n573), .A2(n478), .ZN(n460) );
  XNOR2_X1 U512 ( .A(KEYINPUT55), .B(KEYINPUT119), .ZN(n459) );
  XNOR2_X1 U513 ( .A(n460), .B(n459), .ZN(n461) );
  NAND2_X1 U514 ( .A1(n570), .A2(n559), .ZN(n466) );
  XOR2_X1 U515 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n464) );
  XOR2_X1 U516 ( .A(G176GAT), .B(KEYINPUT121), .Z(n463) );
  XNOR2_X1 U517 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U518 ( .A(n466), .B(n465), .ZN(G1349GAT) );
  NAND2_X1 U519 ( .A1(n570), .A2(n582), .ZN(n468) );
  XNOR2_X1 U520 ( .A(G183GAT), .B(KEYINPUT122), .ZN(n467) );
  XNOR2_X1 U521 ( .A(n468), .B(n467), .ZN(G1350GAT) );
  NAND2_X1 U522 ( .A1(n566), .A2(n570), .ZN(n471) );
  XOR2_X1 U523 ( .A(KEYINPUT58), .B(KEYINPUT123), .Z(n469) );
  XOR2_X1 U524 ( .A(KEYINPUT102), .B(KEYINPUT34), .Z(n492) );
  NAND2_X1 U525 ( .A1(n578), .A2(n574), .ZN(n502) );
  XNOR2_X1 U526 ( .A(KEYINPUT28), .B(n478), .ZN(n533) );
  XOR2_X1 U527 ( .A(n528), .B(KEYINPUT27), .Z(n482) );
  NOR2_X1 U528 ( .A1(n533), .A2(n482), .ZN(n472) );
  NAND2_X1 U529 ( .A1(n555), .A2(n472), .ZN(n540) );
  XOR2_X1 U530 ( .A(KEYINPUT89), .B(n541), .Z(n473) );
  NOR2_X1 U531 ( .A1(n540), .A2(n473), .ZN(n487) );
  NOR2_X1 U532 ( .A1(n479), .A2(n474), .ZN(n475) );
  XOR2_X1 U533 ( .A(KEYINPUT101), .B(n475), .Z(n476) );
  NOR2_X1 U534 ( .A1(n478), .A2(n476), .ZN(n477) );
  XOR2_X1 U535 ( .A(KEYINPUT25), .B(n477), .Z(n484) );
  XOR2_X1 U536 ( .A(KEYINPUT26), .B(KEYINPUT99), .Z(n481) );
  NAND2_X1 U537 ( .A1(n479), .A2(n478), .ZN(n480) );
  XNOR2_X1 U538 ( .A(n481), .B(n480), .ZN(n572) );
  NOR2_X1 U539 ( .A1(n572), .A2(n482), .ZN(n554) );
  XNOR2_X1 U540 ( .A(n554), .B(KEYINPUT100), .ZN(n483) );
  NOR2_X1 U541 ( .A1(n484), .A2(n483), .ZN(n485) );
  NOR2_X1 U542 ( .A1(n555), .A2(n485), .ZN(n486) );
  NOR2_X1 U543 ( .A1(n487), .A2(n486), .ZN(n499) );
  XOR2_X1 U544 ( .A(KEYINPUT16), .B(KEYINPUT81), .Z(n489) );
  NAND2_X1 U545 ( .A1(n582), .A2(n551), .ZN(n488) );
  XNOR2_X1 U546 ( .A(n489), .B(n488), .ZN(n490) );
  OR2_X1 U547 ( .A1(n499), .A2(n490), .ZN(n515) );
  NOR2_X1 U548 ( .A1(n502), .A2(n515), .ZN(n497) );
  NAND2_X1 U549 ( .A1(n497), .A2(n555), .ZN(n491) );
  XNOR2_X1 U550 ( .A(n492), .B(n491), .ZN(n493) );
  XOR2_X1 U551 ( .A(G1GAT), .B(n493), .Z(G1324GAT) );
  NAND2_X1 U552 ( .A1(n528), .A2(n497), .ZN(n494) );
  XNOR2_X1 U553 ( .A(n494), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U554 ( .A(G15GAT), .B(KEYINPUT35), .Z(n496) );
  NAND2_X1 U555 ( .A1(n497), .A2(n541), .ZN(n495) );
  XNOR2_X1 U556 ( .A(n496), .B(n495), .ZN(G1326GAT) );
  NAND2_X1 U557 ( .A1(n497), .A2(n533), .ZN(n498) );
  XNOR2_X1 U558 ( .A(n498), .B(G22GAT), .ZN(G1327GAT) );
  NOR2_X1 U559 ( .A1(n587), .A2(n499), .ZN(n500) );
  NAND2_X1 U560 ( .A1(n500), .A2(n397), .ZN(n501) );
  XOR2_X1 U561 ( .A(KEYINPUT37), .B(n501), .Z(n526) );
  NOR2_X1 U562 ( .A1(n526), .A2(n502), .ZN(n503) );
  XNOR2_X1 U563 ( .A(KEYINPUT38), .B(n503), .ZN(n512) );
  NAND2_X1 U564 ( .A1(n555), .A2(n512), .ZN(n505) );
  XOR2_X1 U565 ( .A(G29GAT), .B(KEYINPUT39), .Z(n504) );
  XNOR2_X1 U566 ( .A(n505), .B(n504), .ZN(G1328GAT) );
  XNOR2_X1 U567 ( .A(G36GAT), .B(KEYINPUT104), .ZN(n507) );
  NAND2_X1 U568 ( .A1(n528), .A2(n512), .ZN(n506) );
  XNOR2_X1 U569 ( .A(n507), .B(n506), .ZN(G1329GAT) );
  XNOR2_X1 U570 ( .A(G43GAT), .B(KEYINPUT105), .ZN(n511) );
  XOR2_X1 U571 ( .A(KEYINPUT106), .B(KEYINPUT40), .Z(n509) );
  NAND2_X1 U572 ( .A1(n512), .A2(n541), .ZN(n508) );
  XNOR2_X1 U573 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U574 ( .A(n511), .B(n510), .ZN(G1330GAT) );
  XOR2_X1 U575 ( .A(G50GAT), .B(KEYINPUT107), .Z(n514) );
  NAND2_X1 U576 ( .A1(n533), .A2(n512), .ZN(n513) );
  XNOR2_X1 U577 ( .A(n514), .B(n513), .ZN(G1331GAT) );
  XOR2_X1 U578 ( .A(KEYINPUT108), .B(KEYINPUT42), .Z(n517) );
  NAND2_X1 U579 ( .A1(n543), .A2(n559), .ZN(n525) );
  NOR2_X1 U580 ( .A1(n525), .A2(n515), .ZN(n522) );
  NAND2_X1 U581 ( .A1(n522), .A2(n555), .ZN(n516) );
  XNOR2_X1 U582 ( .A(n517), .B(n516), .ZN(n518) );
  XOR2_X1 U583 ( .A(G57GAT), .B(n518), .Z(G1332GAT) );
  XOR2_X1 U584 ( .A(G64GAT), .B(KEYINPUT109), .Z(n520) );
  NAND2_X1 U585 ( .A1(n522), .A2(n528), .ZN(n519) );
  XNOR2_X1 U586 ( .A(n520), .B(n519), .ZN(G1333GAT) );
  NAND2_X1 U587 ( .A1(n541), .A2(n522), .ZN(n521) );
  XNOR2_X1 U588 ( .A(n521), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U589 ( .A(G78GAT), .B(KEYINPUT43), .Z(n524) );
  NAND2_X1 U590 ( .A1(n522), .A2(n533), .ZN(n523) );
  XNOR2_X1 U591 ( .A(n524), .B(n523), .ZN(G1335GAT) );
  NOR2_X1 U592 ( .A1(n526), .A2(n525), .ZN(n534) );
  NAND2_X1 U593 ( .A1(n555), .A2(n534), .ZN(n527) );
  XNOR2_X1 U594 ( .A(G85GAT), .B(n527), .ZN(G1336GAT) );
  XOR2_X1 U595 ( .A(KEYINPUT110), .B(KEYINPUT111), .Z(n530) );
  NAND2_X1 U596 ( .A1(n534), .A2(n528), .ZN(n529) );
  XNOR2_X1 U597 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U598 ( .A(G92GAT), .B(n531), .ZN(G1337GAT) );
  NAND2_X1 U599 ( .A1(n541), .A2(n534), .ZN(n532) );
  XNOR2_X1 U600 ( .A(n532), .B(G99GAT), .ZN(G1338GAT) );
  XNOR2_X1 U601 ( .A(G106GAT), .B(KEYINPUT112), .ZN(n538) );
  XOR2_X1 U602 ( .A(KEYINPUT113), .B(KEYINPUT44), .Z(n536) );
  NAND2_X1 U603 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U604 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U605 ( .A(n538), .B(n537), .ZN(G1339GAT) );
  NOR2_X1 U606 ( .A1(n539), .A2(n540), .ZN(n542) );
  NAND2_X1 U607 ( .A1(n542), .A2(n541), .ZN(n550) );
  NOR2_X1 U608 ( .A1(n543), .A2(n550), .ZN(n544) );
  XOR2_X1 U609 ( .A(G113GAT), .B(n544), .Z(G1340GAT) );
  INV_X1 U610 ( .A(n559), .ZN(n545) );
  NOR2_X1 U611 ( .A1(n545), .A2(n550), .ZN(n547) );
  XNOR2_X1 U612 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n547), .B(n546), .ZN(G1341GAT) );
  NOR2_X1 U614 ( .A1(n397), .A2(n550), .ZN(n548) );
  XOR2_X1 U615 ( .A(KEYINPUT50), .B(n548), .Z(n549) );
  XNOR2_X1 U616 ( .A(G127GAT), .B(n549), .ZN(G1342GAT) );
  NOR2_X1 U617 ( .A1(n551), .A2(n550), .ZN(n553) );
  XNOR2_X1 U618 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n553), .B(n552), .ZN(G1343GAT) );
  NAND2_X1 U620 ( .A1(n555), .A2(n554), .ZN(n556) );
  NOR2_X1 U621 ( .A1(n539), .A2(n556), .ZN(n557) );
  XOR2_X1 U622 ( .A(KEYINPUT115), .B(n557), .Z(n567) );
  NAND2_X1 U623 ( .A1(n574), .A2(n567), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n558), .B(G141GAT), .ZN(G1344GAT) );
  XNOR2_X1 U625 ( .A(G148GAT), .B(KEYINPUT116), .ZN(n563) );
  XOR2_X1 U626 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n561) );
  NAND2_X1 U627 ( .A1(n567), .A2(n559), .ZN(n560) );
  XNOR2_X1 U628 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(G1345GAT) );
  XOR2_X1 U630 ( .A(G155GAT), .B(KEYINPUT117), .Z(n565) );
  NAND2_X1 U631 ( .A1(n567), .A2(n582), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n565), .B(n564), .ZN(G1346GAT) );
  NAND2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n568), .B(KEYINPUT118), .ZN(n569) );
  XNOR2_X1 U635 ( .A(G162GAT), .B(n569), .ZN(G1347GAT) );
  NAND2_X1 U636 ( .A1(n570), .A2(n574), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n571), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n576) );
  NOR2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n583) );
  NAND2_X1 U640 ( .A1(n583), .A2(n574), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(n577), .ZN(G1352GAT) );
  XOR2_X1 U643 ( .A(KEYINPUT61), .B(KEYINPUT124), .Z(n580) );
  INV_X1 U644 ( .A(n583), .ZN(n586) );
  OR2_X1 U645 ( .A1(n586), .A2(n578), .ZN(n579) );
  XNOR2_X1 U646 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U647 ( .A(G204GAT), .B(n581), .ZN(G1353GAT) );
  XOR2_X1 U648 ( .A(G211GAT), .B(KEYINPUT125), .Z(n585) );
  NAND2_X1 U649 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n585), .B(n584), .ZN(G1354GAT) );
  NOR2_X1 U651 ( .A1(n587), .A2(n586), .ZN(n589) );
  XNOR2_X1 U652 ( .A(KEYINPUT62), .B(KEYINPUT126), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n589), .B(n588), .ZN(n590) );
  XOR2_X1 U654 ( .A(G218GAT), .B(n590), .Z(G1355GAT) );
endmodule

