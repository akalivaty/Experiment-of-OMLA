//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 1 0 0 1 0 1 0 0 1 0 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 0 1 1 0 0 1 1 1 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:18 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1294, new_n1295, new_n1296,
    new_n1297, new_n1298, new_n1299, new_n1300, new_n1302, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(G353));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n211));
  INV_X1    g0011(.A(G77), .ZN(new_n212));
  INV_X1    g0012(.A(G244), .ZN(new_n213));
  INV_X1    g0013(.A(G264), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n211), .B1(new_n212), .B2(new_n213), .C1(new_n207), .C2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n210), .B1(new_n215), .B2(new_n218), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT1), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n210), .A2(G13), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n221), .B(G250), .C1(G257), .C2(G264), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  XNOR2_X1  g0023(.A(KEYINPUT65), .B(KEYINPUT0), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  INV_X1    g0025(.A(G20), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(new_n201), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n228), .A2(G50), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  AOI22_X1  g0030(.A1(new_n223), .A2(new_n224), .B1(new_n227), .B2(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n231), .B1(new_n223), .B2(new_n224), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n220), .A2(new_n232), .ZN(G361));
  XOR2_X1   g0033(.A(G238), .B(G244), .Z(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G226), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G264), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G358));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n243), .B(new_n244), .Z(new_n245));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  XNOR2_X1  g0049(.A(KEYINPUT3), .B(G33), .ZN(new_n250));
  INV_X1    g0050(.A(G1698), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n250), .A2(G222), .A3(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n250), .A2(G1698), .ZN(new_n253));
  INV_X1    g0053(.A(G223), .ZN(new_n254));
  OAI221_X1 g0054(.A(new_n252), .B1(new_n212), .B2(new_n250), .C1(new_n253), .C2(new_n254), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n225), .B1(G33), .B2(G41), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT68), .ZN(new_n258));
  INV_X1    g0058(.A(G1), .ZN(new_n259));
  INV_X1    g0059(.A(G41), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(KEYINPUT67), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT67), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G41), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  OAI211_X1 g0064(.A(new_n258), .B(new_n259), .C1(new_n264), .C2(G45), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n259), .A2(G45), .ZN(new_n266));
  XNOR2_X1  g0066(.A(KEYINPUT67), .B(G41), .ZN(new_n267));
  OAI211_X1 g0067(.A(KEYINPUT68), .B(new_n266), .C1(new_n267), .C2(G1), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G274), .ZN(new_n270));
  AND2_X1   g0070(.A1(G1), .A2(G13), .ZN(new_n271));
  NAND2_X1  g0071(.A1(G33), .A2(G41), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n270), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n269), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n271), .A2(new_n272), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n259), .B1(G41), .B2(G45), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G226), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n257), .A2(new_n274), .A3(new_n279), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n280), .A2(KEYINPUT69), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n280), .A2(KEYINPUT69), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G190), .ZN(new_n285));
  INV_X1    g0085(.A(new_n283), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n286), .A2(new_n281), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G200), .ZN(new_n288));
  NOR2_X1   g0088(.A1(G20), .A2(G33), .ZN(new_n289));
  AOI22_X1  g0089(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n289), .ZN(new_n290));
  NOR2_X1   g0090(.A1(KEYINPUT8), .A2(G58), .ZN(new_n291));
  XNOR2_X1  g0091(.A(KEYINPUT70), .B(G58), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n291), .B1(new_n292), .B2(KEYINPUT8), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n226), .A2(G33), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n290), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(new_n225), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(KEYINPUT71), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT71), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n296), .A2(new_n301), .A3(new_n298), .ZN(new_n302));
  INV_X1    g0102(.A(G13), .ZN(new_n303));
  NOR3_X1   g0103(.A1(new_n303), .A2(new_n226), .A3(G1), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n304), .A2(new_n298), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n202), .B1(new_n259), .B2(G20), .ZN(new_n306));
  AOI22_X1  g0106(.A1(new_n305), .A2(new_n306), .B1(new_n202), .B2(new_n304), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n300), .A2(new_n302), .A3(new_n307), .ZN(new_n308));
  XNOR2_X1  g0108(.A(new_n308), .B(KEYINPUT9), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n285), .A2(new_n288), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(KEYINPUT10), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT10), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n285), .A2(new_n288), .A3(new_n309), .A4(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n308), .B1(new_n287), .B2(G179), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n284), .A2(G169), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n314), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT76), .ZN(new_n320));
  INV_X1    g0120(.A(G232), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n320), .B1(new_n277), .B2(new_n321), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n275), .A2(KEYINPUT76), .A3(G232), .A4(new_n276), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(G33), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(KEYINPUT3), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT3), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(G33), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n326), .A2(new_n328), .A3(G226), .A4(G1698), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n326), .A2(new_n328), .A3(G223), .A4(new_n251), .ZN(new_n330));
  INV_X1    g0130(.A(G87), .ZN(new_n331));
  OAI211_X1 g0131(.A(new_n329), .B(new_n330), .C1(new_n325), .C2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(new_n256), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n324), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n273), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n335), .B1(new_n265), .B2(new_n268), .ZN(new_n336));
  OAI21_X1  g0136(.A(G169), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  AOI22_X1  g0137(.A1(new_n322), .A2(new_n323), .B1(new_n332), .B2(new_n256), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n338), .A2(G179), .A3(new_n274), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n292), .A2(G68), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n228), .ZN(new_n341));
  AOI22_X1  g0141(.A1(new_n341), .A2(G20), .B1(G159), .B2(new_n289), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT7), .ZN(new_n343));
  NOR3_X1   g0143(.A1(new_n250), .A2(new_n343), .A3(G20), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n327), .A2(G33), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n325), .A2(KEYINPUT3), .ZN(new_n346));
  OAI21_X1  g0146(.A(KEYINPUT74), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT74), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n326), .A2(new_n328), .A3(new_n348), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n347), .A2(new_n226), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n344), .B1(new_n350), .B2(new_n343), .ZN(new_n351));
  INV_X1    g0151(.A(G68), .ZN(new_n352));
  OAI211_X1 g0152(.A(KEYINPUT16), .B(new_n342), .C1(new_n351), .C2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT16), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n201), .B1(new_n292), .B2(G68), .ZN(new_n355));
  INV_X1    g0155(.A(G159), .ZN(new_n356));
  INV_X1    g0156(.A(new_n289), .ZN(new_n357));
  OAI22_X1  g0157(.A1(new_n355), .A2(new_n226), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n343), .B1(new_n250), .B2(G20), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n326), .A2(new_n328), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n360), .A2(KEYINPUT7), .A3(new_n226), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n352), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n354), .B1(new_n358), .B2(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n353), .A2(new_n298), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n259), .A2(G20), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n293), .A2(new_n365), .ZN(new_n366));
  OR2_X1    g0166(.A1(new_n366), .A2(KEYINPUT75), .ZN(new_n367));
  INV_X1    g0167(.A(new_n305), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n368), .B1(new_n366), .B2(KEYINPUT75), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n367), .A2(new_n369), .B1(new_n304), .B2(new_n294), .ZN(new_n370));
  AOI221_X4 g0170(.A(KEYINPUT18), .B1(new_n337), .B2(new_n339), .C1(new_n364), .C2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT18), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n364), .A2(new_n370), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n337), .A2(new_n339), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n372), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n371), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(G200), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n377), .B1(new_n334), .B2(new_n336), .ZN(new_n378));
  INV_X1    g0178(.A(G190), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n338), .A2(new_n379), .A3(new_n274), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  XOR2_X1   g0181(.A(KEYINPUT77), .B(KEYINPUT17), .Z(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n381), .A2(new_n364), .A3(new_n370), .A4(new_n383), .ZN(new_n384));
  AND3_X1   g0184(.A1(new_n381), .A2(new_n364), .A3(new_n370), .ZN(new_n385));
  NOR2_X1   g0185(.A1(KEYINPUT77), .A2(KEYINPUT17), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n384), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n305), .A2(G77), .A3(new_n365), .ZN(new_n388));
  XNOR2_X1  g0188(.A(new_n388), .B(KEYINPUT73), .ZN(new_n389));
  XOR2_X1   g0189(.A(KEYINPUT8), .B(G58), .Z(new_n390));
  OR2_X1    g0190(.A1(new_n289), .A2(KEYINPUT72), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n289), .A2(KEYINPUT72), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  XNOR2_X1  g0193(.A(KEYINPUT15), .B(G87), .ZN(new_n394));
  OAI221_X1 g0194(.A(new_n393), .B1(new_n226), .B2(new_n212), .C1(new_n295), .C2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(new_n298), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n304), .A2(new_n212), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n389), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(G238), .ZN(new_n399));
  OAI22_X1  g0199(.A1(new_n253), .A2(new_n399), .B1(new_n207), .B2(new_n250), .ZN(new_n400));
  NOR3_X1   g0200(.A1(new_n360), .A2(new_n321), .A3(G1698), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n256), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n278), .A2(G244), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n402), .A2(new_n274), .A3(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n398), .B1(G190), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n404), .A2(G200), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(G169), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n404), .A2(new_n409), .ZN(new_n410));
  AND2_X1   g0210(.A1(new_n398), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(G179), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n405), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n376), .A2(new_n387), .A3(new_n408), .A4(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n304), .A2(new_n352), .ZN(new_n416));
  XNOR2_X1  g0216(.A(new_n416), .B(KEYINPUT12), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n305), .A2(G68), .A3(new_n365), .ZN(new_n418));
  OAI22_X1  g0218(.A1(new_n357), .A2(new_n202), .B1(new_n226), .B2(G68), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n295), .A2(new_n212), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n298), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT11), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n417), .B(new_n418), .C1(new_n421), .C2(new_n422), .ZN(new_n423));
  AND2_X1   g0223(.A1(new_n421), .A2(new_n422), .ZN(new_n424));
  OR2_X1    g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT14), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n277), .A2(new_n399), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n427), .B1(new_n269), .B2(new_n273), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT13), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n250), .A2(G232), .A3(G1698), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n250), .A2(G226), .A3(new_n251), .ZN(new_n431));
  NAND2_X1  g0231(.A1(G33), .A2(G97), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n430), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(new_n256), .ZN(new_n434));
  AND3_X1   g0234(.A1(new_n428), .A2(new_n429), .A3(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n429), .B1(new_n428), .B2(new_n434), .ZN(new_n436));
  OAI211_X1 g0236(.A(new_n426), .B(G169), .C1(new_n435), .C2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n427), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n274), .A2(new_n434), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(KEYINPUT13), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n428), .A2(new_n429), .A3(new_n434), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n440), .A2(G179), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n437), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n440), .A2(new_n441), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n426), .B1(new_n444), .B2(G169), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n425), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n444), .A2(G200), .ZN(new_n447));
  INV_X1    g0247(.A(new_n425), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n447), .B(new_n448), .C1(new_n379), .C2(new_n444), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  NOR3_X1   g0250(.A1(new_n319), .A2(new_n415), .A3(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT89), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n250), .A2(G257), .A3(new_n251), .ZN(new_n453));
  XNOR2_X1  g0253(.A(KEYINPUT86), .B(G303), .ZN(new_n454));
  OAI221_X1 g0254(.A(new_n453), .B1(new_n250), .B2(new_n454), .C1(new_n253), .C2(new_n214), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(new_n256), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(KEYINPUT5), .B1(new_n261), .B2(new_n263), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT5), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n259), .B(G45), .C1(new_n459), .C2(G41), .ZN(new_n460));
  OAI211_X1 g0260(.A(G270), .B(new_n275), .C1(new_n458), .C2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT84), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n459), .A2(G41), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n464), .A2(new_n266), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n465), .B1(KEYINPUT5), .B2(new_n267), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n466), .A2(KEYINPUT84), .A3(G270), .A4(new_n275), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n465), .B(new_n273), .C1(KEYINPUT5), .C2(new_n267), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n463), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(KEYINPUT85), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT85), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n463), .A2(new_n467), .A3(new_n471), .A4(new_n468), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n457), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n303), .A2(G1), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(G20), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n259), .A2(G33), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n475), .A2(new_n476), .A3(new_n225), .A4(new_n297), .ZN(new_n477));
  INV_X1    g0277(.A(G116), .ZN(new_n478));
  OR3_X1    g0278(.A1(new_n477), .A2(KEYINPUT87), .A3(new_n478), .ZN(new_n479));
  OAI21_X1  g0279(.A(KEYINPUT87), .B1(new_n477), .B2(new_n478), .ZN(new_n480));
  AND2_X1   g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(G33), .A2(G283), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n482), .B(new_n226), .C1(G33), .C2(new_n206), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n483), .B(new_n298), .C1(new_n226), .C2(G116), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT20), .ZN(new_n485));
  XNOR2_X1  g0285(.A(new_n484), .B(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n474), .A2(G20), .A3(new_n478), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g0288(.A(G169), .B1(new_n481), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n452), .B1(new_n473), .B2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT21), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n452), .B(KEYINPUT21), .C1(new_n473), .C2(new_n489), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n479), .A2(new_n480), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n495), .A2(new_n487), .A3(new_n486), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n412), .B1(new_n455), .B2(new_n256), .ZN(new_n497));
  INV_X1    g0297(.A(new_n468), .ZN(new_n498));
  INV_X1    g0298(.A(new_n461), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n498), .B1(new_n499), .B2(KEYINPUT84), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n471), .B1(new_n500), .B2(new_n463), .ZN(new_n501));
  INV_X1    g0301(.A(new_n472), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n496), .B(new_n497), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT88), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n456), .A2(G179), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n506), .B1(new_n470), .B2(new_n472), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n507), .A2(KEYINPUT88), .A3(new_n496), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n470), .A2(new_n472), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n456), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(G200), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n496), .B1(new_n473), .B2(G190), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT90), .ZN(new_n515));
  AND3_X1   g0315(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n515), .B1(new_n513), .B2(new_n514), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n494), .B(new_n510), .C1(new_n516), .C2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n326), .A2(new_n328), .A3(G257), .A4(G1698), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n326), .A2(new_n328), .A3(G250), .A4(new_n251), .ZN(new_n521));
  NAND2_X1  g0321(.A1(G33), .A2(G294), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n523), .A2(KEYINPUT91), .A3(new_n256), .ZN(new_n524));
  OAI211_X1 g0324(.A(G264), .B(new_n275), .C1(new_n458), .C2(new_n460), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n524), .A2(new_n468), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g0326(.A(KEYINPUT91), .B1(new_n523), .B2(new_n256), .ZN(new_n527));
  OAI21_X1  g0327(.A(G169), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n523), .A2(new_n256), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n529), .A2(G179), .A3(new_n468), .A4(new_n525), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n326), .A2(new_n328), .A3(new_n226), .A4(G87), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(KEYINPUT22), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT22), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n250), .A2(new_n534), .A3(new_n226), .A4(G87), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT24), .ZN(new_n537));
  NAND2_X1  g0337(.A1(G33), .A2(G116), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n538), .A2(G20), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT23), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n540), .B1(new_n226), .B2(G107), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n207), .A2(KEYINPUT23), .A3(G20), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n539), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  AND3_X1   g0343(.A1(new_n536), .A2(new_n537), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n537), .B1(new_n536), .B2(new_n543), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n298), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(new_n477), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT25), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(new_n475), .B2(G107), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n304), .A2(KEYINPUT25), .A3(new_n207), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n547), .A2(G107), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n546), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n531), .A2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT91), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n529), .A2(new_n554), .ZN(new_n555));
  AND2_X1   g0355(.A1(new_n525), .A2(new_n468), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n555), .A2(new_n556), .A3(new_n379), .A4(new_n524), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n529), .A2(new_n468), .A3(new_n525), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n377), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n560), .A2(new_n546), .A3(new_n551), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n553), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(KEYINPUT92), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT83), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n304), .A2(new_n206), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n565), .B1(new_n477), .B2(new_n206), .ZN(new_n566));
  XNOR2_X1  g0366(.A(G97), .B(G107), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT6), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NOR3_X1   g0369(.A1(new_n568), .A2(new_n206), .A3(G107), .ZN(new_n570));
  INV_X1    g0370(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n572), .A2(G20), .B1(G77), .B2(new_n289), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n359), .A2(new_n361), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(G107), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n566), .B1(new_n576), .B2(new_n298), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n326), .A2(new_n328), .A3(G244), .A4(new_n251), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT4), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n250), .A2(KEYINPUT4), .A3(G244), .A4(new_n251), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n250), .A2(G250), .A3(G1698), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n580), .A2(new_n581), .A3(new_n482), .A4(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n256), .ZN(new_n584));
  OAI211_X1 g0384(.A(G257), .B(new_n275), .C1(new_n458), .C2(new_n460), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n468), .ZN(new_n586));
  INV_X1    g0386(.A(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n584), .A2(new_n587), .A3(G190), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT78), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n585), .A2(KEYINPUT78), .A3(new_n468), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n590), .A2(new_n591), .B1(new_n256), .B2(new_n583), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n577), .B(new_n588), .C1(new_n592), .C2(new_n377), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n584), .A2(new_n587), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n409), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n570), .B1(new_n568), .B2(new_n567), .ZN(new_n596));
  OAI22_X1  g0396(.A1(new_n596), .A2(new_n226), .B1(new_n212), .B2(new_n357), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n207), .B1(new_n359), .B2(new_n361), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n298), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n547), .A2(G97), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n599), .A2(new_n565), .A3(new_n600), .ZN(new_n601));
  AND3_X1   g0401(.A1(new_n585), .A2(KEYINPUT78), .A3(new_n468), .ZN(new_n602));
  AOI21_X1  g0402(.A(KEYINPUT78), .B1(new_n585), .B2(new_n468), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n412), .B(new_n584), .C1(new_n602), .C2(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n595), .A2(new_n601), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n593), .A2(new_n605), .ZN(new_n606));
  NOR3_X1   g0406(.A1(new_n360), .A2(new_n213), .A3(new_n251), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n326), .A2(new_n328), .A3(G238), .A4(new_n251), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n538), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n256), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT79), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n266), .A2(G250), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n611), .B1(new_n256), .B2(new_n612), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n275), .A2(KEYINPUT79), .A3(G250), .A4(new_n266), .ZN(new_n614));
  INV_X1    g0414(.A(new_n266), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n613), .A2(new_n614), .B1(new_n273), .B2(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n610), .A2(new_n616), .A3(G179), .ZN(new_n617));
  AND2_X1   g0417(.A1(new_n610), .A2(new_n616), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n617), .B1(new_n618), .B2(new_n409), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT19), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(KEYINPUT80), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT80), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(KEYINPUT19), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n432), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  OAI22_X1  g0424(.A1(new_n624), .A2(G20), .B1(G87), .B2(new_n208), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n226), .A2(G33), .A3(G97), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT81), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n626), .A2(new_n621), .A3(new_n623), .A4(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n250), .A2(new_n226), .A3(G68), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n626), .A2(new_n621), .A3(new_n623), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(KEYINPUT81), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n625), .A2(new_n628), .A3(new_n629), .A4(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n298), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n394), .A2(new_n304), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT82), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n635), .B1(new_n477), .B2(new_n394), .ZN(new_n636));
  INV_X1    g0436(.A(new_n394), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n305), .A2(KEYINPUT82), .A3(new_n637), .A4(new_n476), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n633), .A2(new_n634), .A3(new_n636), .A4(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n619), .A2(new_n639), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n377), .B1(new_n610), .B2(new_n616), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n632), .A2(new_n298), .B1(new_n304), .B2(new_n394), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n547), .A2(G87), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n610), .A2(new_n616), .A3(G190), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n642), .A2(new_n643), .A3(new_n644), .A4(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n640), .A2(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n564), .B1(new_n606), .B2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT92), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n553), .A2(new_n561), .A3(new_n649), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n643), .A2(new_n644), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n641), .B1(G190), .B2(new_n618), .ZN(new_n652));
  AOI22_X1  g0452(.A1(new_n651), .A2(new_n652), .B1(new_n619), .B2(new_n639), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n653), .A2(KEYINPUT83), .A3(new_n593), .A4(new_n605), .ZN(new_n654));
  AND4_X1   g0454(.A1(new_n563), .A2(new_n648), .A3(new_n650), .A4(new_n654), .ZN(new_n655));
  AND3_X1   g0455(.A1(new_n451), .A2(new_n519), .A3(new_n655), .ZN(G372));
  INV_X1    g0456(.A(new_n414), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n449), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n446), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n387), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n373), .A2(new_n374), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(KEYINPUT18), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n373), .A2(new_n372), .A3(new_n374), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n662), .A2(KEYINPUT93), .A3(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT93), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n665), .B1(new_n371), .B2(new_n375), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n660), .A2(new_n667), .ZN(new_n668));
  OR2_X1    g0468(.A1(new_n668), .A2(KEYINPUT94), .ZN(new_n669));
  AOI22_X1  g0469(.A1(new_n668), .A2(KEYINPUT94), .B1(new_n311), .B2(new_n313), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n317), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n451), .ZN(new_n672));
  INV_X1    g0472(.A(new_n605), .ZN(new_n673));
  AND3_X1   g0473(.A1(new_n653), .A2(KEYINPUT26), .A3(new_n673), .ZN(new_n674));
  AOI21_X1  g0474(.A(KEYINPUT26), .B1(new_n653), .B2(new_n673), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n640), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n494), .A2(new_n510), .A3(new_n553), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n606), .A2(new_n647), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(new_n561), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n676), .B1(new_n677), .B2(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n671), .B1(new_n672), .B2(new_n681), .ZN(new_n682));
  XOR2_X1   g0482(.A(new_n682), .B(KEYINPUT95), .Z(G369));
  INV_X1    g0483(.A(G330), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n474), .A2(new_n226), .ZN(new_n685));
  OR2_X1    g0485(.A1(new_n685), .A2(KEYINPUT27), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(KEYINPUT27), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n686), .A2(G213), .A3(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(G343), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n496), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g0491(.A(new_n691), .B(KEYINPUT96), .Z(new_n692));
  NAND2_X1  g0492(.A1(new_n519), .A2(new_n692), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n509), .B1(new_n492), .B2(new_n493), .ZN(new_n694));
  OR2_X1    g0494(.A1(new_n694), .A2(new_n692), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n684), .B1(new_n693), .B2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  AND3_X1   g0497(.A1(new_n553), .A2(new_n649), .A3(new_n561), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n649), .B1(new_n553), .B2(new_n561), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n552), .A2(new_n690), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n690), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n553), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n702), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT97), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n702), .A2(KEYINPUT97), .A3(new_n705), .ZN(new_n709));
  AND2_X1   g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n697), .A2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n694), .A2(new_n690), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n714), .B1(new_n708), .B2(new_n709), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n553), .A2(new_n690), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n712), .A2(new_n717), .ZN(G399));
  INV_X1    g0518(.A(new_n221), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(new_n264), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n208), .A2(G87), .A3(G116), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n721), .A2(G1), .A3(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n723), .B1(new_n229), .B2(new_n721), .ZN(new_n724));
  XNOR2_X1  g0524(.A(new_n724), .B(KEYINPUT28), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT100), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT99), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n584), .B1(new_n602), .B2(new_n603), .ZN(new_n728));
  AOI21_X1  g0528(.A(G179), .B1(new_n610), .B2(new_n616), .ZN(new_n729));
  AND3_X1   g0529(.A1(new_n728), .A2(new_n558), .A3(new_n729), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n727), .B1(new_n512), .B2(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n728), .A2(new_n558), .A3(new_n729), .ZN(new_n732));
  NOR3_X1   g0532(.A1(new_n473), .A2(new_n732), .A3(KEYINPUT99), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n610), .A2(new_n616), .A3(new_n529), .A4(new_n525), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n594), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT30), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(KEYINPUT98), .ZN(new_n738));
  AND4_X1   g0538(.A1(new_n511), .A2(new_n736), .A3(new_n497), .A4(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n738), .B1(new_n507), .B2(new_n736), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n703), .B1(new_n734), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n726), .B1(new_n742), .B2(KEYINPUT31), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n511), .A2(new_n736), .A3(new_n497), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n744), .A2(KEYINPUT98), .A3(new_n737), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n512), .A2(new_n730), .A3(new_n727), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n507), .A2(new_n738), .A3(new_n736), .ZN(new_n747));
  OAI21_X1  g0547(.A(KEYINPUT99), .B1(new_n473), .B2(new_n732), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n745), .A2(new_n746), .A3(new_n747), .A4(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(KEYINPUT31), .B1(new_n749), .B2(new_n690), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(KEYINPUT100), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n743), .A2(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n741), .B1(new_n473), .B2(new_n732), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n753), .A2(KEYINPUT31), .A3(new_n690), .ZN(new_n754));
  NAND4_X1  g0554(.A1(new_n700), .A2(new_n648), .A3(new_n654), .A4(new_n703), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n754), .B1(new_n755), .B2(new_n518), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n752), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(new_n684), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n679), .B1(new_n694), .B2(new_n553), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n703), .B1(new_n759), .B2(new_n676), .ZN(new_n760));
  XNOR2_X1  g0560(.A(KEYINPUT101), .B(KEYINPUT29), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n760), .A2(KEYINPUT102), .A3(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n681), .A2(new_n690), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(KEYINPUT29), .ZN(new_n765));
  AND2_X1   g0565(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(KEYINPUT102), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n767), .B1(new_n764), .B2(new_n761), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n758), .B1(new_n766), .B2(new_n768), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n725), .B1(new_n769), .B2(G1), .ZN(G364));
  NOR2_X1   g0570(.A1(new_n303), .A2(G20), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n259), .B1(new_n771), .B2(G45), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n720), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n693), .A2(new_n684), .A3(new_n695), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n697), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(G13), .A2(G33), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(G20), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n693), .A2(new_n695), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n250), .A2(new_n221), .ZN(new_n782));
  INV_X1    g0582(.A(G355), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n782), .A2(new_n783), .B1(G116), .B2(new_n221), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n347), .A2(new_n349), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(new_n719), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(G45), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n787), .B1(new_n788), .B2(new_n230), .ZN(new_n789));
  OR2_X1    g0589(.A1(new_n245), .A2(new_n788), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n784), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n226), .B1(KEYINPUT103), .B2(new_n409), .ZN(new_n792));
  OR2_X1    g0592(.A1(new_n409), .A2(KEYINPUT103), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n225), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(new_n780), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n774), .B1(new_n791), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n226), .A2(new_n412), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(G200), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(G190), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  OR2_X1    g0601(.A1(KEYINPUT33), .A2(G317), .ZN(new_n802));
  NAND2_X1  g0602(.A1(KEYINPUT33), .A2(G317), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n801), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n799), .A2(new_n379), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(G326), .ZN(new_n807));
  INV_X1    g0607(.A(G294), .ZN(new_n808));
  NOR3_X1   g0608(.A1(new_n379), .A2(G179), .A3(G200), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n809), .A2(new_n226), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n806), .A2(new_n807), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n804), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n377), .A2(G179), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n813), .A2(G20), .A3(G190), .ZN(new_n814));
  INV_X1    g0614(.A(G303), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n360), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n798), .A2(G190), .A3(new_n377), .ZN(new_n817));
  INV_X1    g0617(.A(G322), .ZN(new_n818));
  NOR2_X1   g0618(.A1(G190), .A2(G200), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n798), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(G311), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n817), .A2(new_n818), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n379), .A2(G20), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT104), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n823), .B(new_n824), .ZN(new_n825));
  NOR3_X1   g0625(.A1(new_n825), .A2(G179), .A3(new_n377), .ZN(new_n826));
  AOI211_X1 g0626(.A(new_n816), .B(new_n822), .C1(new_n826), .C2(G283), .ZN(new_n827));
  NOR3_X1   g0627(.A1(new_n825), .A2(G179), .A3(G200), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  OR2_X1    g0629(.A1(new_n829), .A2(KEYINPUT107), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(KEYINPUT107), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(G329), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n812), .B(new_n827), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n292), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n835), .A2(new_n817), .B1(new_n820), .B2(new_n212), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n806), .A2(new_n202), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n836), .B(new_n837), .C1(G68), .C2(new_n800), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n250), .B1(new_n814), .B2(new_n331), .ZN(new_n839));
  OR2_X1    g0639(.A1(new_n839), .A2(KEYINPUT105), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n826), .A2(G107), .B1(new_n839), .B2(KEYINPUT105), .ZN(new_n841));
  XOR2_X1   g0641(.A(new_n810), .B(KEYINPUT106), .Z(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(G97), .ZN(new_n843));
  NAND4_X1  g0643(.A1(new_n838), .A2(new_n840), .A3(new_n841), .A4(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n828), .A2(G159), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n845), .B(KEYINPUT32), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n834), .B1(new_n844), .B2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT108), .ZN(new_n848));
  OR2_X1    g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n794), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n850), .B1(new_n847), .B2(new_n848), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n797), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n781), .A2(new_n852), .ZN(new_n853));
  AND2_X1   g0653(.A1(new_n777), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(G396));
  NAND2_X1  g0655(.A1(new_n398), .A2(new_n690), .ZN(new_n856));
  AOI22_X1  g0656(.A1(new_n408), .A2(new_n856), .B1(new_n411), .B2(new_n413), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n414), .A2(new_n690), .ZN(new_n858));
  OR2_X1    g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n760), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n857), .A2(new_n858), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n703), .B(new_n861), .C1(new_n759), .C2(new_n676), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n517), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n655), .A2(new_n694), .A3(new_n866), .A4(new_n703), .ZN(new_n867));
  NAND4_X1  g0667(.A1(new_n867), .A2(new_n754), .A3(new_n743), .A4(new_n751), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(G330), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n775), .B1(new_n863), .B2(new_n869), .ZN(new_n870));
  AND2_X1   g0670(.A1(new_n863), .A2(new_n869), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n870), .B1(KEYINPUT109), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n872), .B1(KEYINPUT109), .B2(new_n871), .ZN(new_n873));
  INV_X1    g0673(.A(new_n832), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(G311), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n826), .A2(G87), .ZN(new_n876));
  INV_X1    g0676(.A(G283), .ZN(new_n877));
  OAI22_X1  g0677(.A1(new_n877), .A2(new_n801), .B1(new_n806), .B2(new_n815), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n360), .B1(new_n817), .B2(new_n808), .ZN(new_n879));
  OAI22_X1  g0679(.A1(new_n207), .A2(new_n814), .B1(new_n820), .B2(new_n478), .ZN(new_n880));
  NOR3_X1   g0680(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  NAND4_X1  g0681(.A1(new_n875), .A2(new_n843), .A3(new_n876), .A4(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n874), .A2(G132), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n826), .A2(G68), .ZN(new_n884));
  INV_X1    g0684(.A(new_n810), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n292), .ZN(new_n886));
  INV_X1    g0686(.A(new_n785), .ZN(new_n887));
  INV_X1    g0687(.A(new_n814), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n887), .B1(G50), .B2(new_n888), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n883), .A2(new_n884), .A3(new_n886), .A4(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n817), .ZN(new_n891));
  INV_X1    g0691(.A(new_n820), .ZN(new_n892));
  AOI22_X1  g0692(.A1(new_n891), .A2(G143), .B1(new_n892), .B2(G159), .ZN(new_n893));
  INV_X1    g0693(.A(G137), .ZN(new_n894));
  INV_X1    g0694(.A(G150), .ZN(new_n895));
  OAI221_X1 g0695(.A(new_n893), .B1(new_n806), .B2(new_n894), .C1(new_n895), .C2(new_n801), .ZN(new_n896));
  XOR2_X1   g0696(.A(new_n896), .B(KEYINPUT34), .Z(new_n897));
  OAI21_X1  g0697(.A(new_n882), .B1(new_n890), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n794), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n794), .A2(new_n778), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n775), .B1(new_n900), .B2(new_n212), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n899), .B(new_n901), .C1(new_n861), .C2(new_n779), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n873), .A2(new_n902), .ZN(G384));
  INV_X1    g0703(.A(KEYINPUT40), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT38), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT37), .ZN(new_n906));
  INV_X1    g0706(.A(new_n688), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n373), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n381), .A2(new_n364), .A3(new_n370), .ZN(new_n909));
  AND4_X1   g0709(.A1(new_n906), .A2(new_n661), .A3(new_n908), .A4(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n353), .A2(new_n298), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n342), .B1(new_n351), .B2(new_n352), .ZN(new_n912));
  AOI21_X1  g0712(.A(KEYINPUT16), .B1(new_n912), .B2(KEYINPUT111), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT111), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n914), .B(new_n342), .C1(new_n351), .C2(new_n352), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n911), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(new_n370), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n907), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n374), .B1(new_n916), .B2(new_n917), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n918), .A2(new_n919), .A3(new_n909), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n910), .B1(KEYINPUT37), .B2(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n918), .B1(new_n376), .B2(new_n387), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n905), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n387), .A2(new_n662), .A3(new_n663), .ZN(new_n924));
  INV_X1    g0724(.A(new_n918), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n912), .A2(KEYINPUT111), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n927), .A2(new_n354), .A3(new_n915), .ZN(new_n928));
  INV_X1    g0728(.A(new_n911), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n370), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n385), .B1(new_n931), .B2(new_n374), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n906), .B1(new_n932), .B2(new_n918), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n926), .B(KEYINPUT38), .C1(new_n933), .C2(new_n910), .ZN(new_n934));
  AND2_X1   g0734(.A1(new_n923), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n425), .A2(new_n690), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n936), .B1(new_n446), .B2(new_n449), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n446), .A2(new_n449), .A3(new_n936), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n859), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n750), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n749), .A2(KEYINPUT31), .A3(new_n690), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n755), .A2(new_n518), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n940), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n904), .B1(new_n935), .B2(new_n945), .ZN(new_n946));
  AND3_X1   g0746(.A1(new_n446), .A2(new_n449), .A3(new_n936), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n861), .B1(new_n947), .B2(new_n937), .ZN(new_n948));
  INV_X1    g0748(.A(new_n942), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n949), .A2(new_n750), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n948), .B1(new_n867), .B2(new_n950), .ZN(new_n951));
  NOR3_X1   g0751(.A1(new_n371), .A2(new_n375), .A3(new_n665), .ZN(new_n952));
  AOI21_X1  g0752(.A(KEYINPUT93), .B1(new_n662), .B2(new_n663), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n387), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(new_n908), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n661), .A2(new_n908), .A3(new_n909), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(new_n906), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(KEYINPUT38), .B1(new_n956), .B2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n934), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n951), .B(KEYINPUT40), .C1(new_n960), .C2(new_n961), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n946), .A2(new_n962), .A3(G330), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n867), .A2(new_n950), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n451), .A2(G330), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  OR2_X1    g0766(.A1(new_n966), .A2(KEYINPUT112), .ZN(new_n967));
  NAND4_X1  g0767(.A1(new_n946), .A2(new_n962), .A3(new_n451), .A4(new_n964), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n966), .A2(KEYINPUT112), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n967), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n908), .B1(new_n667), .B2(new_n387), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n905), .B1(new_n971), .B2(new_n958), .ZN(new_n972));
  AOI21_X1  g0772(.A(KEYINPUT39), .B1(new_n972), .B2(new_n934), .ZN(new_n973));
  AND3_X1   g0773(.A1(new_n923), .A2(new_n934), .A3(KEYINPUT39), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n659), .A2(new_n703), .ZN(new_n975));
  NOR3_X1   g0775(.A1(new_n973), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n923), .A2(new_n934), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n947), .A2(new_n937), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  NOR3_X1   g0779(.A1(new_n681), .A2(new_n690), .A3(new_n859), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n977), .B(new_n979), .C1(new_n980), .C2(new_n858), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n664), .A2(new_n666), .A3(new_n688), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n976), .A2(new_n983), .ZN(new_n984));
  NAND4_X1  g0784(.A1(new_n768), .A2(new_n451), .A3(new_n765), .A4(new_n763), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(new_n671), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n984), .B(new_n986), .Z(new_n987));
  OAI22_X1  g0787(.A1(new_n970), .A2(new_n987), .B1(new_n259), .B2(new_n771), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n988), .A2(KEYINPUT113), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n970), .A2(new_n987), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n988), .A2(KEYINPUT113), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n989), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  OAI211_X1 g0792(.A(G116), .B(new_n227), .C1(new_n572), .C2(KEYINPUT35), .ZN(new_n993));
  AOI22_X1  g0793(.A1(new_n993), .A2(KEYINPUT110), .B1(KEYINPUT35), .B2(new_n572), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(KEYINPUT110), .B2(new_n993), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT36), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n230), .A2(new_n340), .A3(G77), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n997), .B1(G50), .B2(new_n352), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n998), .A2(G1), .A3(new_n303), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n992), .A2(new_n996), .A3(new_n999), .ZN(G367));
  OAI21_X1  g0800(.A(new_n653), .B1(new_n651), .B2(new_n703), .ZN(new_n1001));
  OR3_X1    g0801(.A1(new_n640), .A2(new_n651), .A3(new_n703), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT43), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1003), .A2(KEYINPUT43), .ZN(new_n1007));
  OAI211_X1 g0807(.A(new_n593), .B(new_n605), .C1(new_n577), .C2(new_n703), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n673), .A2(new_n690), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n715), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(KEYINPUT42), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT114), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n593), .A2(new_n531), .A3(new_n552), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n690), .B1(new_n1014), .B2(new_n605), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1015), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1012), .A2(new_n1013), .A3(new_n1016), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1011), .A2(KEYINPUT42), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1015), .B1(new_n1011), .B2(KEYINPUT42), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1021), .A2(new_n1013), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n1006), .B(new_n1007), .C1(new_n1020), .C2(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1010), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n712), .A2(new_n1024), .ZN(new_n1025));
  OR2_X1    g0825(.A1(new_n1021), .A2(new_n1013), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1018), .B1(new_n1021), .B2(new_n1013), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n1026), .A2(new_n1027), .A3(new_n1005), .A4(new_n1004), .ZN(new_n1028));
  AND3_X1   g0828(.A1(new_n1023), .A2(new_n1025), .A3(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1025), .B1(new_n1023), .B2(new_n1028), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n720), .B(KEYINPUT41), .Z(new_n1032));
  INV_X1    g0832(.A(KEYINPUT45), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n708), .A2(new_n709), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1034), .A2(new_n713), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n716), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1033), .B1(new_n1037), .B2(new_n1024), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n717), .A2(KEYINPUT45), .A3(new_n1010), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1037), .A2(KEYINPUT44), .A3(new_n1024), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT44), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n717), .B2(new_n1010), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1040), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT115), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1045), .A2(new_n1046), .A3(new_n711), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n769), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT116), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n697), .B(new_n1049), .C1(new_n1034), .C2(new_n713), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n1034), .A2(new_n713), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n696), .B1(new_n1051), .B2(KEYINPUT116), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1053), .A2(new_n1035), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1050), .A2(new_n1052), .A3(new_n715), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1048), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1040), .B(new_n1044), .C1(KEYINPUT115), .C2(new_n712), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1047), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1032), .B1(new_n1058), .B2(new_n769), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1031), .B1(new_n1059), .B2(new_n773), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n787), .A2(new_n241), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n795), .B1(new_n221), .B2(new_n394), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n774), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n826), .A2(G97), .ZN(new_n1064));
  INV_X1    g0864(.A(G317), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1064), .B1(new_n829), .B2(new_n1065), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n887), .B1(new_n877), .B2(new_n820), .C1(new_n454), .C2(new_n817), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n814), .A2(new_n478), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT46), .ZN(new_n1069));
  NOR3_X1   g0869(.A1(new_n1066), .A2(new_n1067), .A3(new_n1069), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(G107), .A2(new_n885), .B1(new_n805), .B2(G311), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1070), .B(new_n1071), .C1(new_n808), .C2(new_n801), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n842), .A2(G68), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n828), .A2(G137), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n835), .A2(new_n814), .B1(new_n817), .B2(new_n895), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1075), .B1(G50), .B2(new_n892), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n800), .A2(G159), .B1(new_n805), .B2(G143), .ZN(new_n1077));
  NAND4_X1  g0877(.A1(new_n1073), .A2(new_n1074), .A3(new_n1076), .A4(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n826), .A2(G77), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n250), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1080), .B(KEYINPUT117), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1072), .B1(new_n1078), .B2(new_n1081), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT47), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1063), .B1(new_n1083), .B2(new_n794), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n780), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1084), .B1(new_n1085), .B2(new_n1003), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1060), .A2(new_n1086), .ZN(G387));
  NOR2_X1   g0887(.A1(new_n1056), .A2(new_n721), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1088), .B1(new_n769), .B2(new_n1089), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n782), .A2(new_n722), .B1(G107), .B2(new_n221), .ZN(new_n1091));
  XOR2_X1   g0891(.A(new_n1091), .B(KEYINPUT118), .Z(new_n1092));
  AND2_X1   g0892(.A1(new_n238), .A2(G45), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n390), .A2(new_n202), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(KEYINPUT119), .B(KEYINPUT50), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1094), .B(new_n1095), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n722), .B(new_n788), .C1(new_n352), .C2(new_n212), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n786), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1092), .B1(new_n1093), .B2(new_n1098), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n1099), .A2(KEYINPUT120), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1099), .A2(KEYINPUT120), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n795), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n1064), .B1(new_n801), .B2(new_n294), .C1(new_n829), .C2(new_n895), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n842), .A2(new_n637), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(G77), .A2(new_n888), .B1(new_n892), .B2(G68), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1106), .B1(new_n202), .B2(new_n817), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n785), .B1(new_n806), .B2(new_n356), .ZN(new_n1108));
  NOR4_X1   g0908(.A1(new_n1103), .A2(new_n1105), .A3(new_n1107), .A4(new_n1108), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n810), .A2(new_n877), .B1(new_n814), .B2(new_n808), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n454), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n891), .A2(G317), .B1(new_n892), .B2(new_n1111), .ZN(new_n1112));
  OAI221_X1 g0912(.A(new_n1112), .B1(new_n806), .B2(new_n818), .C1(new_n821), .C2(new_n801), .ZN(new_n1113));
  INV_X1    g0913(.A(KEYINPUT48), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1110), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1115), .B1(new_n1114), .B2(new_n1113), .ZN(new_n1116));
  XOR2_X1   g0916(.A(new_n1116), .B(KEYINPUT121), .Z(new_n1117));
  OR2_X1    g0917(.A1(new_n1117), .A2(KEYINPUT49), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n826), .ZN(new_n1119));
  OAI221_X1 g0919(.A(new_n887), .B1(new_n829), .B2(new_n807), .C1(new_n478), .C2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1120), .B1(new_n1117), .B2(KEYINPUT49), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1109), .B1(new_n1118), .B2(new_n1121), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n774), .B1(new_n1100), .B2(new_n1102), .C1(new_n1122), .C2(new_n850), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1123), .B1(new_n710), .B2(new_n780), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1124), .B1(new_n1089), .B2(new_n773), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1090), .A2(new_n1125), .ZN(G393));
  XNOR2_X1  g0926(.A(new_n1045), .B(new_n712), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n1058), .B(new_n720), .C1(new_n1127), .C2(new_n1056), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n787), .A2(new_n248), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n795), .B1(new_n206), .B2(new_n221), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n876), .B(new_n785), .C1(new_n352), .C2(new_n814), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(G150), .A2(new_n805), .B1(new_n891), .B2(G159), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n1132), .B(KEYINPUT51), .ZN(new_n1133));
  AOI211_X1 g0933(.A(new_n1131), .B(new_n1133), .C1(G143), .C2(new_n828), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n842), .A2(G77), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n800), .A2(G50), .B1(new_n892), .B2(new_n390), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1135), .B1(KEYINPUT122), .B2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1137), .B1(KEYINPUT122), .B2(new_n1136), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n806), .A2(new_n1065), .B1(new_n821), .B2(new_n817), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n1139), .B(KEYINPUT52), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n207), .A2(new_n1119), .B1(new_n829), .B2(new_n818), .ZN(new_n1141));
  OAI221_X1 g0941(.A(new_n360), .B1(new_n820), .B2(new_n808), .C1(new_n877), .C2(new_n814), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n801), .A2(new_n454), .B1(new_n478), .B2(new_n810), .ZN(new_n1143));
  NOR3_X1   g0943(.A1(new_n1141), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n1134), .A2(new_n1138), .B1(new_n1140), .B2(new_n1144), .ZN(new_n1145));
  OAI221_X1 g0945(.A(new_n774), .B1(new_n1129), .B2(new_n1130), .C1(new_n1145), .C2(new_n850), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1146), .B1(new_n1024), .B2(new_n780), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1147), .B1(new_n1127), .B2(new_n773), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1128), .A2(new_n1148), .ZN(G390));
  INV_X1    g0949(.A(new_n858), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n978), .B1(new_n862), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n975), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n973), .A2(new_n974), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n979), .B1(new_n980), .B2(new_n858), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n972), .A2(new_n934), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1154), .A2(new_n975), .A3(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1153), .A2(new_n1156), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n859), .A2(new_n684), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n964), .A2(new_n979), .A3(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1157), .A2(new_n1160), .ZN(new_n1161));
  OAI211_X1 g0961(.A(G330), .B(new_n940), .C1(new_n752), .C2(new_n756), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(KEYINPUT123), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT123), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n868), .A2(new_n1164), .A3(G330), .A4(new_n940), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1153), .A2(new_n1166), .A3(new_n1156), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1161), .A2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n985), .A2(new_n671), .A3(new_n965), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n862), .A2(new_n1150), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n964), .A2(new_n1158), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1171), .B1(new_n1172), .B2(new_n978), .ZN(new_n1173));
  AND2_X1   g0973(.A1(new_n1166), .A2(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1171), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n978), .B1(new_n869), .B2(new_n859), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1175), .B1(new_n1176), .B2(new_n1159), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1170), .B1(new_n1174), .B2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n721), .B1(new_n1168), .B2(new_n1178), .ZN(new_n1179));
  AND3_X1   g0979(.A1(new_n1153), .A2(new_n1166), .A3(new_n1156), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1159), .B1(new_n1153), .B2(new_n1156), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1176), .A2(new_n1159), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1183), .A2(new_n1171), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1166), .A2(new_n1173), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1182), .A2(new_n1170), .A3(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1179), .A2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1161), .A2(new_n773), .A3(new_n1167), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n778), .B1(new_n973), .B2(new_n974), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n900), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n774), .B1(new_n1191), .B2(new_n293), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(KEYINPUT54), .B(G143), .ZN(new_n1193));
  INV_X1    g0993(.A(G132), .ZN(new_n1194));
  OAI221_X1 g0994(.A(new_n250), .B1(new_n820), .B2(new_n1193), .C1(new_n1194), .C2(new_n817), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n801), .A2(new_n894), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n1195), .B(new_n1196), .C1(G128), .C2(new_n805), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n842), .A2(G159), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT53), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1199), .B1(new_n814), .B2(new_n895), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n888), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n826), .A2(G50), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1197), .A2(new_n1198), .A3(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(G125), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n832), .A2(new_n1204), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n832), .A2(new_n808), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n207), .A2(new_n801), .B1(new_n806), .B2(new_n877), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n360), .B1(new_n814), .B2(new_n331), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n817), .A2(new_n478), .B1(new_n820), .B2(new_n206), .ZN(new_n1209));
  NOR3_X1   g1009(.A1(new_n1207), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1210), .A2(new_n884), .A3(new_n1135), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n1203), .A2(new_n1205), .B1(new_n1206), .B2(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1192), .B1(new_n1212), .B2(new_n794), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1190), .A2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1189), .A2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1188), .A2(new_n1216), .ZN(G378));
  XNOR2_X1  g1017(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n308), .A2(new_n907), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n314), .A2(new_n318), .A3(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1220), .B1(new_n314), .B2(new_n318), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1219), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1223), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1225), .A2(new_n1221), .A3(new_n1218), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1224), .A2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n963), .A2(new_n1228), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1227), .A2(new_n946), .A3(G330), .A4(new_n962), .ZN(new_n1230));
  AND3_X1   g1030(.A1(new_n1229), .A2(new_n984), .A3(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n984), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n773), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n774), .B1(new_n1191), .B2(G50), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(new_n887), .B2(new_n267), .ZN(new_n1236));
  OAI221_X1 g1036(.A(new_n887), .B1(new_n806), .B2(new_n478), .C1(new_n206), .C2(new_n801), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1119), .A2(new_n835), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n267), .B1(new_n814), .B2(new_n212), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n817), .A2(new_n207), .B1(new_n820), .B2(new_n394), .ZN(new_n1240));
  NOR4_X1   g1040(.A1(new_n1237), .A2(new_n1238), .A3(new_n1239), .A4(new_n1240), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1241), .B(new_n1073), .C1(new_n877), .C2(new_n832), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT58), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1236), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n1204), .A2(new_n806), .B1(new_n801), .B2(new_n1194), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n891), .A2(G128), .ZN(new_n1246));
  OAI221_X1 g1046(.A(new_n1246), .B1(new_n814), .B2(new_n1193), .C1(new_n894), .C2(new_n820), .ZN(new_n1247));
  AOI211_X1 g1047(.A(new_n1245), .B(new_n1247), .C1(G150), .C2(new_n842), .ZN(new_n1248));
  XNOR2_X1  g1048(.A(new_n1248), .B(KEYINPUT124), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1250), .A2(KEYINPUT59), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n325), .B(new_n260), .C1(new_n1119), .C2(new_n356), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1252), .B1(G124), .B2(new_n828), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT59), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1253), .B1(new_n1249), .B2(new_n1254), .ZN(new_n1255));
  OAI221_X1 g1055(.A(new_n1244), .B1(new_n1243), .B2(new_n1242), .C1(new_n1251), .C2(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1234), .B1(new_n1256), .B2(new_n794), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1257), .B1(new_n1227), .B2(new_n779), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1233), .A2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  OAI21_X1  g1060(.A(KEYINPUT57), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1169), .B1(new_n1182), .B2(new_n1186), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n720), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1170), .B1(new_n1168), .B2(new_n1178), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n984), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1229), .A2(new_n984), .A3(new_n1230), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(KEYINPUT57), .B1(new_n1264), .B2(new_n1269), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1260), .B1(new_n1263), .B2(new_n1270), .ZN(G375));
  NAND3_X1  g1071(.A1(new_n1184), .A2(new_n1169), .A3(new_n1185), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1032), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1272), .A2(new_n1178), .A3(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1186), .A2(new_n773), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n774), .B1(new_n1191), .B2(G68), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n874), .A2(G128), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n842), .A2(G50), .ZN(new_n1278));
  OAI22_X1  g1078(.A1(new_n356), .A2(new_n814), .B1(new_n820), .B2(new_n895), .ZN(new_n1279));
  AOI211_X1 g1079(.A(new_n1279), .B(new_n1238), .C1(G137), .C2(new_n891), .ZN(new_n1280));
  OAI221_X1 g1080(.A(new_n785), .B1(new_n806), .B2(new_n1194), .C1(new_n801), .C2(new_n1193), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1277), .A2(new_n1278), .A3(new_n1280), .A4(new_n1282), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n832), .A2(new_n815), .ZN(new_n1284));
  OAI22_X1  g1084(.A1(new_n478), .A2(new_n801), .B1(new_n806), .B2(new_n808), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n360), .B1(new_n817), .B2(new_n877), .ZN(new_n1286));
  OAI22_X1  g1086(.A1(new_n206), .A2(new_n814), .B1(new_n820), .B2(new_n207), .ZN(new_n1287));
  NOR3_X1   g1087(.A1(new_n1285), .A2(new_n1286), .A3(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1288), .A2(new_n1079), .A3(new_n1104), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1283), .B1(new_n1284), .B2(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1276), .B1(new_n1290), .B2(new_n794), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1291), .B1(new_n979), .B2(new_n779), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1274), .A2(new_n1275), .A3(new_n1292), .ZN(G381));
  NOR2_X1   g1093(.A1(G393), .A2(G396), .ZN(new_n1294));
  INV_X1    g1094(.A(G384), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  NOR3_X1   g1096(.A1(new_n1296), .A2(G390), .A3(G381), .ZN(new_n1297));
  INV_X1    g1097(.A(G387), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1215), .B1(new_n1179), .B2(new_n1187), .ZN(new_n1299));
  INV_X1    g1099(.A(G375), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1297), .A2(new_n1298), .A3(new_n1299), .A4(new_n1300), .ZN(G407));
  NAND2_X1  g1101(.A1(new_n1299), .A2(new_n689), .ZN(new_n1302));
  OAI211_X1 g1102(.A(G407), .B(G213), .C1(G375), .C2(new_n1302), .ZN(G409));
  OAI21_X1  g1103(.A(new_n1273), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1304));
  NOR2_X1   g1104(.A1(new_n1304), .A2(new_n1262), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1299), .B1(new_n1305), .B2(new_n1259), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT125), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  OAI211_X1 g1108(.A(G378), .B(new_n1260), .C1(new_n1263), .C2(new_n1270), .ZN(new_n1309));
  OAI211_X1 g1109(.A(new_n1299), .B(KEYINPUT125), .C1(new_n1305), .C2(new_n1259), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1308), .A2(new_n1309), .A3(new_n1310), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1184), .A2(new_n1185), .A3(KEYINPUT60), .A4(new_n1169), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1312), .A2(new_n720), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1178), .A2(KEYINPUT60), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1313), .B1(new_n1272), .B2(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1275), .A2(new_n1292), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1295), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1316), .ZN(new_n1318));
  AND2_X1   g1118(.A1(new_n1314), .A2(new_n1272), .ZN(new_n1319));
  OAI211_X1 g1119(.A(G384), .B(new_n1318), .C1(new_n1319), .C2(new_n1313), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1317), .A2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n689), .A2(G213), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1311), .A2(new_n1322), .A3(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1324), .A2(KEYINPUT62), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1311), .A2(new_n1323), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n689), .A2(G213), .A3(G2897), .ZN(new_n1327));
  AND3_X1   g1127(.A1(new_n1317), .A2(new_n1320), .A3(new_n1327), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1327), .B1(new_n1317), .B2(new_n1320), .ZN(new_n1329));
  NOR2_X1   g1129(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1326), .A2(new_n1330), .ZN(new_n1331));
  INV_X1    g1131(.A(KEYINPUT61), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT62), .ZN(new_n1333));
  NAND4_X1  g1133(.A1(new_n1311), .A2(new_n1333), .A3(new_n1322), .A4(new_n1323), .ZN(new_n1334));
  NAND4_X1  g1134(.A1(new_n1325), .A2(new_n1331), .A3(new_n1332), .A4(new_n1334), .ZN(new_n1335));
  AND3_X1   g1135(.A1(new_n1060), .A2(G390), .A3(new_n1086), .ZN(new_n1336));
  AOI21_X1  g1136(.A(G390), .B1(new_n1060), .B2(new_n1086), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n854), .B1(new_n1090), .B2(new_n1125), .ZN(new_n1338));
  OAI22_X1  g1138(.A1(new_n1336), .A2(new_n1337), .B1(new_n1294), .B2(new_n1338), .ZN(new_n1339));
  INV_X1    g1139(.A(G390), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(G387), .A2(new_n1340), .ZN(new_n1341));
  NOR2_X1   g1141(.A1(new_n1294), .A2(new_n1338), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1060), .A2(G390), .A3(new_n1086), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1341), .A2(new_n1342), .A3(new_n1343), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1339), .A2(new_n1344), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1335), .A2(new_n1345), .ZN(new_n1346));
  AND2_X1   g1146(.A1(new_n1339), .A2(new_n1344), .ZN(new_n1347));
  AOI21_X1  g1147(.A(KEYINPUT61), .B1(new_n1326), .B2(new_n1330), .ZN(new_n1348));
  INV_X1    g1148(.A(KEYINPUT63), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1324), .A2(new_n1349), .ZN(new_n1350));
  NAND4_X1  g1150(.A1(new_n1311), .A2(KEYINPUT63), .A3(new_n1322), .A4(new_n1323), .ZN(new_n1351));
  NAND4_X1  g1151(.A1(new_n1347), .A2(new_n1348), .A3(new_n1350), .A4(new_n1351), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1346), .A2(new_n1352), .ZN(G405));
  INV_X1    g1153(.A(KEYINPUT126), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1309), .A2(new_n1354), .ZN(new_n1355));
  NAND3_X1  g1155(.A1(new_n1322), .A2(new_n1299), .A3(G375), .ZN(new_n1356));
  OAI21_X1  g1156(.A(new_n1321), .B1(new_n1300), .B2(G378), .ZN(new_n1357));
  AOI21_X1  g1157(.A(new_n1355), .B1(new_n1356), .B2(new_n1357), .ZN(new_n1358));
  INV_X1    g1158(.A(new_n1358), .ZN(new_n1359));
  NAND3_X1  g1159(.A1(new_n1356), .A2(new_n1355), .A3(new_n1357), .ZN(new_n1360));
  NAND3_X1  g1160(.A1(new_n1347), .A2(new_n1359), .A3(new_n1360), .ZN(new_n1361));
  INV_X1    g1161(.A(new_n1360), .ZN(new_n1362));
  OAI21_X1  g1162(.A(new_n1345), .B1(new_n1362), .B2(new_n1358), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(new_n1361), .A2(new_n1363), .ZN(G402));
endmodule


