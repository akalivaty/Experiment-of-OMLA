

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821;

  AND2_X1 U370 ( .A1(n464), .A2(n417), .ZN(n380) );
  BUF_X1 U371 ( .A(n656), .Z(n491) );
  BUF_X1 U372 ( .A(G116), .Z(n433) );
  INV_X1 U373 ( .A(G101), .ZN(n595) );
  XNOR2_X1 U374 ( .A(KEYINPUT85), .B(KEYINPUT8), .ZN(n557) );
  XNOR2_X1 U375 ( .A(G119), .B(G116), .ZN(n436) );
  XOR2_X2 U376 ( .A(n552), .B(KEYINPUT21), .Z(n753) );
  AND2_X2 U377 ( .A1(n434), .A2(n524), .ZN(n523) );
  NOR2_X2 U378 ( .A1(n667), .A2(n531), .ZN(n520) );
  XNOR2_X2 U379 ( .A(KEYINPUT90), .B(KEYINPUT46), .ZN(n698) );
  XNOR2_X1 U380 ( .A(n347), .B(n409), .ZN(n422) );
  NAND2_X1 U381 ( .A1(n462), .A2(n463), .ZN(n347) );
  OR2_X2 U382 ( .A1(n794), .A2(n469), .ZN(n349) );
  NOR2_X1 U383 ( .A1(n348), .A2(n793), .ZN(G63) );
  XNOR2_X2 U384 ( .A(n787), .B(n788), .ZN(n348) );
  NOR2_X1 U385 ( .A1(n709), .A2(n781), .ZN(n437) );
  XNOR2_X1 U386 ( .A(G119), .B(G116), .ZN(n538) );
  XNOR2_X1 U387 ( .A(G119), .B(G137), .ZN(n533) );
  XNOR2_X1 U388 ( .A(G104), .B(G107), .ZN(n360) );
  NOR2_X1 U389 ( .A1(n640), .A2(n428), .ZN(n697) );
  BUF_X1 U390 ( .A(G122), .Z(n368) );
  NOR2_X2 U391 ( .A1(n754), .A2(n636), .ZN(n448) );
  AND2_X2 U392 ( .A1(n525), .A2(n527), .ZN(n485) );
  XNOR2_X1 U393 ( .A(KEYINPUT38), .B(n491), .ZN(n693) );
  NOR2_X1 U394 ( .A1(n699), .A2(n775), .ZN(n692) );
  XNOR2_X1 U395 ( .A(n400), .B(KEYINPUT22), .ZN(n634) );
  AND2_X1 U396 ( .A1(n387), .A2(KEYINPUT41), .ZN(n382) );
  NOR2_X1 U397 ( .A1(n745), .A2(n388), .ZN(n387) );
  AND2_X1 U398 ( .A1(n705), .A2(KEYINPUT64), .ZN(n359) );
  OR2_X1 U399 ( .A1(n705), .A2(KEYINPUT64), .ZN(n358) );
  NAND2_X1 U400 ( .A1(G214), .A2(n584), .ZN(n742) );
  INV_X1 U401 ( .A(G146), .ZN(n486) );
  INV_X1 U402 ( .A(G472), .ZN(n367) );
  INV_X1 U403 ( .A(KEYINPUT45), .ZN(n505) );
  INV_X1 U404 ( .A(KEYINPUT66), .ZN(n403) );
  INV_X1 U405 ( .A(KEYINPUT41), .ZN(n389) );
  AND2_X1 U406 ( .A1(n413), .A2(n378), .ZN(n376) );
  NAND2_X1 U407 ( .A1(n391), .A2(n396), .ZN(n390) );
  NAND2_X1 U408 ( .A1(n380), .A2(n419), .ZN(n375) );
  NAND2_X1 U409 ( .A1(n460), .A2(n406), .ZN(n459) );
  NAND2_X1 U410 ( .A1(n356), .A2(n355), .ZN(n353) );
  NOR2_X2 U411 ( .A1(n352), .A2(n350), .ZN(n354) );
  XNOR2_X1 U412 ( .A(n461), .B(KEYINPUT87), .ZN(n460) );
  NAND2_X1 U413 ( .A1(n351), .A2(n358), .ZN(n350) );
  NAND2_X1 U414 ( .A1(n466), .A2(n359), .ZN(n351) );
  XNOR2_X1 U415 ( .A(n618), .B(n617), .ZN(n819) );
  NAND2_X1 U416 ( .A1(n490), .A2(n488), .ZN(n618) );
  XNOR2_X1 U417 ( .A(n440), .B(n441), .ZN(n816) );
  NOR2_X2 U418 ( .A1(n634), .A2(n643), .ZN(n632) );
  NAND2_X1 U419 ( .A1(n383), .A2(n381), .ZN(n775) );
  AND2_X1 U420 ( .A1(n739), .A2(n730), .ZN(n702) );
  NAND2_X1 U421 ( .A1(n743), .A2(n382), .ZN(n381) );
  AND2_X1 U422 ( .A1(n394), .A2(n420), .ZN(n393) );
  AND2_X1 U423 ( .A1(n386), .A2(n384), .ZN(n383) );
  NAND2_X1 U424 ( .A1(n396), .A2(n395), .ZN(n394) );
  NAND2_X1 U425 ( .A1(n503), .A2(n408), .ZN(n479) );
  INV_X1 U426 ( .A(n693), .ZN(n743) );
  INV_X1 U427 ( .A(n410), .ZN(n396) );
  NAND2_X1 U428 ( .A1(n385), .A2(n389), .ZN(n384) );
  INV_X1 U429 ( .A(n387), .ZN(n385) );
  XNOR2_X1 U430 ( .A(n686), .B(KEYINPUT6), .ZN(n667) );
  NOR2_X1 U431 ( .A1(n415), .A2(n419), .ZN(n379) );
  NOR2_X1 U432 ( .A1(n720), .A2(G902), .ZN(n551) );
  INV_X1 U433 ( .A(n742), .ZN(n388) );
  XNOR2_X1 U434 ( .A(n404), .B(n581), .ZN(n512) );
  XNOR2_X1 U435 ( .A(n444), .B(n360), .ZN(n476) );
  XNOR2_X1 U436 ( .A(n511), .B(n510), .ZN(n509) );
  XOR2_X1 U437 ( .A(G146), .B(G125), .Z(n404) );
  XNOR2_X1 U438 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n511) );
  XNOR2_X1 U439 ( .A(KEYINPUT4), .B(KEYINPUT97), .ZN(n510) );
  INV_X4 U440 ( .A(G953), .ZN(n812) );
  NAND2_X1 U441 ( .A1(G234), .A2(G237), .ZN(n591) );
  XOR2_X1 U442 ( .A(KEYINPUT72), .B(G110), .Z(n594) );
  XOR2_X1 U443 ( .A(KEYINPUT76), .B(G113), .Z(n546) );
  INV_X1 U444 ( .A(G122), .ZN(n449) );
  XNOR2_X2 U445 ( .A(KEYINPUT100), .B(KEYINPUT101), .ZN(n535) );
  INV_X1 U446 ( .A(KEYINPUT16), .ZN(n481) );
  INV_X1 U447 ( .A(KEYINPUT34), .ZN(n532) );
  AND2_X2 U448 ( .A1(n357), .A2(n359), .ZN(n352) );
  NAND2_X1 U449 ( .A1(n349), .A2(n809), .ZN(n357) );
  NAND2_X2 U450 ( .A1(n354), .A2(n353), .ZN(n709) );
  INV_X1 U451 ( .A(n357), .ZN(n355) );
  NOR2_X1 U452 ( .A1(n466), .A2(KEYINPUT64), .ZN(n356) );
  XNOR2_X2 U453 ( .A(G140), .B(KEYINPUT68), .ZN(n444) );
  INV_X2 U454 ( .A(KEYINPUT69), .ZN(n362) );
  XNOR2_X2 U455 ( .A(n361), .B(G146), .ZN(n604) );
  XNOR2_X2 U456 ( .A(G125), .B(KEYINPUT10), .ZN(n361) );
  XNOR2_X2 U457 ( .A(n362), .B(G131), .ZN(n365) );
  XNOR2_X2 U458 ( .A(n555), .B(n363), .ZN(n806) );
  XNOR2_X2 U459 ( .A(n365), .B(n364), .ZN(n363) );
  XNOR2_X2 U460 ( .A(G137), .B(KEYINPUT4), .ZN(n364) );
  XNOR2_X2 U461 ( .A(n571), .B(G134), .ZN(n555) );
  XNOR2_X2 U462 ( .A(G143), .B(G128), .ZN(n571) );
  NAND2_X1 U463 ( .A1(n366), .A2(n514), .ZN(n513) );
  XNOR2_X1 U464 ( .A(n454), .B(n698), .ZN(n366) );
  XNOR2_X1 U465 ( .A(n427), .B(n457), .ZN(n426) );
  NAND2_X1 U466 ( .A1(n686), .A2(n742), .ZN(n676) );
  XNOR2_X2 U467 ( .A(n551), .B(n367), .ZN(n686) );
  INV_X1 U468 ( .A(n622), .ZN(n645) );
  AND2_X1 U469 ( .A1(n622), .A2(KEYINPUT34), .ZN(n524) );
  XNOR2_X2 U470 ( .A(n479), .B(n478), .ZN(n622) );
  NOR2_X1 U471 ( .A1(n639), .A2(n638), .ZN(n653) );
  XNOR2_X2 U472 ( .A(n806), .B(n486), .ZN(n599) );
  NOR2_X2 U473 ( .A1(n709), .A2(n781), .ZN(n464) );
  XNOR2_X2 U474 ( .A(n369), .B(KEYINPUT19), .ZN(n503) );
  NAND2_X2 U475 ( .A1(n656), .A2(n742), .ZN(n369) );
  XNOR2_X2 U476 ( .A(n588), .B(n587), .ZN(n656) );
  NAND2_X1 U477 ( .A1(n372), .A2(n370), .ZN(G60) );
  NAND2_X1 U478 ( .A1(n371), .A2(n377), .ZN(n370) );
  AND2_X1 U479 ( .A1(n413), .A2(n379), .ZN(n371) );
  NAND2_X1 U480 ( .A1(n374), .A2(n373), .ZN(n372) );
  NAND2_X1 U481 ( .A1(n375), .A2(KEYINPUT60), .ZN(n373) );
  NAND2_X1 U482 ( .A1(n376), .A2(n375), .ZN(n374) );
  INV_X1 U483 ( .A(n380), .ZN(n377) );
  INV_X1 U484 ( .A(n415), .ZN(n378) );
  NAND2_X1 U485 ( .A1(n693), .A2(n389), .ZN(n386) );
  NAND2_X1 U486 ( .A1(n743), .A2(n742), .ZN(n746) );
  XNOR2_X2 U487 ( .A(n604), .B(n444), .ZN(n805) );
  NAND2_X1 U488 ( .A1(n392), .A2(n390), .ZN(n399) );
  INV_X1 U489 ( .A(n438), .ZN(n391) );
  AND2_X1 U490 ( .A1(n397), .A2(n393), .ZN(n392) );
  INV_X1 U491 ( .A(G210), .ZN(n395) );
  NAND2_X1 U492 ( .A1(n438), .A2(n398), .ZN(n397) );
  AND2_X1 U493 ( .A1(n410), .A2(G210), .ZN(n398) );
  XNOR2_X1 U494 ( .A(n399), .B(n412), .ZN(G51) );
  XNOR2_X1 U495 ( .A(n632), .B(KEYINPUT91), .ZN(n603) );
  NAND2_X1 U496 ( .A1(n622), .A2(n593), .ZN(n400) );
  XNOR2_X2 U497 ( .A(n542), .B(n482), .ZN(n401) );
  XNOR2_X1 U498 ( .A(n542), .B(n482), .ZN(n574) );
  NAND2_X2 U499 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U500 ( .A(n805), .B(n611), .ZN(n473) );
  BUF_X1 U501 ( .A(n689), .Z(n446) );
  XNOR2_X1 U502 ( .A(n473), .B(n609), .ZN(n791) );
  NOR2_X1 U503 ( .A1(n791), .A2(G902), .ZN(n616) );
  NOR2_X2 U504 ( .A1(n694), .A2(n693), .ZN(n696) );
  BUF_X1 U505 ( .A(n503), .Z(n402) );
  XNOR2_X1 U506 ( .A(n403), .B(n635), .ZN(n636) );
  BUF_X1 U507 ( .A(n817), .Z(n405) );
  NOR2_X1 U508 ( .A1(n706), .A2(n794), .ZN(n779) );
  INV_X1 U509 ( .A(n577), .ZN(n576) );
  XNOR2_X1 U510 ( .A(n465), .B(n516), .ZN(n612) );
  XNOR2_X1 U511 ( .A(KEYINPUT20), .B(KEYINPUT102), .ZN(n516) );
  NAND2_X1 U512 ( .A1(n655), .A2(G234), .ZN(n465) );
  XNOR2_X1 U513 ( .A(G902), .B(KEYINPUT15), .ZN(n655) );
  OR2_X1 U514 ( .A1(G237), .A2(G902), .ZN(n584) );
  XNOR2_X1 U515 ( .A(n487), .B(n583), .ZN(n710) );
  XNOR2_X1 U516 ( .A(n512), .B(n509), .ZN(n582) );
  INV_X1 U517 ( .A(KEYINPUT78), .ZN(n707) );
  XNOR2_X1 U518 ( .A(n718), .B(n717), .ZN(n719) );
  NOR2_X1 U519 ( .A1(n747), .A2(n731), .ZN(n700) );
  INV_X1 U520 ( .A(KEYINPUT71), .ZN(n482) );
  XNOR2_X1 U521 ( .A(n568), .B(n564), .ZN(n502) );
  XNOR2_X1 U522 ( .A(G140), .B(KEYINPUT105), .ZN(n564) );
  INV_X1 U523 ( .A(KEYINPUT88), .ZN(n457) );
  NAND2_X1 U524 ( .A1(n425), .A2(n424), .ZN(n427) );
  XNOR2_X1 U525 ( .A(n586), .B(n585), .ZN(n587) );
  INV_X1 U526 ( .A(KEYINPUT28), .ZN(n484) );
  XNOR2_X1 U527 ( .A(n616), .B(n615), .ZN(n619) );
  XNOR2_X1 U528 ( .A(n515), .B(n613), .ZN(n614) );
  INV_X1 U529 ( .A(KEYINPUT0), .ZN(n478) );
  XOR2_X1 U530 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n554) );
  XNOR2_X1 U531 ( .A(KEYINPUT108), .B(KEYINPUT109), .ZN(n553) );
  XNOR2_X1 U532 ( .A(n442), .B(n432), .ZN(n431) );
  XNOR2_X1 U533 ( .A(n433), .B(KEYINPUT107), .ZN(n432) );
  XNOR2_X1 U534 ( .A(n672), .B(n499), .ZN(n498) );
  INV_X1 U535 ( .A(KEYINPUT117), .ZN(n499) );
  INV_X1 U536 ( .A(KEYINPUT118), .ZN(n496) );
  XNOR2_X1 U537 ( .A(n560), .B(n493), .ZN(n640) );
  XNOR2_X1 U538 ( .A(n494), .B(G478), .ZN(n493) );
  INV_X1 U539 ( .A(KEYINPUT110), .ZN(n494) );
  NAND2_X1 U540 ( .A1(n416), .A2(n420), .ZN(n415) );
  XNOR2_X1 U541 ( .A(n596), .B(n595), .ZN(n597) );
  XNOR2_X1 U542 ( .A(n476), .B(n594), .ZN(n598) );
  BUF_X1 U543 ( .A(n571), .Z(n577) );
  NAND2_X1 U544 ( .A1(n470), .A2(n471), .ZN(n469) );
  NAND2_X1 U545 ( .A1(n445), .A2(KEYINPUT86), .ZN(n467) );
  INV_X1 U546 ( .A(KEYINPUT48), .ZN(n472) );
  INV_X1 U547 ( .A(KEYINPUT33), .ZN(n531) );
  NAND2_X1 U548 ( .A1(n612), .A2(G217), .ZN(n515) );
  XOR2_X1 U549 ( .A(KEYINPUT81), .B(KEYINPUT80), .Z(n613) );
  XNOR2_X1 U550 ( .A(KEYINPUT5), .B(KEYINPUT75), .ZN(n545) );
  XNOR2_X1 U551 ( .A(n654), .B(KEYINPUT92), .ZN(n508) );
  XNOR2_X1 U552 ( .A(G128), .B(G110), .ZN(n605) );
  XNOR2_X1 U553 ( .A(n534), .B(n533), .ZN(n608) );
  XNOR2_X1 U554 ( .A(n535), .B(KEYINPUT84), .ZN(n534) );
  XNOR2_X1 U555 ( .A(n501), .B(n500), .ZN(n716) );
  XNOR2_X1 U556 ( .A(n475), .B(n567), .ZN(n500) );
  XNOR2_X1 U557 ( .A(n565), .B(n502), .ZN(n501) );
  INV_X1 U558 ( .A(n667), .ZN(n643) );
  XNOR2_X1 U559 ( .A(n688), .B(n483), .ZN(n690) );
  XNOR2_X1 U560 ( .A(n484), .B(KEYINPUT119), .ZN(n483) );
  NOR2_X1 U561 ( .A1(n781), .A2(n367), .ZN(n462) );
  XNOR2_X1 U562 ( .A(n430), .B(n429), .ZN(n788) );
  XNOR2_X1 U563 ( .A(n559), .B(n431), .ZN(n430) );
  NOR2_X1 U564 ( .A1(n781), .A2(n780), .ZN(n461) );
  XNOR2_X1 U565 ( .A(n497), .B(n495), .ZN(n671) );
  XNOR2_X1 U566 ( .A(n496), .B(KEYINPUT43), .ZN(n495) );
  NAND2_X1 U567 ( .A1(n498), .A2(n670), .ZN(n497) );
  XNOR2_X1 U568 ( .A(n456), .B(n455), .ZN(n820) );
  INV_X1 U569 ( .A(KEYINPUT40), .ZN(n455) );
  XNOR2_X1 U570 ( .A(n697), .B(KEYINPUT115), .ZN(n733) );
  INV_X1 U571 ( .A(KEYINPUT113), .ZN(n617) );
  NOR2_X1 U572 ( .A1(n758), .A2(n489), .ZN(n488) );
  XNOR2_X1 U573 ( .A(n790), .B(n474), .ZN(n792) );
  INV_X1 U574 ( .A(KEYINPUT60), .ZN(n419) );
  XNOR2_X1 U575 ( .A(n785), .B(n784), .ZN(n786) );
  AND2_X1 U576 ( .A1(n778), .A2(n777), .ZN(n406) );
  XNOR2_X1 U577 ( .A(n569), .B(n570), .ZN(n641) );
  INV_X1 U578 ( .A(n641), .ZN(n428) );
  AND2_X1 U579 ( .A1(n530), .A2(n529), .ZN(n407) );
  AND2_X1 U580 ( .A1(n592), .A2(n658), .ZN(n408) );
  XOR2_X1 U581 ( .A(n720), .B(KEYINPUT62), .Z(n409) );
  XOR2_X1 U582 ( .A(n713), .B(n712), .Z(n410) );
  INV_X1 U583 ( .A(KEYINPUT86), .ZN(n471) );
  XNOR2_X1 U584 ( .A(KEYINPUT96), .B(n714), .ZN(n793) );
  INV_X1 U585 ( .A(n793), .ZN(n420) );
  XOR2_X1 U586 ( .A(n721), .B(KEYINPUT94), .Z(n411) );
  XOR2_X1 U587 ( .A(n715), .B(KEYINPUT89), .Z(n412) );
  NAND2_X1 U588 ( .A1(n414), .A2(n719), .ZN(n413) );
  INV_X1 U589 ( .A(n464), .ZN(n414) );
  NAND2_X1 U590 ( .A1(n719), .A2(n418), .ZN(n416) );
  NOR2_X1 U591 ( .A1(n719), .A2(n418), .ZN(n417) );
  INV_X1 U592 ( .A(G475), .ZN(n418) );
  XNOR2_X1 U593 ( .A(n421), .B(n411), .ZN(G57) );
  NAND2_X1 U594 ( .A1(n422), .A2(n420), .ZN(n421) );
  INV_X1 U595 ( .A(n741), .ZN(n424) );
  XNOR2_X1 U596 ( .A(n513), .B(n472), .ZN(n425) );
  NAND2_X1 U597 ( .A1(n426), .A2(n740), .ZN(n706) );
  XNOR2_X1 U598 ( .A(n555), .B(n556), .ZN(n429) );
  NAND2_X1 U599 ( .A1(n521), .A2(n520), .ZN(n434) );
  NAND2_X1 U600 ( .A1(n521), .A2(n520), .ZN(n528) );
  INV_X1 U601 ( .A(G107), .ZN(n450) );
  BUF_X1 U602 ( .A(n805), .Z(n435) );
  NAND2_X1 U603 ( .A1(n450), .A2(G122), .ZN(n451) );
  NAND2_X1 U604 ( .A1(n449), .A2(G107), .ZN(n452) );
  XNOR2_X1 U605 ( .A(n689), .B(KEYINPUT1), .ZN(n620) );
  NAND2_X1 U606 ( .A1(n517), .A2(n620), .ZN(n453) );
  BUF_X1 U607 ( .A(n620), .Z(n758) );
  NOR2_X2 U608 ( .A1(n709), .A2(n781), .ZN(n438) );
  BUF_X1 U609 ( .A(n791), .Z(n439) );
  AND2_X1 U610 ( .A1(n652), .A2(n508), .ZN(n507) );
  XOR2_X1 U611 ( .A(n630), .B(KEYINPUT82), .Z(n440) );
  AND2_X1 U612 ( .A1(n632), .A2(n631), .ZN(n441) );
  BUF_X1 U613 ( .A(n573), .Z(n442) );
  NAND2_X1 U614 ( .A1(n667), .A2(n531), .ZN(n529) );
  BUF_X1 U615 ( .A(n806), .Z(n443) );
  XNOR2_X1 U616 ( .A(n574), .B(n544), .ZN(n549) );
  XNOR2_X2 U617 ( .A(n573), .B(n481), .ZN(n480) );
  XNOR2_X1 U618 ( .A(G902), .B(KEYINPUT15), .ZN(n445) );
  NAND2_X1 U619 ( .A1(n523), .A2(n407), .ZN(n522) );
  NAND2_X1 U620 ( .A1(n530), .A2(n529), .ZN(n518) );
  NOR2_X1 U621 ( .A1(n816), .A2(n448), .ZN(n447) );
  NAND2_X2 U622 ( .A1(n451), .A2(n452), .ZN(n573) );
  BUF_X1 U623 ( .A(n604), .Z(n475) );
  INV_X1 U624 ( .A(n754), .ZN(n489) );
  XNOR2_X1 U625 ( .A(n642), .B(KEYINPUT114), .ZN(n644) );
  XNOR2_X2 U626 ( .A(n453), .B(KEYINPUT74), .ZN(n642) );
  XNOR2_X2 U627 ( .A(n477), .B(KEYINPUT67), .ZN(n517) );
  NOR2_X2 U628 ( .A1(n820), .A2(n821), .ZN(n454) );
  NAND2_X1 U629 ( .A1(n704), .A2(n697), .ZN(n456) );
  XNOR2_X1 U630 ( .A(n459), .B(n458), .ZN(G75) );
  INV_X1 U631 ( .A(KEYINPUT53), .ZN(n458) );
  INV_X1 U632 ( .A(n709), .ZN(n463) );
  NAND2_X1 U633 ( .A1(n437), .A2(G478), .ZN(n787) );
  NAND2_X1 U634 ( .A1(n437), .A2(G469), .ZN(n785) );
  NAND2_X1 U635 ( .A1(n438), .A2(G217), .ZN(n790) );
  NAND2_X1 U636 ( .A1(n468), .A2(n467), .ZN(n466) );
  NAND2_X1 U637 ( .A1(n794), .A2(KEYINPUT86), .ZN(n468) );
  INV_X1 U638 ( .A(n445), .ZN(n470) );
  XNOR2_X2 U639 ( .A(n506), .B(n505), .ZN(n794) );
  XNOR2_X2 U640 ( .A(n599), .B(n600), .ZN(n783) );
  XNOR2_X2 U641 ( .A(n575), .B(n401), .ZN(n799) );
  XNOR2_X1 U642 ( .A(n439), .B(KEYINPUT126), .ZN(n474) );
  NOR2_X2 U643 ( .A1(n783), .A2(G902), .ZN(n602) );
  NAND2_X1 U644 ( .A1(n619), .A2(n753), .ZN(n477) );
  XNOR2_X2 U645 ( .A(n480), .B(n572), .ZN(n575) );
  INV_X1 U646 ( .A(n699), .ZN(n504) );
  NAND2_X1 U647 ( .A1(n485), .A2(n522), .ZN(n646) );
  NAND2_X1 U648 ( .A1(n579), .A2(n580), .ZN(n487) );
  INV_X1 U649 ( .A(n603), .ZN(n490) );
  NAND2_X1 U650 ( .A1(n507), .A2(n653), .ZN(n506) );
  NAND2_X1 U651 ( .A1(n526), .A2(n532), .ZN(n525) );
  XNOR2_X2 U652 ( .A(n492), .B(KEYINPUT35), .ZN(n817) );
  NAND2_X1 U653 ( .A1(n646), .A2(n647), .ZN(n492) );
  NAND2_X1 U654 ( .A1(n504), .A2(n402), .ZN(n731) );
  AND2_X1 U655 ( .A1(n701), .A2(n702), .ZN(n514) );
  NAND2_X1 U656 ( .A1(n517), .A2(n446), .ZN(n677) );
  NOR2_X1 U657 ( .A1(n758), .A2(n517), .ZN(n759) );
  NAND2_X1 U658 ( .A1(n518), .A2(n532), .ZN(n527) );
  NAND2_X1 U659 ( .A1(n528), .A2(n622), .ZN(n526) );
  INV_X1 U660 ( .A(n645), .ZN(n519) );
  INV_X1 U661 ( .A(n644), .ZN(n521) );
  NAND2_X1 U662 ( .A1(n407), .A2(n434), .ZN(n774) );
  NAND2_X1 U663 ( .A1(n644), .A2(n531), .ZN(n530) );
  INV_X1 U664 ( .A(KEYINPUT73), .ZN(n648) );
  XNOR2_X1 U665 ( .A(n549), .B(n548), .ZN(n550) );
  INV_X1 U666 ( .A(n716), .ZN(n718) );
  INV_X1 U667 ( .A(KEYINPUT39), .ZN(n695) );
  INV_X1 U668 ( .A(KEYINPUT63), .ZN(n721) );
  XNOR2_X1 U669 ( .A(n783), .B(n782), .ZN(n784) );
  XNOR2_X1 U670 ( .A(n696), .B(n695), .ZN(n704) );
  XNOR2_X2 U671 ( .A(G101), .B(KEYINPUT3), .ZN(n536) );
  INV_X1 U672 ( .A(n536), .ZN(n537) );
  NAND2_X1 U673 ( .A1(n537), .A2(n436), .ZN(n541) );
  INV_X1 U674 ( .A(n538), .ZN(n539) );
  NAND2_X1 U675 ( .A1(n539), .A2(n536), .ZN(n540) );
  NOR2_X1 U676 ( .A1(G953), .A2(G237), .ZN(n543) );
  XOR2_X1 U677 ( .A(KEYINPUT77), .B(n543), .Z(n566) );
  NAND2_X1 U678 ( .A1(n566), .A2(G210), .ZN(n544) );
  XNOR2_X1 U679 ( .A(n546), .B(n545), .ZN(n547) );
  XOR2_X1 U680 ( .A(KEYINPUT103), .B(n547), .Z(n548) );
  XNOR2_X1 U681 ( .A(n599), .B(n550), .ZN(n720) );
  NAND2_X1 U682 ( .A1(n612), .A2(G221), .ZN(n552) );
  XNOR2_X1 U683 ( .A(n554), .B(n553), .ZN(n556) );
  NAND2_X1 U684 ( .A1(n812), .A2(G234), .ZN(n558) );
  XNOR2_X1 U685 ( .A(n558), .B(n557), .ZN(n610) );
  NAND2_X1 U686 ( .A1(G217), .A2(n610), .ZN(n559) );
  NOR2_X1 U687 ( .A1(G902), .A2(n788), .ZN(n560) );
  XNOR2_X1 U688 ( .A(KEYINPUT13), .B(G475), .ZN(n570) );
  XOR2_X1 U689 ( .A(KEYINPUT12), .B(KEYINPUT106), .Z(n562) );
  XNOR2_X1 U690 ( .A(G131), .B(KEYINPUT11), .ZN(n561) );
  XNOR2_X1 U691 ( .A(n562), .B(n561), .ZN(n568) );
  XOR2_X2 U692 ( .A(G113), .B(G104), .Z(n572) );
  XNOR2_X1 U693 ( .A(G143), .B(n572), .ZN(n563) );
  XNOR2_X1 U694 ( .A(n563), .B(n368), .ZN(n565) );
  NAND2_X1 U695 ( .A1(G214), .A2(n566), .ZN(n567) );
  NOR2_X1 U696 ( .A1(G902), .A2(n716), .ZN(n569) );
  NOR2_X1 U697 ( .A1(n640), .A2(n641), .ZN(n691) );
  AND2_X1 U698 ( .A1(n753), .A2(n691), .ZN(n593) );
  NAND2_X1 U699 ( .A1(n799), .A2(n576), .ZN(n580) );
  INV_X1 U700 ( .A(n799), .ZN(n578) );
  NAND2_X1 U701 ( .A1(n578), .A2(n577), .ZN(n579) );
  NAND2_X1 U702 ( .A1(G224), .A2(n812), .ZN(n581) );
  XOR2_X1 U703 ( .A(n582), .B(n594), .Z(n583) );
  NAND2_X1 U704 ( .A1(n710), .A2(n445), .ZN(n588) );
  NAND2_X1 U705 ( .A1(G210), .A2(n584), .ZN(n586) );
  INV_X1 U706 ( .A(KEYINPUT98), .ZN(n585) );
  NOR2_X1 U707 ( .A1(G898), .A2(n812), .ZN(n589) );
  XOR2_X1 U708 ( .A(KEYINPUT99), .B(n589), .Z(n802) );
  NAND2_X1 U709 ( .A1(n802), .A2(G902), .ZN(n590) );
  NAND2_X1 U710 ( .A1(G952), .A2(n812), .ZN(n657) );
  NAND2_X1 U711 ( .A1(n590), .A2(n657), .ZN(n592) );
  XOR2_X1 U712 ( .A(KEYINPUT14), .B(n591), .Z(n771) );
  INV_X1 U713 ( .A(n771), .ZN(n658) );
  NAND2_X1 U714 ( .A1(G227), .A2(n812), .ZN(n596) );
  INV_X1 U715 ( .A(n595), .ZN(n818) );
  XNOR2_X2 U716 ( .A(n598), .B(n597), .ZN(n600) );
  INV_X1 U717 ( .A(G469), .ZN(n601) );
  XNOR2_X2 U718 ( .A(n602), .B(n601), .ZN(n689) );
  XOR2_X1 U719 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n606) );
  XNOR2_X1 U720 ( .A(n606), .B(n605), .ZN(n607) );
  XNOR2_X1 U721 ( .A(n608), .B(n607), .ZN(n609) );
  NAND2_X1 U722 ( .A1(n610), .A2(G221), .ZN(n611) );
  XNOR2_X1 U723 ( .A(KEYINPUT25), .B(n614), .ZN(n615) );
  BUF_X1 U724 ( .A(n619), .Z(n754) );
  NAND2_X1 U725 ( .A1(n428), .A2(n640), .ZN(n735) );
  XNOR2_X1 U726 ( .A(KEYINPUT111), .B(n735), .ZN(n703) );
  NOR2_X1 U727 ( .A1(n703), .A2(n697), .ZN(n747) );
  INV_X1 U728 ( .A(n747), .ZN(n627) );
  XOR2_X1 U729 ( .A(KEYINPUT104), .B(KEYINPUT31), .Z(n624) );
  BUF_X1 U730 ( .A(n642), .Z(n621) );
  INV_X1 U731 ( .A(n686), .ZN(n757) );
  NOR2_X1 U732 ( .A1(n621), .A2(n757), .ZN(n763) );
  NAND2_X1 U733 ( .A1(n519), .A2(n763), .ZN(n623) );
  XNOR2_X1 U734 ( .A(n624), .B(n623), .ZN(n736) );
  NOR2_X1 U735 ( .A1(n645), .A2(n677), .ZN(n625) );
  NAND2_X1 U736 ( .A1(n625), .A2(n757), .ZN(n725) );
  NAND2_X1 U737 ( .A1(n736), .A2(n725), .ZN(n626) );
  NAND2_X1 U738 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U739 ( .A(n628), .B(KEYINPUT112), .ZN(n629) );
  NAND2_X1 U740 ( .A1(n819), .A2(n629), .ZN(n639) );
  XNOR2_X1 U741 ( .A(KEYINPUT65), .B(KEYINPUT32), .ZN(n630) );
  INV_X1 U742 ( .A(n758), .ZN(n670) );
  NOR2_X1 U743 ( .A1(n754), .A2(n670), .ZN(n631) );
  NAND2_X1 U744 ( .A1(n670), .A2(n757), .ZN(n633) );
  NOR2_X1 U745 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U746 ( .A1(n816), .A2(n448), .ZN(n650) );
  NOR2_X1 U747 ( .A1(KEYINPUT73), .A2(KEYINPUT44), .ZN(n637) );
  NOR2_X1 U748 ( .A1(n650), .A2(n637), .ZN(n638) );
  NAND2_X1 U749 ( .A1(n641), .A2(n640), .ZN(n683) );
  INV_X1 U750 ( .A(n683), .ZN(n647) );
  NOR2_X2 U751 ( .A1(n817), .A2(KEYINPUT44), .ZN(n649) );
  XNOR2_X1 U752 ( .A(n649), .B(n648), .ZN(n651) );
  NAND2_X1 U753 ( .A1(n651), .A2(n447), .ZN(n652) );
  NAND2_X1 U754 ( .A1(n817), .A2(KEYINPUT44), .ZN(n654) );
  NOR2_X1 U755 ( .A1(n771), .A2(n657), .ZN(n663) );
  NAND2_X1 U756 ( .A1(G902), .A2(n658), .ZN(n659) );
  NOR2_X1 U757 ( .A1(G900), .A2(n659), .ZN(n660) );
  NAND2_X1 U758 ( .A1(G953), .A2(n660), .ZN(n661) );
  XOR2_X1 U759 ( .A(KEYINPUT116), .B(n661), .Z(n662) );
  NOR2_X1 U760 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U761 ( .A(KEYINPUT83), .B(n664), .ZN(n678) );
  AND2_X1 U762 ( .A1(n753), .A2(n678), .ZN(n665) );
  XNOR2_X1 U763 ( .A(n665), .B(KEYINPUT70), .ZN(n685) );
  NAND2_X1 U764 ( .A1(n742), .A2(n685), .ZN(n666) );
  NOR2_X1 U765 ( .A1(n733), .A2(n666), .ZN(n669) );
  NOR2_X1 U766 ( .A1(n754), .A2(n667), .ZN(n668) );
  AND2_X1 U767 ( .A1(n669), .A2(n668), .ZN(n672) );
  NOR2_X1 U768 ( .A1(n491), .A2(n671), .ZN(n741) );
  NAND2_X1 U769 ( .A1(n672), .A2(n491), .ZN(n674) );
  XNOR2_X1 U770 ( .A(KEYINPUT93), .B(KEYINPUT36), .ZN(n673) );
  XNOR2_X1 U771 ( .A(n674), .B(n673), .ZN(n675) );
  NAND2_X1 U772 ( .A1(n675), .A2(n758), .ZN(n739) );
  XOR2_X1 U773 ( .A(KEYINPUT30), .B(n676), .Z(n682) );
  INV_X1 U774 ( .A(n677), .ZN(n679) );
  NAND2_X1 U775 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U776 ( .A(n680), .B(KEYINPUT79), .ZN(n681) );
  NAND2_X1 U777 ( .A1(n682), .A2(n681), .ZN(n694) );
  NOR2_X1 U778 ( .A1(n694), .A2(n683), .ZN(n684) );
  NAND2_X1 U779 ( .A1(n684), .A2(n491), .ZN(n730) );
  NAND2_X1 U780 ( .A1(n686), .A2(n685), .ZN(n687) );
  NOR2_X1 U781 ( .A1(n687), .A2(n754), .ZN(n688) );
  NAND2_X1 U782 ( .A1(n690), .A2(n446), .ZN(n699) );
  INV_X1 U783 ( .A(n691), .ZN(n745) );
  XNOR2_X1 U784 ( .A(n692), .B(KEYINPUT42), .ZN(n821) );
  XNOR2_X1 U785 ( .A(n700), .B(KEYINPUT47), .ZN(n701) );
  NAND2_X1 U786 ( .A1(n704), .A2(n703), .ZN(n740) );
  INV_X1 U787 ( .A(n706), .ZN(n809) );
  NAND2_X1 U788 ( .A1(n470), .A2(KEYINPUT2), .ZN(n705) );
  NAND2_X1 U789 ( .A1(n779), .A2(KEYINPUT2), .ZN(n708) );
  XNOR2_X2 U790 ( .A(n708), .B(n707), .ZN(n781) );
  XOR2_X1 U791 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n713) );
  BUF_X1 U792 ( .A(n710), .Z(n711) );
  XNOR2_X1 U793 ( .A(n711), .B(KEYINPUT95), .ZN(n712) );
  NOR2_X1 U794 ( .A1(G952), .A2(n812), .ZN(n714) );
  INV_X1 U795 ( .A(KEYINPUT56), .ZN(n715) );
  XOR2_X1 U796 ( .A(KEYINPUT59), .B(KEYINPUT125), .Z(n717) );
  NOR2_X1 U797 ( .A1(n733), .A2(n725), .ZN(n722) );
  XOR2_X1 U798 ( .A(G104), .B(n722), .Z(G6) );
  XOR2_X1 U799 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n724) );
  XNOR2_X1 U800 ( .A(G107), .B(KEYINPUT120), .ZN(n723) );
  XNOR2_X1 U801 ( .A(n724), .B(n723), .ZN(n727) );
  NOR2_X1 U802 ( .A1(n735), .A2(n725), .ZN(n726) );
  XOR2_X1 U803 ( .A(n727), .B(n726), .Z(G9) );
  XOR2_X1 U804 ( .A(G110), .B(n448), .Z(G12) );
  NOR2_X1 U805 ( .A1(n735), .A2(n731), .ZN(n729) );
  XNOR2_X1 U806 ( .A(G128), .B(KEYINPUT29), .ZN(n728) );
  XNOR2_X1 U807 ( .A(n729), .B(n728), .ZN(G30) );
  XNOR2_X1 U808 ( .A(G143), .B(n730), .ZN(G45) );
  NOR2_X1 U809 ( .A1(n733), .A2(n731), .ZN(n732) );
  XOR2_X1 U810 ( .A(G146), .B(n732), .Z(G48) );
  NOR2_X1 U811 ( .A1(n736), .A2(n733), .ZN(n734) );
  XOR2_X1 U812 ( .A(G113), .B(n734), .Z(G15) );
  NOR2_X1 U813 ( .A1(n736), .A2(n735), .ZN(n737) );
  XOR2_X1 U814 ( .A(n433), .B(n737), .Z(G18) );
  XOR2_X1 U815 ( .A(G125), .B(KEYINPUT37), .Z(n738) );
  XNOR2_X1 U816 ( .A(n739), .B(n738), .ZN(G27) );
  XNOR2_X1 U817 ( .A(G134), .B(n740), .ZN(G36) );
  XOR2_X1 U818 ( .A(G140), .B(n741), .Z(G42) );
  NOR2_X1 U819 ( .A1(n743), .A2(n742), .ZN(n744) );
  NOR2_X1 U820 ( .A1(n745), .A2(n744), .ZN(n750) );
  NOR2_X1 U821 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U822 ( .A(n748), .B(KEYINPUT122), .ZN(n749) );
  NOR2_X1 U823 ( .A1(n750), .A2(n749), .ZN(n751) );
  XOR2_X1 U824 ( .A(KEYINPUT123), .B(n751), .Z(n752) );
  NOR2_X1 U825 ( .A1(n774), .A2(n752), .ZN(n768) );
  NOR2_X1 U826 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U827 ( .A(n755), .B(KEYINPUT49), .ZN(n756) );
  NAND2_X1 U828 ( .A1(n757), .A2(n756), .ZN(n761) );
  XNOR2_X1 U829 ( .A(n759), .B(KEYINPUT50), .ZN(n760) );
  NOR2_X1 U830 ( .A1(n761), .A2(n760), .ZN(n762) );
  NOR2_X1 U831 ( .A1(n763), .A2(n762), .ZN(n764) );
  XOR2_X1 U832 ( .A(KEYINPUT51), .B(n764), .Z(n765) );
  NOR2_X1 U833 ( .A1(n775), .A2(n765), .ZN(n766) );
  XOR2_X1 U834 ( .A(KEYINPUT121), .B(n766), .Z(n767) );
  NOR2_X1 U835 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U836 ( .A(n769), .B(KEYINPUT52), .ZN(n770) );
  NOR2_X1 U837 ( .A1(n771), .A2(n770), .ZN(n772) );
  NAND2_X1 U838 ( .A1(n772), .A2(G952), .ZN(n773) );
  XNOR2_X1 U839 ( .A(n773), .B(KEYINPUT124), .ZN(n778) );
  NOR2_X1 U840 ( .A1(n775), .A2(n774), .ZN(n776) );
  NOR2_X1 U841 ( .A1(G953), .A2(n776), .ZN(n777) );
  NOR2_X1 U842 ( .A1(KEYINPUT2), .A2(n779), .ZN(n780) );
  XOR2_X1 U843 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n782) );
  NOR2_X1 U844 ( .A1(n793), .A2(n786), .ZN(G54) );
  NOR2_X1 U845 ( .A1(n793), .A2(n792), .ZN(G66) );
  OR2_X1 U846 ( .A1(n794), .A2(G953), .ZN(n798) );
  NAND2_X1 U847 ( .A1(G953), .A2(G224), .ZN(n795) );
  XNOR2_X1 U848 ( .A(KEYINPUT61), .B(n795), .ZN(n796) );
  NAND2_X1 U849 ( .A1(n796), .A2(G898), .ZN(n797) );
  NAND2_X1 U850 ( .A1(n798), .A2(n797), .ZN(n804) );
  BUF_X1 U851 ( .A(n799), .Z(n800) );
  XNOR2_X1 U852 ( .A(n800), .B(G110), .ZN(n801) );
  NOR2_X1 U853 ( .A1(n802), .A2(n801), .ZN(n803) );
  XNOR2_X1 U854 ( .A(n804), .B(n803), .ZN(G69) );
  XOR2_X1 U855 ( .A(n435), .B(n443), .Z(n810) );
  XNOR2_X1 U856 ( .A(G227), .B(n810), .ZN(n807) );
  NAND2_X1 U857 ( .A1(n807), .A2(G900), .ZN(n808) );
  NAND2_X1 U858 ( .A1(n808), .A2(G953), .ZN(n815) );
  XNOR2_X1 U859 ( .A(n810), .B(n809), .ZN(n811) );
  XNOR2_X1 U860 ( .A(n811), .B(KEYINPUT127), .ZN(n813) );
  NAND2_X1 U861 ( .A1(n813), .A2(n812), .ZN(n814) );
  NAND2_X1 U862 ( .A1(n815), .A2(n814), .ZN(G72) );
  XOR2_X1 U863 ( .A(G119), .B(n816), .Z(G21) );
  XOR2_X1 U864 ( .A(n405), .B(n368), .Z(G24) );
  XNOR2_X1 U865 ( .A(n819), .B(n818), .ZN(G3) );
  XOR2_X1 U866 ( .A(n820), .B(G131), .Z(G33) );
  XOR2_X1 U867 ( .A(G137), .B(n821), .Z(G39) );
endmodule

