//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 1 0 1 1 0 1 0 0 1 1 0 1 0 1 0 0 0 0 1 1 0 1 0 1 0 1 1 1 0 0 0 1 1 1 0 0 1 0 0 1 0 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:31 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1254, new_n1255,
    new_n1256, new_n1257, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  AOI21_X1  g0005(.A(G50), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G77), .ZN(new_n207));
  AND2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(G353));
  OAI21_X1  g0008(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(KEYINPUT66), .ZN(new_n211));
  INV_X1    g0011(.A(KEYINPUT66), .ZN(new_n212));
  NAND3_X1  g0012(.A1(new_n212), .A2(G1), .A3(G13), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(G20), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n204), .A2(new_n205), .ZN(new_n218));
  INV_X1    g0018(.A(G50), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  XOR2_X1   g0021(.A(KEYINPUT67), .B(G238), .Z(new_n222));
  OR2_X1    g0022(.A1(new_n222), .A2(new_n203), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G107), .A2(G264), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n227));
  AND4_X1   g0027(.A1(new_n224), .A2(new_n225), .A3(new_n226), .A4(new_n227), .ZN(new_n228));
  AOI22_X1  g0028(.A1(new_n223), .A2(new_n228), .B1(G1), .B2(G20), .ZN(new_n229));
  INV_X1    g0029(.A(KEYINPUT1), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n221), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  INV_X1    g0031(.A(G1), .ZN(new_n232));
  NOR3_X1   g0032(.A1(new_n232), .A2(new_n216), .A3(G13), .ZN(new_n233));
  OAI211_X1 g0033(.A(new_n233), .B(G250), .C1(G257), .C2(G264), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n234), .B(KEYINPUT65), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT0), .ZN(new_n236));
  AOI211_X1 g0036(.A(new_n231), .B(new_n236), .C1(new_n230), .C2(new_n229), .ZN(G361));
  XOR2_X1   g0037(.A(G238), .B(G244), .Z(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT68), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(KEYINPUT2), .B(G226), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G264), .B(G270), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G358));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n219), .A2(G68), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n203), .A2(G50), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(G58), .B(G77), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n249), .B(new_n254), .ZN(G351));
  XNOR2_X1  g0055(.A(KEYINPUT15), .B(G87), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n216), .A2(G33), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  AOI22_X1  g0059(.A1(new_n257), .A2(new_n259), .B1(G20), .B2(G77), .ZN(new_n260));
  NOR2_X1   g0060(.A1(G20), .A2(G33), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n262), .A2(KEYINPUT71), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n202), .A2(KEYINPUT8), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT8), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G58), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT71), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n267), .B1(new_n268), .B2(new_n261), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n260), .B1(new_n263), .B2(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n211), .A2(new_n213), .A3(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n232), .A2(G13), .A3(G20), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  AOI22_X1  g0074(.A1(new_n270), .A2(new_n272), .B1(new_n207), .B2(new_n274), .ZN(new_n275));
  NAND4_X1  g0075(.A1(new_n211), .A2(new_n213), .A3(new_n273), .A4(new_n271), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n232), .A2(G20), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n277), .A2(G77), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n275), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n210), .B1(G33), .B2(G41), .ZN(new_n281));
  INV_X1    g0081(.A(G41), .ZN(new_n282));
  INV_X1    g0082(.A(G45), .ZN(new_n283));
  AOI21_X1  g0083(.A(G1), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n281), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G244), .ZN(new_n286));
  INV_X1    g0086(.A(G274), .ZN(new_n287));
  INV_X1    g0087(.A(new_n210), .ZN(new_n288));
  NAND2_X1  g0088(.A1(G33), .A2(G41), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n287), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(new_n284), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n286), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g0092(.A(KEYINPUT3), .B(G33), .ZN(new_n293));
  INV_X1    g0093(.A(G1698), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n293), .A2(G232), .A3(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G107), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n293), .A2(G1698), .ZN(new_n297));
  OAI221_X1 g0097(.A(new_n295), .B1(new_n296), .B2(new_n293), .C1(new_n297), .C2(new_n222), .ZN(new_n298));
  AND2_X1   g0098(.A1(new_n214), .A2(new_n289), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n292), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n280), .B1(G190), .B2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G200), .ZN(new_n302));
  OR2_X1    g0102(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G179), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n300), .A2(new_n305), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n280), .B(new_n306), .C1(G169), .C2(new_n300), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n285), .A2(G226), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(new_n291), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n293), .A2(G222), .A3(new_n294), .ZN(new_n310));
  INV_X1    g0110(.A(G223), .ZN(new_n311));
  OAI221_X1 g0111(.A(new_n310), .B1(new_n207), .B2(new_n293), .C1(new_n297), .C2(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n309), .B1(new_n312), .B2(new_n299), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G169), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  XNOR2_X1  g0116(.A(KEYINPUT8), .B(G58), .ZN(new_n317));
  INV_X1    g0117(.A(G150), .ZN(new_n318));
  OAI22_X1  g0118(.A1(new_n317), .A2(new_n258), .B1(new_n318), .B2(new_n262), .ZN(new_n319));
  OAI22_X1  g0119(.A1(new_n319), .A2(KEYINPUT69), .B1(new_n216), .B2(new_n206), .ZN(new_n320));
  AOI22_X1  g0120(.A1(new_n267), .A2(new_n259), .B1(G150), .B2(new_n261), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT69), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n272), .B1(new_n320), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n278), .A2(G50), .ZN(new_n325));
  OAI22_X1  g0125(.A1(new_n276), .A2(new_n325), .B1(G50), .B2(new_n273), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(KEYINPUT70), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT70), .ZN(new_n328));
  OAI221_X1 g0128(.A(new_n328), .B1(G50), .B2(new_n273), .C1(new_n276), .C2(new_n325), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n324), .A2(new_n330), .ZN(new_n331));
  OAI211_X1 g0131(.A(new_n316), .B(new_n331), .C1(G179), .C2(new_n314), .ZN(new_n332));
  AND3_X1   g0132(.A1(new_n304), .A2(new_n307), .A3(new_n332), .ZN(new_n333));
  AOI22_X1  g0133(.A1(new_n261), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n334), .B1(new_n207), .B2(new_n258), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(new_n272), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT11), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n274), .A2(new_n203), .ZN(new_n339));
  XNOR2_X1  g0139(.A(new_n339), .B(KEYINPUT12), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n335), .A2(KEYINPUT11), .A3(new_n272), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n277), .A2(G68), .A3(new_n278), .ZN(new_n342));
  AND4_X1   g0142(.A1(new_n338), .A2(new_n340), .A3(new_n341), .A4(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(G33), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(KEYINPUT3), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT3), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(G33), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n346), .A2(new_n348), .A3(G232), .A4(G1698), .ZN(new_n349));
  NAND4_X1  g0149(.A1(new_n346), .A2(new_n348), .A3(G226), .A4(new_n294), .ZN(new_n350));
  INV_X1    g0150(.A(G97), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n349), .B(new_n350), .C1(new_n345), .C2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n299), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT13), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n285), .A2(G238), .B1(new_n290), .B2(new_n284), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n354), .B1(new_n353), .B2(new_n355), .ZN(new_n358));
  OAI21_X1  g0158(.A(G169), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  XNOR2_X1  g0159(.A(new_n359), .B(KEYINPUT14), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n353), .A2(new_n355), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(KEYINPUT13), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n362), .A2(G179), .A3(new_n356), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT74), .ZN(new_n364));
  XNOR2_X1  g0164(.A(new_n363), .B(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n344), .B1(new_n360), .B2(new_n365), .ZN(new_n366));
  OAI21_X1  g0166(.A(G200), .B1(new_n357), .B2(new_n358), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n362), .A2(G190), .A3(new_n356), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n367), .A2(new_n368), .A3(new_n343), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT73), .ZN(new_n370));
  XNOR2_X1  g0170(.A(new_n369), .B(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n333), .A2(new_n366), .A3(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT72), .ZN(new_n373));
  AND3_X1   g0173(.A1(new_n324), .A2(new_n330), .A3(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n373), .B1(new_n324), .B2(new_n330), .ZN(new_n375));
  OAI21_X1  g0175(.A(KEYINPUT9), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n331), .A2(KEYINPUT72), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT9), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n324), .A2(new_n330), .A3(new_n373), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n377), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n376), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT10), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n313), .A2(new_n302), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n383), .B1(G190), .B2(new_n313), .ZN(new_n384));
  AND3_X1   g0184(.A1(new_n381), .A2(new_n382), .A3(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n382), .B1(new_n381), .B2(new_n384), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n372), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT79), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n267), .A2(new_n278), .ZN(new_n390));
  OAI22_X1  g0190(.A1(new_n390), .A2(new_n276), .B1(new_n267), .B2(new_n273), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(G226), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n297), .A2(new_n393), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n346), .A2(new_n348), .A3(G223), .A4(new_n294), .ZN(new_n395));
  INV_X1    g0195(.A(G87), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n395), .B1(new_n345), .B2(new_n396), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n299), .B1(new_n394), .B2(new_n397), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n285), .A2(G232), .B1(new_n290), .B2(new_n284), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(new_n302), .ZN(new_n401));
  AND2_X1   g0201(.A1(KEYINPUT77), .A2(G190), .ZN(new_n402));
  NOR2_X1   g0202(.A1(KEYINPUT77), .A2(G190), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n401), .B1(new_n400), .B2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n272), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT7), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n408), .B1(new_n293), .B2(G20), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n347), .A2(G33), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n345), .A2(KEYINPUT3), .ZN(new_n411));
  OAI211_X1 g0211(.A(KEYINPUT7), .B(new_n216), .C1(new_n410), .C2(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n203), .B1(new_n409), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(G58), .A2(G68), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n204), .A2(new_n205), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(G20), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n261), .A2(G159), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n413), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n407), .B1(new_n419), .B2(KEYINPUT16), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT16), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n421), .B1(new_n413), .B2(new_n418), .ZN(new_n422));
  AOI21_X1  g0222(.A(KEYINPUT75), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n346), .A2(new_n348), .ZN(new_n424));
  AOI21_X1  g0224(.A(KEYINPUT7), .B1(new_n424), .B2(new_n216), .ZN(new_n425));
  AOI211_X1 g0225(.A(new_n408), .B(G20), .C1(new_n346), .C2(new_n348), .ZN(new_n426));
  OAI21_X1  g0226(.A(G68), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  AOI22_X1  g0227(.A1(new_n415), .A2(G20), .B1(G159), .B2(new_n261), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n427), .A2(KEYINPUT16), .A3(new_n428), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n429), .A2(new_n422), .A3(KEYINPUT75), .A4(new_n272), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n392), .B(new_n406), .C1(new_n423), .C2(new_n431), .ZN(new_n432));
  AND2_X1   g0232(.A1(KEYINPUT78), .A2(KEYINPUT17), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NOR2_X1   g0234(.A1(KEYINPUT78), .A2(KEYINPUT17), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n429), .A2(new_n422), .A3(new_n272), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT75), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n391), .B1(new_n439), .B2(new_n430), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n436), .B1(new_n440), .B2(new_n406), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n434), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT18), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n392), .B1(new_n423), .B2(new_n431), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n400), .A2(G169), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n445), .B1(new_n305), .B2(new_n400), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n443), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n446), .ZN(new_n448));
  NOR3_X1   g0248(.A1(new_n440), .A2(KEYINPUT18), .A3(new_n448), .ZN(new_n449));
  OAI21_X1  g0249(.A(KEYINPUT76), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n444), .A2(new_n443), .A3(new_n446), .ZN(new_n451));
  OAI21_X1  g0251(.A(KEYINPUT18), .B1(new_n440), .B2(new_n448), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT76), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n442), .B1(new_n450), .B2(new_n454), .ZN(new_n455));
  AND3_X1   g0255(.A1(new_n388), .A2(new_n389), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n389), .B1(new_n388), .B2(new_n455), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n232), .A2(G33), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n277), .A2(G116), .A3(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(G116), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n274), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g0263(.A(G20), .B1(G33), .B2(G283), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n345), .A2(G97), .ZN(new_n465));
  AOI22_X1  g0265(.A1(new_n464), .A2(new_n465), .B1(G20), .B2(new_n462), .ZN(new_n466));
  AND3_X1   g0266(.A1(new_n466), .A2(new_n272), .A3(KEYINPUT20), .ZN(new_n467));
  AOI21_X1  g0267(.A(KEYINPUT20), .B1(new_n466), .B2(new_n272), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n461), .B(new_n463), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n346), .A2(new_n348), .A3(G264), .A4(G1698), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n346), .A2(new_n348), .A3(G257), .A4(new_n294), .ZN(new_n471));
  INV_X1    g0271(.A(G303), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n470), .B(new_n471), .C1(new_n472), .C2(new_n293), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(new_n299), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT82), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT5), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n475), .B1(new_n476), .B2(G41), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n282), .A2(KEYINPUT82), .A3(KEYINPUT5), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n283), .A2(G1), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n476), .A2(G41), .ZN(new_n480));
  AND4_X1   g0280(.A1(new_n477), .A2(new_n478), .A3(new_n479), .A4(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(new_n290), .ZN(new_n482));
  INV_X1    g0282(.A(new_n281), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n479), .A2(new_n480), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n476), .A2(G41), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n483), .B(G270), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n474), .A2(new_n482), .A3(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n469), .A2(new_n487), .A3(G169), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT21), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n487), .A2(G200), .ZN(new_n491));
  INV_X1    g0291(.A(new_n469), .ZN(new_n492));
  AND2_X1   g0292(.A1(new_n482), .A2(new_n486), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n493), .A2(new_n405), .A3(new_n474), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n491), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n469), .A2(G179), .A3(new_n474), .A4(new_n493), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n469), .A2(new_n487), .A3(KEYINPUT21), .A4(G169), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n490), .A2(new_n495), .A3(new_n496), .A4(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT88), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AND2_X1   g0300(.A1(new_n497), .A2(new_n496), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n501), .A2(KEYINPUT88), .A3(new_n490), .A4(new_n495), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n261), .A2(G77), .ZN(new_n504));
  XNOR2_X1  g0304(.A(new_n504), .B(KEYINPUT80), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT6), .ZN(new_n506));
  NOR3_X1   g0306(.A1(new_n506), .A2(new_n351), .A3(G107), .ZN(new_n507));
  XNOR2_X1  g0307(.A(G97), .B(G107), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n507), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n505), .B1(new_n216), .B2(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n296), .B1(new_n409), .B2(new_n412), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n272), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n273), .A2(G97), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT81), .ZN(new_n514));
  XNOR2_X1  g0314(.A(new_n513), .B(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n276), .B1(new_n232), .B2(G33), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n515), .B1(G97), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n512), .A2(new_n517), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n346), .A2(new_n348), .A3(G244), .A4(new_n294), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT4), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n293), .A2(KEYINPUT4), .A3(G244), .A4(new_n294), .ZN(new_n522));
  NAND2_X1  g0322(.A1(G33), .A2(G283), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n293), .A2(G250), .A3(G1698), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n521), .A2(new_n522), .A3(new_n523), .A4(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n299), .ZN(new_n526));
  INV_X1    g0326(.A(new_n484), .ZN(new_n527));
  INV_X1    g0327(.A(new_n485), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n281), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n529), .A2(G257), .B1(new_n290), .B2(new_n481), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n526), .A2(new_n530), .A3(new_n305), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n518), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n526), .A2(new_n530), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT83), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n526), .A2(new_n530), .A3(KEYINPUT83), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n532), .B1(new_n537), .B2(new_n315), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT84), .ZN(new_n539));
  AND3_X1   g0339(.A1(new_n526), .A2(new_n530), .A3(KEYINPUT83), .ZN(new_n540));
  AOI21_X1  g0340(.A(KEYINPUT83), .B1(new_n526), .B2(new_n530), .ZN(new_n541));
  INV_X1    g0341(.A(G190), .ZN(new_n542));
  NOR3_X1   g0342(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n533), .A2(G200), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n544), .A2(new_n512), .A3(new_n517), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n539), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n535), .A2(G190), .A3(new_n536), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n302), .B1(new_n526), .B2(new_n530), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n518), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n547), .A2(new_n549), .A3(KEYINPUT84), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n538), .B1(new_n546), .B2(new_n550), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n346), .A2(new_n348), .A3(G257), .A4(G1698), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n346), .A2(new_n348), .A3(G250), .A4(new_n294), .ZN(new_n553));
  NAND2_X1  g0353(.A1(G33), .A2(G294), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n299), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n483), .B(G264), .C1(new_n484), .C2(new_n485), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n556), .A2(new_n482), .A3(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n558), .A2(KEYINPUT90), .A3(G169), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n556), .A2(G179), .A3(new_n482), .A4(new_n557), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(KEYINPUT90), .B1(new_n558), .B2(G169), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT24), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n346), .A2(new_n348), .A3(new_n216), .A4(G87), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(KEYINPUT22), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT22), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n293), .A2(new_n566), .A3(new_n216), .A4(G87), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT89), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n569), .B1(new_n216), .B2(G107), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(KEYINPUT23), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT23), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n569), .B(new_n572), .C1(new_n216), .C2(G107), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n571), .A2(new_n573), .B1(G116), .B2(new_n259), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n563), .B1(new_n568), .B2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n568), .A2(new_n563), .A3(new_n574), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n407), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n516), .A2(G107), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n274), .A2(new_n296), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT25), .ZN(new_n581));
  XNOR2_X1  g0381(.A(new_n580), .B(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  OAI22_X1  g0383(.A1(new_n561), .A2(new_n562), .B1(new_n578), .B2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n577), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n272), .B1(new_n585), .B2(new_n575), .ZN(new_n586));
  OR2_X1    g0386(.A1(new_n558), .A2(new_n542), .ZN(new_n587));
  INV_X1    g0387(.A(new_n583), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n558), .A2(G200), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n586), .A2(new_n587), .A3(new_n588), .A4(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n584), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n346), .A2(new_n348), .A3(G244), .A4(G1698), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n346), .A2(new_n348), .A3(G238), .A4(new_n294), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n592), .B(new_n593), .C1(new_n345), .C2(new_n462), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n299), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n479), .A2(new_n287), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n483), .B(new_n596), .C1(G250), .C2(new_n479), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n595), .A2(new_n305), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(KEYINPUT85), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n595), .A2(new_n597), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n315), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT85), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n595), .A2(new_n602), .A3(new_n305), .A4(new_n597), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n293), .A2(new_n216), .A3(G68), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT19), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n605), .B1(new_n258), .B2(new_n351), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n608));
  AND2_X1   g0408(.A1(new_n608), .A2(new_n216), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n396), .A2(new_n351), .A3(new_n296), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT86), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n396), .A2(new_n351), .A3(new_n296), .A4(KEYINPUT86), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n609), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n272), .B1(new_n607), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n516), .A2(new_n257), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n257), .A2(new_n273), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n615), .A2(new_n616), .A3(new_n618), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n599), .A2(new_n601), .A3(new_n603), .A4(new_n619), .ZN(new_n620));
  AND2_X1   g0420(.A1(new_n615), .A2(new_n618), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n600), .A2(G200), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n516), .A2(G87), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n595), .A2(G190), .A3(new_n597), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n621), .A2(new_n622), .A3(new_n623), .A4(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT87), .ZN(new_n626));
  AND3_X1   g0426(.A1(new_n620), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n626), .B1(new_n620), .B2(new_n625), .ZN(new_n628));
  NOR3_X1   g0428(.A1(new_n591), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  AND4_X1   g0429(.A1(new_n459), .A2(new_n503), .A3(new_n551), .A4(new_n629), .ZN(G372));
  NAND3_X1  g0430(.A1(new_n601), .A2(new_n619), .A3(new_n598), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n590), .A2(new_n625), .A3(new_n631), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n501), .A2(new_n490), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n633), .B1(new_n634), .B2(new_n584), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n632), .B1(new_n635), .B2(new_n551), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n625), .A2(new_n631), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n538), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT26), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n620), .A2(new_n625), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(KEYINPUT87), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n620), .A2(new_n625), .A3(new_n626), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n643), .A2(new_n538), .A3(KEYINPUT26), .A4(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n636), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n459), .A2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT91), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n649), .B1(new_n385), .B2(new_n386), .ZN(new_n650));
  NOR3_X1   g0450(.A1(new_n374), .A2(new_n375), .A3(KEYINPUT9), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n378), .B1(new_n377), .B2(new_n379), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n384), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(KEYINPUT10), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n381), .A2(new_n382), .A3(new_n384), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n654), .A2(KEYINPUT91), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n650), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g0457(.A(new_n369), .B(KEYINPUT73), .ZN(new_n658));
  OR2_X1    g0458(.A1(new_n658), .A2(new_n307), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n442), .B1(new_n659), .B2(new_n366), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n451), .A2(new_n452), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n657), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n662), .A2(new_n332), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n648), .A2(new_n663), .ZN(G369));
  NAND3_X1  g0464(.A1(new_n500), .A2(KEYINPUT93), .A3(new_n502), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n232), .A2(new_n216), .A3(G13), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n666), .A2(KEYINPUT27), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(KEYINPUT27), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n667), .A2(new_n668), .A3(G213), .ZN(new_n669));
  XOR2_X1   g0469(.A(KEYINPUT92), .B(G343), .Z(new_n670));
  NOR2_X1   g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n492), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT93), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n673), .B1(new_n503), .B2(new_n674), .ZN(new_n675));
  AOI22_X1  g0475(.A1(new_n665), .A2(new_n675), .B1(new_n634), .B2(new_n673), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(G330), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n584), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(new_n671), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n671), .B1(new_n578), .B2(new_n583), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n584), .A2(new_n590), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n678), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n501), .A2(new_n490), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(new_n672), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n686), .A2(new_n591), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n687), .B1(new_n679), .B2(new_n672), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n684), .A2(new_n688), .ZN(G399));
  AND2_X1   g0489(.A1(new_n612), .A2(new_n613), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(new_n462), .ZN(new_n691));
  INV_X1    g0491(.A(new_n233), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(G41), .ZN(new_n693));
  NOR3_X1   g0493(.A1(new_n691), .A2(new_n232), .A3(new_n693), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n694), .B1(new_n220), .B2(new_n693), .ZN(new_n695));
  XOR2_X1   g0495(.A(new_n695), .B(KEYINPUT28), .Z(new_n696));
  NAND2_X1  g0496(.A1(new_n647), .A2(new_n672), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT29), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(KEYINPUT94), .A3(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT94), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n671), .B1(new_n636), .B2(new_n646), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n700), .B1(new_n701), .B2(KEYINPUT29), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n640), .B1(new_n538), .B2(new_n638), .ZN(new_n703));
  INV_X1    g0503(.A(new_n538), .ZN(new_n704));
  NOR3_X1   g0504(.A1(new_n704), .A2(new_n627), .A3(new_n628), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n703), .B1(new_n705), .B2(new_n640), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n671), .B1(new_n706), .B2(new_n636), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(KEYINPUT29), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n699), .A2(new_n702), .A3(new_n708), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n629), .A2(new_n551), .A3(new_n503), .A4(new_n672), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n474), .A2(G179), .A3(new_n482), .A4(new_n486), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n556), .A2(new_n557), .ZN(new_n712));
  NOR3_X1   g0512(.A1(new_n711), .A2(new_n600), .A3(new_n712), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n713), .A2(new_n535), .A3(new_n536), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT30), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n713), .A2(new_n535), .A3(KEYINPUT30), .A4(new_n536), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n533), .A2(new_n558), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n487), .A2(new_n305), .A3(new_n600), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n716), .A2(new_n717), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(new_n671), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT31), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n720), .B1(new_n714), .B2(new_n715), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n672), .B1(new_n726), .B2(new_n717), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(KEYINPUT31), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n710), .A2(new_n725), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(G330), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n709), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT95), .ZN(new_n732));
  XNOR2_X1  g0532(.A(new_n731), .B(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n696), .B1(new_n733), .B2(G1), .ZN(G364));
  AND2_X1   g0534(.A1(new_n216), .A2(G13), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n232), .B1(new_n735), .B2(G45), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n693), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n678), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n676), .A2(G330), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(G13), .A2(G33), .ZN(new_n742));
  XNOR2_X1  g0542(.A(new_n742), .B(KEYINPUT98), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(G20), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  OR2_X1    g0545(.A1(new_n676), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n738), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n216), .A2(new_n305), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(G200), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(G190), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR3_X1   g0551(.A1(new_n542), .A2(G179), .A3(G200), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(new_n216), .ZN(new_n753));
  OAI22_X1  g0553(.A1(new_n751), .A2(new_n203), .B1(new_n753), .B2(new_n351), .ZN(new_n754));
  OR2_X1    g0554(.A1(new_n754), .A2(KEYINPUT100), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(KEYINPUT100), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n216), .A2(G179), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n757), .A2(new_n542), .A3(G200), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n296), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n749), .A2(new_n404), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n759), .B1(G50), .B2(new_n760), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n757), .A2(G190), .A3(G200), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(new_n396), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G190), .A2(G200), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n757), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(G159), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n763), .B1(new_n768), .B2(KEYINPUT32), .ZN(new_n769));
  NAND4_X1  g0569(.A1(new_n755), .A2(new_n756), .A3(new_n761), .A4(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(KEYINPUT32), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n424), .B1(new_n767), .B2(new_n771), .ZN(new_n772));
  XOR2_X1   g0572(.A(new_n748), .B(KEYINPUT99), .Z(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(new_n764), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n404), .A2(G200), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  OAI221_X1 g0576(.A(new_n772), .B1(new_n774), .B2(new_n207), .C1(new_n202), .C2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n765), .ZN(new_n778));
  AND2_X1   g0578(.A1(new_n778), .A2(G329), .ZN(new_n779));
  AOI211_X1 g0579(.A(new_n293), .B(new_n779), .C1(G326), .C2(new_n760), .ZN(new_n780));
  INV_X1    g0580(.A(new_n776), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G322), .ZN(new_n782));
  INV_X1    g0582(.A(G311), .ZN(new_n783));
  OAI211_X1 g0583(.A(new_n780), .B(new_n782), .C1(new_n783), .C2(new_n774), .ZN(new_n784));
  INV_X1    g0584(.A(new_n753), .ZN(new_n785));
  INV_X1    g0585(.A(new_n762), .ZN(new_n786));
  AOI22_X1  g0586(.A1(new_n785), .A2(G294), .B1(new_n786), .B2(G303), .ZN(new_n787));
  INV_X1    g0587(.A(G283), .ZN(new_n788));
  XOR2_X1   g0588(.A(KEYINPUT33), .B(G317), .Z(new_n789));
  OAI221_X1 g0589(.A(new_n787), .B1(new_n788), .B2(new_n758), .C1(new_n751), .C2(new_n789), .ZN(new_n790));
  OAI22_X1  g0590(.A1(new_n770), .A2(new_n777), .B1(new_n784), .B2(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n215), .B1(G20), .B2(new_n315), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n747), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n792), .A2(new_n744), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n293), .A2(new_n233), .ZN(new_n796));
  XOR2_X1   g0596(.A(new_n796), .B(KEYINPUT96), .Z(new_n797));
  AOI22_X1  g0597(.A1(new_n797), .A2(G355), .B1(new_n462), .B2(new_n692), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n220), .A2(new_n283), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n692), .A2(new_n293), .ZN(new_n800));
  OAI211_X1 g0600(.A(new_n799), .B(new_n800), .C1(new_n254), .C2(new_n283), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n795), .B1(new_n802), .B2(KEYINPUT97), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n803), .B1(KEYINPUT97), .B2(new_n802), .ZN(new_n804));
  AND2_X1   g0604(.A1(new_n793), .A2(new_n804), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n739), .A2(new_n741), .B1(new_n746), .B2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(G396));
  NAND2_X1  g0607(.A1(new_n280), .A2(new_n671), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n304), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(new_n307), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n307), .A2(new_n671), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n697), .A2(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n811), .B1(new_n809), .B2(new_n307), .ZN(new_n815));
  INV_X1    g0615(.A(new_n550), .ZN(new_n816));
  AOI21_X1  g0616(.A(KEYINPUT84), .B1(new_n547), .B2(new_n549), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n704), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  OAI211_X1 g0618(.A(new_n590), .B(new_n638), .C1(new_n679), .C2(new_n685), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n631), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  AND2_X1   g0620(.A1(new_n641), .A2(new_n645), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n672), .B(new_n815), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n814), .A2(new_n822), .ZN(new_n823));
  OR2_X1    g0623(.A1(new_n823), .A2(new_n730), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n738), .B1(new_n823), .B2(new_n730), .ZN(new_n825));
  AND2_X1   g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n743), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n792), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n747), .B1(new_n828), .B2(new_n207), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n753), .A2(new_n351), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n424), .B1(new_n765), .B2(new_n783), .ZN(new_n831));
  INV_X1    g0631(.A(new_n774), .ZN(new_n832));
  AOI211_X1 g0632(.A(new_n830), .B(new_n831), .C1(new_n832), .C2(G116), .ZN(new_n833));
  INV_X1    g0633(.A(G294), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n833), .B1(new_n834), .B2(new_n776), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n396), .A2(new_n758), .B1(new_n762), .B2(new_n296), .ZN(new_n836));
  INV_X1    g0636(.A(new_n760), .ZN(new_n837));
  OAI22_X1  g0637(.A1(new_n788), .A2(new_n751), .B1(new_n837), .B2(new_n472), .ZN(new_n838));
  NOR3_X1   g0638(.A1(new_n835), .A2(new_n836), .A3(new_n838), .ZN(new_n839));
  AOI22_X1  g0639(.A1(G137), .A2(new_n760), .B1(new_n750), .B2(G150), .ZN(new_n840));
  INV_X1    g0640(.A(G143), .ZN(new_n841));
  OAI221_X1 g0641(.A(new_n840), .B1(new_n776), .B2(new_n841), .C1(new_n766), .C2(new_n774), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n842), .B(KEYINPUT34), .ZN(new_n843));
  INV_X1    g0643(.A(G132), .ZN(new_n844));
  OAI221_X1 g0644(.A(new_n293), .B1(new_n765), .B2(new_n844), .C1(new_n753), .C2(new_n202), .ZN(new_n845));
  OAI22_X1  g0645(.A1(new_n219), .A2(new_n762), .B1(new_n758), .B2(new_n203), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n839), .B1(new_n843), .B2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n792), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n829), .B1(new_n848), .B2(new_n849), .C1(new_n743), .C2(new_n815), .ZN(new_n850));
  XOR2_X1   g0650(.A(new_n850), .B(KEYINPUT101), .Z(new_n851));
  NOR2_X1   g0651(.A1(new_n826), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(G384));
  INV_X1    g0653(.A(new_n509), .ZN(new_n854));
  OR2_X1    g0654(.A1(new_n854), .A2(KEYINPUT35), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(KEYINPUT35), .ZN(new_n856));
  NAND4_X1  g0656(.A1(new_n855), .A2(G116), .A3(new_n217), .A4(new_n856), .ZN(new_n857));
  XOR2_X1   g0657(.A(new_n857), .B(KEYINPUT36), .Z(new_n858));
  NAND3_X1  g0658(.A1(new_n220), .A2(G77), .A3(new_n414), .ZN(new_n859));
  AOI211_X1 g0659(.A(new_n232), .B(G13), .C1(new_n859), .C2(new_n250), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT105), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n661), .A2(new_n669), .ZN(new_n863));
  XOR2_X1   g0663(.A(new_n811), .B(KEYINPUT102), .Z(new_n864));
  NAND2_X1  g0664(.A1(new_n822), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n343), .A2(new_n672), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT14), .ZN(new_n867));
  XNOR2_X1  g0667(.A(new_n359), .B(new_n867), .ZN(new_n868));
  XNOR2_X1  g0668(.A(new_n363), .B(KEYINPUT74), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n343), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n866), .B1(new_n870), .B2(new_n658), .ZN(new_n871));
  INV_X1    g0671(.A(new_n866), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n366), .A2(new_n371), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n865), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n444), .A2(new_n446), .ZN(new_n876));
  INV_X1    g0676(.A(new_n669), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n444), .A2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT37), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n876), .A2(new_n878), .A3(new_n879), .A4(new_n432), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n429), .A2(new_n272), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n427), .A2(new_n428), .ZN(new_n882));
  OR2_X1    g0682(.A1(new_n882), .A2(KEYINPUT103), .ZN(new_n883));
  AOI21_X1  g0683(.A(KEYINPUT16), .B1(new_n882), .B2(KEYINPUT103), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n881), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  OAI22_X1  g0685(.A1(new_n885), .A2(new_n391), .B1(new_n446), .B2(new_n877), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n432), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(KEYINPUT37), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n880), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n885), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n669), .B1(new_n890), .B2(new_n392), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n889), .B1(new_n455), .B2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT38), .ZN(new_n894));
  OR2_X1    g0694(.A1(new_n434), .A2(new_n441), .ZN(new_n895));
  AND3_X1   g0695(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n453), .B1(new_n451), .B2(new_n452), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n895), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n891), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n894), .B1(new_n880), .B2(new_n888), .ZN(new_n900));
  AOI22_X1  g0700(.A1(new_n893), .A2(new_n894), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n863), .B1(new_n875), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n900), .B1(new_n455), .B2(new_n892), .ZN(new_n903));
  INV_X1    g0703(.A(new_n889), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n904), .B1(new_n898), .B2(new_n891), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n903), .B1(new_n905), .B2(KEYINPUT38), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(KEYINPUT39), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n440), .A2(new_n669), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n908), .B1(new_n442), .B2(new_n661), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n432), .B1(new_n440), .B2(new_n448), .ZN(new_n910));
  OAI21_X1  g0710(.A(KEYINPUT37), .B1(new_n910), .B2(new_n908), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n880), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n909), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n894), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT39), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n914), .A2(new_n903), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(KEYINPUT104), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT104), .ZN(new_n918));
  NAND4_X1  g0718(.A1(new_n914), .A2(new_n903), .A3(new_n918), .A4(new_n915), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n907), .A2(new_n917), .A3(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n366), .A2(new_n671), .ZN(new_n921));
  AOI211_X1 g0721(.A(new_n862), .B(new_n902), .C1(new_n920), .C2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n919), .B1(new_n901), .B2(new_n915), .ZN(new_n923));
  AOI21_X1  g0723(.A(KEYINPUT38), .B1(new_n909), .B2(new_n912), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n924), .B1(new_n899), .B2(new_n900), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n918), .B1(new_n925), .B2(new_n915), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n921), .B1(new_n923), .B2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(new_n902), .ZN(new_n928));
  AOI21_X1  g0728(.A(KEYINPUT105), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n922), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n663), .B1(new_n709), .B2(new_n458), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n930), .B(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT106), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n723), .A2(new_n933), .A3(new_n724), .ZN(new_n934));
  OAI21_X1  g0734(.A(KEYINPUT106), .B1(new_n727), .B2(KEYINPUT31), .ZN(new_n935));
  NAND4_X1  g0735(.A1(new_n710), .A2(new_n934), .A3(new_n935), .A4(new_n728), .ZN(new_n936));
  AND2_X1   g0736(.A1(new_n459), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n813), .B1(new_n871), .B2(new_n873), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n939), .B1(new_n903), .B2(new_n914), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT40), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n936), .A2(new_n938), .A3(new_n941), .ZN(new_n942));
  OAI22_X1  g0742(.A1(new_n940), .A2(new_n941), .B1(new_n901), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(G330), .B1(new_n937), .B2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n945), .A2(KEYINPUT107), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n937), .A2(new_n943), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n945), .A2(KEYINPUT107), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n946), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n932), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n232), .B2(new_n735), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n932), .A2(new_n949), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n861), .B1(new_n951), .B2(new_n952), .ZN(G367));
  XNOR2_X1  g0753(.A(new_n731), .B(KEYINPUT95), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n518), .A2(new_n671), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n551), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n538), .A2(new_n671), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n688), .A2(new_n958), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n959), .B(KEYINPUT45), .Z(new_n960));
  NOR2_X1   g0760(.A1(new_n688), .A2(new_n958), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT44), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(new_n684), .ZN(new_n964));
  INV_X1    g0764(.A(new_n683), .ZN(new_n965));
  AOI21_X1  g0765(.A(KEYINPUT109), .B1(new_n965), .B2(new_n686), .ZN(new_n966));
  MUX2_X1   g0766(.A(new_n966), .B(KEYINPUT109), .S(new_n687), .Z(new_n967));
  XNOR2_X1  g0767(.A(new_n967), .B(new_n677), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n954), .B1(new_n964), .B2(new_n968), .ZN(new_n969));
  XNOR2_X1  g0769(.A(KEYINPUT108), .B(KEYINPUT41), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n693), .B(new_n970), .Z(new_n971));
  OAI21_X1  g0771(.A(new_n736), .B1(new_n969), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n958), .A2(new_n687), .ZN(new_n973));
  OR2_X1    g0773(.A1(new_n973), .A2(KEYINPUT42), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n679), .B1(new_n816), .B2(new_n817), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n671), .B1(new_n975), .B2(new_n704), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n976), .B1(new_n973), .B2(KEYINPUT42), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n621), .A2(new_n623), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(new_n671), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n638), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n980), .B1(new_n631), .B2(new_n979), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n974), .A2(new_n977), .B1(KEYINPUT43), .B2(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n981), .A2(KEYINPUT43), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n982), .B(new_n983), .Z(new_n984));
  INV_X1    g0784(.A(new_n958), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n684), .A2(new_n985), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n984), .B(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n972), .A2(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n794), .B1(new_n233), .B2(new_n256), .ZN(new_n989));
  AND2_X1   g0789(.A1(new_n245), .A2(new_n800), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n738), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  AOI22_X1  g0791(.A1(G143), .A2(new_n760), .B1(new_n750), .B2(G159), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n785), .A2(G68), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n992), .B(new_n993), .C1(new_n207), .C2(new_n758), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n424), .B1(new_n778), .B2(G137), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n995), .B1(new_n202), .B2(new_n762), .C1(new_n774), .C2(new_n219), .ZN(new_n996));
  AOI211_X1 g0796(.A(new_n994), .B(new_n996), .C1(G150), .C2(new_n781), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n293), .B1(new_n778), .B2(G317), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n998), .B1(new_n296), .B2(new_n753), .C1(new_n776), .C2(new_n472), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT46), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(new_n762), .B2(new_n462), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n786), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1002));
  OAI211_X1 g0802(.A(new_n1001), .B(new_n1002), .C1(new_n774), .C2(new_n788), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n758), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n760), .A2(G311), .B1(new_n1004), .B2(G97), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n834), .B2(new_n751), .ZN(new_n1006));
  NOR3_X1   g0806(.A1(new_n999), .A2(new_n1003), .A3(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n997), .A2(new_n1007), .ZN(new_n1008));
  XOR2_X1   g0808(.A(new_n1008), .B(KEYINPUT47), .Z(new_n1009));
  AOI21_X1  g0809(.A(new_n991), .B1(new_n1009), .B2(new_n792), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1010), .B1(new_n745), .B2(new_n981), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n988), .A2(new_n1011), .ZN(G387));
  NOR2_X1   g0812(.A1(new_n733), .A2(new_n968), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n733), .A2(new_n968), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(new_n693), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1013), .B1(new_n1015), .B2(KEYINPUT112), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(KEYINPUT112), .B2(new_n1015), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n965), .A2(new_n744), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n797), .A2(new_n691), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1019), .B1(G107), .B2(new_n233), .ZN(new_n1020));
  AOI211_X1 g0820(.A(G45), .B(new_n691), .C1(G68), .C2(G77), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT110), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n317), .A2(G50), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT50), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1023), .A2(new_n1024), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n800), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(new_n242), .B2(G45), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1020), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n738), .B1(new_n1030), .B2(new_n795), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n753), .A2(new_n256), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n837), .A2(new_n766), .B1(new_n207), .B2(new_n762), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n1032), .B(new_n1033), .C1(new_n267), .C2(new_n750), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n293), .B1(new_n765), .B2(new_n318), .C1(new_n351), .C2(new_n758), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1035), .B1(new_n781), .B2(G50), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1034), .B(new_n1036), .C1(new_n203), .C2(new_n774), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n293), .B1(new_n778), .B2(G326), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n753), .A2(new_n788), .B1(new_n762), .B2(new_n834), .ZN(new_n1039));
  XOR2_X1   g0839(.A(new_n1039), .B(KEYINPUT111), .Z(new_n1040));
  AOI22_X1  g0840(.A1(G322), .A2(new_n760), .B1(new_n750), .B2(G311), .ZN(new_n1041));
  INV_X1    g0841(.A(G317), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n1041), .B1(new_n776), .B2(new_n1042), .C1(new_n472), .C2(new_n774), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT48), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1040), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1045), .B1(new_n1044), .B2(new_n1043), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT49), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n1038), .B1(new_n462), .B2(new_n758), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1048));
  AND2_X1   g0848(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1037), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1031), .B1(new_n1050), .B2(new_n792), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n968), .A2(new_n737), .B1(new_n1018), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1017), .A2(new_n1052), .ZN(G393));
  OAI22_X1  g0853(.A1(new_n776), .A2(new_n783), .B1(new_n1042), .B2(new_n837), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n1054), .B(KEYINPUT52), .Z(new_n1055));
  OAI22_X1  g0855(.A1(new_n751), .A2(new_n472), .B1(new_n788), .B2(new_n762), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(G116), .B2(new_n785), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n293), .B(new_n759), .C1(G322), .C2(new_n778), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1057), .B(new_n1058), .C1(new_n834), .C2(new_n774), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n776), .A2(new_n766), .B1(new_n318), .B2(new_n837), .ZN(new_n1060));
  XOR2_X1   g0860(.A(new_n1060), .B(KEYINPUT51), .Z(new_n1061));
  OAI221_X1 g0861(.A(new_n293), .B1(new_n765), .B2(new_n841), .C1(new_n396), .C2(new_n758), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(new_n832), .B2(new_n267), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(G77), .A2(new_n785), .B1(new_n750), .B2(G50), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n1063), .B(new_n1064), .C1(new_n203), .C2(new_n762), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n1055), .A2(new_n1059), .B1(new_n1061), .B2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(new_n792), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n249), .A2(new_n1028), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n794), .B1(new_n351), .B2(new_n233), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1067), .B(new_n738), .C1(new_n1068), .C2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(new_n985), .B2(new_n744), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(new_n964), .B2(new_n737), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1014), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1073), .A2(new_n964), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n693), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n1073), .A2(new_n964), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1072), .B1(new_n1075), .B2(new_n1076), .ZN(G390));
  INV_X1    g0877(.A(new_n921), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n864), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1079), .B1(new_n701), .B2(new_n815), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n874), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1078), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n907), .A2(new_n917), .A3(new_n919), .A4(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n889), .A2(KEYINPUT38), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(new_n898), .B2(new_n891), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n811), .B1(new_n707), .B2(new_n810), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n1078), .B1(new_n1085), .B2(new_n924), .C1(new_n1086), .C2(new_n1081), .ZN(new_n1087));
  INV_X1    g0887(.A(G330), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n813), .A2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n729), .A2(new_n874), .A3(new_n1089), .ZN(new_n1090));
  AND3_X1   g0890(.A1(new_n1083), .A2(new_n1087), .A3(new_n1090), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n936), .A2(new_n874), .A3(new_n1089), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(new_n1083), .B2(new_n1087), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  NOR3_X1   g0894(.A1(new_n1085), .A2(KEYINPUT39), .A3(new_n924), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n1095), .A2(new_n918), .B1(new_n906), .B2(KEYINPUT39), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1096), .A2(new_n827), .A3(new_n917), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n747), .B1(new_n828), .B2(new_n317), .ZN(new_n1098));
  XOR2_X1   g0898(.A(new_n1098), .B(KEYINPUT114), .Z(new_n1099));
  AND2_X1   g0899(.A1(new_n778), .A2(G125), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n424), .B(new_n1100), .C1(G128), .C2(new_n760), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n753), .A2(new_n766), .B1(new_n758), .B2(new_n219), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(G137), .B2(new_n750), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1101), .B(new_n1103), .C1(new_n844), .C2(new_n776), .ZN(new_n1104));
  OR3_X1    g0904(.A1(new_n762), .A2(KEYINPUT53), .A3(new_n318), .ZN(new_n1105));
  OAI21_X1  g0905(.A(KEYINPUT53), .B1(new_n762), .B2(new_n318), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(KEYINPUT54), .B(G143), .ZN(new_n1107));
  XOR2_X1   g0907(.A(new_n1107), .B(KEYINPUT115), .Z(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n1105), .B(new_n1106), .C1(new_n1109), .C2(new_n774), .ZN(new_n1110));
  AOI211_X1 g0910(.A(new_n293), .B(new_n763), .C1(G294), .C2(new_n778), .ZN(new_n1111));
  OAI221_X1 g0911(.A(new_n1111), .B1(new_n351), .B2(new_n774), .C1(new_n462), .C2(new_n776), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n785), .A2(G77), .B1(new_n1004), .B2(G68), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n1113), .B1(new_n296), .B2(new_n751), .C1(new_n788), .C2(new_n837), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n1104), .A2(new_n1110), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1099), .B1(new_n1115), .B2(new_n792), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n1094), .A2(new_n737), .B1(new_n1097), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT113), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n693), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1083), .A2(new_n1087), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1092), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1083), .A2(new_n1087), .A3(new_n1090), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n729), .A2(new_n1089), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(new_n1081), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1080), .B1(new_n1126), .B2(new_n1092), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n936), .A2(new_n1089), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(new_n1081), .ZN(new_n1129));
  AND2_X1   g0929(.A1(new_n1086), .A2(new_n1090), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1127), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  OAI211_X1 g0931(.A(G330), .B(new_n936), .C1(new_n456), .C2(new_n457), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n1132), .B(new_n663), .C1(new_n709), .C2(new_n458), .ZN(new_n1133));
  OR2_X1    g0933(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1119), .B1(new_n1124), .B2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1122), .A2(new_n1123), .A3(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1118), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1134), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1139));
  AND4_X1   g0939(.A1(new_n1118), .A2(new_n1139), .A3(new_n1137), .A4(new_n693), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1117), .B1(new_n1138), .B2(new_n1140), .ZN(G378));
  AOI21_X1  g0941(.A(new_n1078), .B1(new_n1096), .B2(new_n917), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n862), .B1(new_n1142), .B2(new_n902), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n936), .B(new_n938), .C1(new_n1085), .C2(new_n924), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n942), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n1144), .A2(KEYINPUT40), .B1(new_n906), .B2(new_n1145), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n669), .B1(new_n377), .B2(new_n379), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1150), .B1(new_n657), .B2(new_n332), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n332), .ZN(new_n1152));
  AOI211_X1 g0952(.A(new_n1152), .B(new_n1149), .C1(new_n650), .C2(new_n656), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1148), .B1(new_n1151), .B2(new_n1153), .ZN(new_n1154));
  NOR3_X1   g0954(.A1(new_n385), .A2(new_n386), .A3(new_n649), .ZN(new_n1155));
  AOI21_X1  g0955(.A(KEYINPUT91), .B1(new_n654), .B2(new_n655), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n332), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(new_n1149), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n657), .A2(new_n332), .A3(new_n1150), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1158), .A2(new_n1159), .A3(new_n1147), .ZN(new_n1160));
  AND2_X1   g0960(.A1(new_n1154), .A2(new_n1160), .ZN(new_n1161));
  NOR3_X1   g0961(.A1(new_n1146), .A2(new_n1161), .A3(new_n1088), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1154), .A2(new_n1160), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(new_n943), .B2(G330), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n927), .A2(KEYINPUT105), .A3(new_n928), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1143), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1161), .B1(new_n1146), .B2(new_n1088), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n943), .A2(G330), .A3(new_n1163), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1170), .B1(new_n922), .B2(new_n929), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1167), .A2(new_n1171), .A3(new_n737), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n747), .B1(new_n828), .B2(new_n219), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n424), .A2(new_n282), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(G283), .B2(new_n778), .ZN(new_n1175));
  OAI221_X1 g0975(.A(new_n1175), .B1(new_n202), .B2(new_n758), .C1(new_n207), .C2(new_n762), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n1176), .B(KEYINPUT116), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n993), .B1(new_n751), .B2(new_n351), .C1(new_n462), .C2(new_n837), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n296), .A2(new_n776), .B1(new_n774), .B2(new_n256), .ZN(new_n1179));
  NOR3_X1   g0979(.A1(new_n1177), .A2(new_n1178), .A3(new_n1179), .ZN(new_n1180));
  XOR2_X1   g0980(.A(new_n1180), .B(KEYINPUT58), .Z(new_n1181));
  OAI211_X1 g0981(.A(new_n1174), .B(new_n219), .C1(G33), .C2(G41), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n760), .A2(G125), .ZN(new_n1183));
  OAI221_X1 g0983(.A(new_n1183), .B1(new_n318), .B2(new_n753), .C1(new_n751), .C2(new_n844), .ZN(new_n1184));
  INV_X1    g0984(.A(G128), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n1109), .A2(new_n762), .B1(new_n776), .B2(new_n1185), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n1184), .B(new_n1186), .C1(G137), .C2(new_n832), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1188), .A2(KEYINPUT59), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1188), .A2(KEYINPUT59), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1004), .A2(G159), .ZN(new_n1191));
  AOI211_X1 g0991(.A(G33), .B(G41), .C1(new_n778), .C2(G124), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1190), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1181), .B(new_n1182), .C1(new_n1189), .C2(new_n1193), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1194), .A2(KEYINPUT117), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(KEYINPUT117), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1196), .A2(new_n792), .ZN(new_n1197));
  OAI221_X1 g0997(.A(new_n1173), .B1(new_n1195), .B2(new_n1197), .C1(new_n1163), .C2(new_n743), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1172), .A2(new_n1198), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(new_n1133), .B(KEYINPUT118), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1137), .A2(new_n1200), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1201), .A2(KEYINPUT57), .A3(new_n1167), .A4(new_n1171), .ZN(new_n1202));
  AND2_X1   g1002(.A1(new_n1202), .A2(new_n693), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT57), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1167), .A2(new_n1171), .ZN(new_n1205));
  INV_X1    g1005(.A(KEYINPUT118), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1133), .B(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(new_n1094), .B2(new_n1136), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1204), .B1(new_n1205), .B2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1199), .B1(new_n1203), .B2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1210), .A2(KEYINPUT119), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1209), .A2(new_n693), .A3(new_n1202), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1199), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT119), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1211), .A2(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(G375));
  OR2_X1    g1018(.A1(new_n1131), .A2(new_n736), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n293), .B1(new_n1004), .B2(G77), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1220), .B1(new_n776), .B2(new_n788), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1032), .B1(G116), .B2(new_n750), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1222), .B1(new_n834), .B2(new_n837), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n762), .A2(new_n351), .B1(new_n765), .B2(new_n472), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1223), .B1(KEYINPUT120), .B2(new_n1224), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1225), .B1(KEYINPUT120), .B2(new_n1224), .ZN(new_n1226));
  AOI211_X1 g1026(.A(new_n1221), .B(new_n1226), .C1(G107), .C2(new_n832), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1228), .A2(KEYINPUT121), .ZN(new_n1229));
  OAI221_X1 g1029(.A(new_n293), .B1(new_n765), .B2(new_n1185), .C1(new_n202), .C2(new_n758), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(new_n832), .B2(G150), .ZN(new_n1231));
  OAI22_X1  g1031(.A1(new_n837), .A2(new_n844), .B1(new_n219), .B2(new_n753), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(G159), .B2(new_n786), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1108), .A2(new_n750), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n781), .A2(G137), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1231), .A2(new_n1233), .A3(new_n1234), .A4(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT121), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1236), .B1(new_n1227), .B2(new_n1237), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n792), .B1(new_n1229), .B2(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n747), .B1(new_n828), .B2(new_n203), .ZN(new_n1240));
  OAI211_X1 g1040(.A(new_n1239), .B(new_n1240), .C1(new_n743), .C2(new_n874), .ZN(new_n1241));
  AND2_X1   g1041(.A1(new_n1219), .A2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n971), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1134), .A2(new_n1243), .A3(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1242), .A2(new_n1245), .ZN(new_n1246));
  XOR2_X1   g1046(.A(new_n1246), .B(KEYINPUT122), .Z(G381));
  NOR4_X1   g1047(.A1(G381), .A2(G387), .A3(G390), .A4(G384), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(new_n1117), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(G393), .A2(G396), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1217), .A2(new_n1248), .A3(new_n1251), .A4(new_n1252), .ZN(G407));
  NAND2_X1  g1053(.A1(new_n670), .A2(G213), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1217), .A2(new_n1251), .A3(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(G407), .A2(G213), .A3(new_n1256), .ZN(new_n1257));
  XNOR2_X1  g1057(.A(new_n1257), .B(KEYINPUT123), .ZN(G409));
  INV_X1    g1058(.A(KEYINPUT60), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1244), .B1(new_n1136), .B2(new_n1259), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1131), .A2(new_n1133), .A3(KEYINPUT60), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1260), .A2(new_n693), .A3(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(new_n1242), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(new_n852), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1262), .A2(G384), .A3(new_n1242), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1255), .A2(G2897), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(new_n1266), .B(new_n1267), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1201), .A2(new_n1243), .A3(new_n1167), .A4(new_n1171), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1250), .B1(new_n1213), .B2(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1270), .B1(new_n1210), .B2(G378), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1268), .B1(new_n1271), .B2(new_n1255), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT61), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1212), .A2(G378), .A3(new_n1213), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1213), .A2(new_n1269), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(new_n1251), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1274), .A2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT62), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1266), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1277), .A2(new_n1278), .A3(new_n1254), .A4(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1272), .A2(new_n1273), .A3(new_n1280), .ZN(new_n1281));
  XOR2_X1   g1081(.A(KEYINPUT125), .B(KEYINPUT62), .Z(new_n1282));
  AOI21_X1  g1082(.A(new_n1255), .B1(new_n1274), .B2(new_n1276), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1282), .B1(new_n1283), .B2(new_n1279), .ZN(new_n1284));
  OAI21_X1  g1084(.A(KEYINPUT126), .B1(new_n1281), .B2(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n806), .B1(new_n1017), .B2(new_n1052), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1252), .A2(new_n1286), .ZN(new_n1287));
  XNOR2_X1  g1087(.A(G387), .B(G390), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(G387), .ZN(new_n1290));
  AND2_X1   g1090(.A1(new_n1290), .A2(G390), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1290), .A2(G390), .ZN(new_n1292));
  OAI22_X1  g1092(.A1(new_n1291), .A2(new_n1292), .B1(new_n1252), .B2(new_n1286), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1289), .A2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1283), .A2(new_n1279), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1282), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1277), .A2(new_n1254), .ZN(new_n1298));
  AOI21_X1  g1098(.A(KEYINPUT61), .B1(new_n1298), .B2(new_n1268), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT126), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1297), .A2(new_n1299), .A3(new_n1300), .A4(new_n1280), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1285), .A2(new_n1294), .A3(new_n1301), .ZN(new_n1302));
  XNOR2_X1  g1102(.A(KEYINPUT124), .B(KEYINPUT63), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1294), .B1(new_n1295), .B2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT63), .ZN(new_n1305));
  OAI211_X1 g1105(.A(new_n1304), .B(new_n1299), .C1(new_n1305), .C2(new_n1295), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1302), .A2(new_n1306), .ZN(G405));
  AND3_X1   g1107(.A1(new_n1212), .A2(KEYINPUT119), .A3(new_n1213), .ZN(new_n1308));
  AOI21_X1  g1108(.A(KEYINPUT119), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1309));
  NOR3_X1   g1109(.A1(new_n1308), .A2(new_n1309), .A3(new_n1250), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1274), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1266), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1312));
  AND2_X1   g1112(.A1(new_n1289), .A2(new_n1293), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1211), .A2(new_n1216), .A3(new_n1251), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1314), .A2(new_n1279), .A3(new_n1274), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1312), .A2(new_n1313), .A3(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(KEYINPUT127), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT127), .ZN(new_n1318));
  NAND4_X1  g1118(.A1(new_n1312), .A2(new_n1313), .A3(new_n1315), .A4(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1312), .A2(new_n1315), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1320), .A2(new_n1294), .ZN(new_n1321));
  AND3_X1   g1121(.A1(new_n1317), .A2(new_n1319), .A3(new_n1321), .ZN(G402));
endmodule


