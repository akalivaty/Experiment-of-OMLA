

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582;

  XOR2_X1 U321 ( .A(KEYINPUT100), .B(n399), .Z(n289) );
  XOR2_X1 U322 ( .A(G127GAT), .B(KEYINPUT78), .Z(n290) );
  OR2_X1 U323 ( .A1(n521), .A2(n519), .ZN(n397) );
  INV_X1 U324 ( .A(n576), .ZN(n443) );
  NAND2_X1 U325 ( .A1(n443), .A2(n547), .ZN(n444) );
  XNOR2_X1 U326 ( .A(n380), .B(G176GAT), .ZN(n381) );
  INV_X1 U327 ( .A(n419), .ZN(n420) );
  XNOR2_X1 U328 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U329 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U330 ( .A(n391), .B(n390), .ZN(n392) );
  XOR2_X1 U331 ( .A(n551), .B(KEYINPUT73), .Z(n476) );
  XNOR2_X1 U332 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U333 ( .A(n393), .B(n392), .ZN(n395) );
  NOR2_X1 U334 ( .A1(n521), .A2(n470), .ZN(n560) );
  INV_X1 U335 ( .A(G106GAT), .ZN(n448) );
  XOR2_X1 U336 ( .A(KEYINPUT94), .B(n405), .Z(n565) );
  XOR2_X1 U337 ( .A(n395), .B(n394), .Z(n521) );
  XNOR2_X1 U338 ( .A(KEYINPUT58), .B(G190GAT), .ZN(n471) );
  XNOR2_X1 U339 ( .A(n448), .B(KEYINPUT44), .ZN(n449) );
  XNOR2_X1 U340 ( .A(n472), .B(n471), .ZN(G1351GAT) );
  XOR2_X1 U341 ( .A(KEYINPUT2), .B(KEYINPUT86), .Z(n292) );
  XNOR2_X1 U342 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n291) );
  XNOR2_X1 U343 ( .A(n292), .B(n291), .ZN(n293) );
  XOR2_X1 U344 ( .A(G141GAT), .B(n293), .Z(n360) );
  XOR2_X1 U345 ( .A(G211GAT), .B(KEYINPUT21), .Z(n295) );
  XNOR2_X1 U346 ( .A(G197GAT), .B(KEYINPUT85), .ZN(n294) );
  XNOR2_X1 U347 ( .A(n295), .B(n294), .ZN(n374) );
  XOR2_X1 U348 ( .A(G50GAT), .B(G162GAT), .Z(n419) );
  XOR2_X1 U349 ( .A(n374), .B(n419), .Z(n297) );
  XNOR2_X1 U350 ( .A(G218GAT), .B(G106GAT), .ZN(n296) );
  XNOR2_X1 U351 ( .A(n297), .B(n296), .ZN(n298) );
  XNOR2_X1 U352 ( .A(n360), .B(n298), .ZN(n311) );
  XOR2_X1 U353 ( .A(KEYINPUT88), .B(KEYINPUT84), .Z(n300) );
  XNOR2_X1 U354 ( .A(KEYINPUT87), .B(KEYINPUT23), .ZN(n299) );
  XNOR2_X1 U355 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U356 ( .A(G78GAT), .B(KEYINPUT22), .Z(n302) );
  XNOR2_X1 U357 ( .A(G22GAT), .B(G148GAT), .ZN(n301) );
  XNOR2_X1 U358 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U359 ( .A(n304), .B(n303), .Z(n309) );
  XOR2_X1 U360 ( .A(KEYINPUT24), .B(G204GAT), .Z(n306) );
  NAND2_X1 U361 ( .A1(G228GAT), .A2(G233GAT), .ZN(n305) );
  XNOR2_X1 U362 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U363 ( .A(KEYINPUT89), .B(n307), .ZN(n308) );
  XNOR2_X1 U364 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U365 ( .A(n311), .B(n310), .ZN(n466) );
  XOR2_X1 U366 ( .A(n466), .B(KEYINPUT28), .Z(n514) );
  XOR2_X1 U367 ( .A(KEYINPUT69), .B(G141GAT), .Z(n313) );
  XNOR2_X1 U368 ( .A(G113GAT), .B(G197GAT), .ZN(n312) );
  XNOR2_X1 U369 ( .A(n313), .B(n312), .ZN(n329) );
  XOR2_X1 U370 ( .A(G43GAT), .B(G50GAT), .Z(n315) );
  XNOR2_X1 U371 ( .A(G169GAT), .B(G36GAT), .ZN(n314) );
  XNOR2_X1 U372 ( .A(n315), .B(n314), .ZN(n318) );
  XOR2_X1 U373 ( .A(G1GAT), .B(G8GAT), .Z(n317) );
  XNOR2_X1 U374 ( .A(G15GAT), .B(G22GAT), .ZN(n316) );
  XNOR2_X1 U375 ( .A(n317), .B(n316), .ZN(n429) );
  XOR2_X1 U376 ( .A(n318), .B(n429), .Z(n327) );
  XOR2_X1 U377 ( .A(KEYINPUT71), .B(KEYINPUT30), .Z(n320) );
  XNOR2_X1 U378 ( .A(KEYINPUT68), .B(KEYINPUT70), .ZN(n319) );
  XNOR2_X1 U379 ( .A(n320), .B(n319), .ZN(n325) );
  XNOR2_X1 U380 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n321) );
  XNOR2_X1 U381 ( .A(n321), .B(KEYINPUT7), .ZN(n418) );
  XOR2_X1 U382 ( .A(n418), .B(KEYINPUT29), .Z(n323) );
  NAND2_X1 U383 ( .A1(G229GAT), .A2(G233GAT), .ZN(n322) );
  XNOR2_X1 U384 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U385 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U386 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U387 ( .A(n329), .B(n328), .ZN(n540) );
  XOR2_X1 U388 ( .A(G92GAT), .B(G85GAT), .Z(n331) );
  XNOR2_X1 U389 ( .A(G99GAT), .B(G106GAT), .ZN(n330) );
  XNOR2_X1 U390 ( .A(n331), .B(n330), .ZN(n411) );
  XOR2_X1 U391 ( .A(n411), .B(KEYINPUT31), .Z(n333) );
  NAND2_X1 U392 ( .A1(G230GAT), .A2(G233GAT), .ZN(n332) );
  XNOR2_X1 U393 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U394 ( .A(n334), .B(KEYINPUT32), .ZN(n336) );
  XOR2_X1 U395 ( .A(G148GAT), .B(G57GAT), .Z(n346) );
  XOR2_X1 U396 ( .A(n346), .B(KEYINPUT33), .Z(n335) );
  XNOR2_X1 U397 ( .A(n336), .B(n335), .ZN(n338) );
  XNOR2_X1 U398 ( .A(G176GAT), .B(G204GAT), .ZN(n337) );
  XNOR2_X1 U399 ( .A(n337), .B(G64GAT), .ZN(n369) );
  XNOR2_X1 U400 ( .A(n338), .B(n369), .ZN(n340) );
  XOR2_X1 U401 ( .A(G120GAT), .B(G71GAT), .Z(n386) );
  XOR2_X1 U402 ( .A(G78GAT), .B(KEYINPUT13), .Z(n428) );
  XNOR2_X1 U403 ( .A(n386), .B(n428), .ZN(n339) );
  XNOR2_X1 U404 ( .A(n340), .B(n339), .ZN(n570) );
  XNOR2_X1 U405 ( .A(n570), .B(KEYINPUT41), .ZN(n341) );
  XNOR2_X1 U406 ( .A(KEYINPUT64), .B(n341), .ZN(n544) );
  XNOR2_X1 U407 ( .A(KEYINPUT107), .B(n544), .ZN(n557) );
  NAND2_X1 U408 ( .A1(n540), .A2(n557), .ZN(n342) );
  XOR2_X1 U409 ( .A(KEYINPUT108), .B(n342), .Z(n504) );
  XNOR2_X1 U410 ( .A(KEYINPUT37), .B(KEYINPUT102), .ZN(n446) );
  XOR2_X1 U411 ( .A(G85GAT), .B(G162GAT), .Z(n344) );
  XNOR2_X1 U412 ( .A(G29GAT), .B(G134GAT), .ZN(n343) );
  XNOR2_X1 U413 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U414 ( .A(n346), .B(n345), .Z(n348) );
  NAND2_X1 U415 ( .A1(G225GAT), .A2(G233GAT), .ZN(n347) );
  XNOR2_X1 U416 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U417 ( .A(n349), .B(KEYINPUT1), .Z(n352) );
  XNOR2_X1 U418 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n350) );
  XNOR2_X1 U419 ( .A(n290), .B(n350), .ZN(n382) );
  XNOR2_X1 U420 ( .A(n382), .B(KEYINPUT5), .ZN(n351) );
  XNOR2_X1 U421 ( .A(n352), .B(n351), .ZN(n356) );
  XOR2_X1 U422 ( .A(KEYINPUT91), .B(KEYINPUT90), .Z(n354) );
  XNOR2_X1 U423 ( .A(G1GAT), .B(G120GAT), .ZN(n353) );
  XNOR2_X1 U424 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U425 ( .A(n356), .B(n355), .Z(n362) );
  XOR2_X1 U426 ( .A(KEYINPUT4), .B(KEYINPUT92), .Z(n358) );
  XNOR2_X1 U427 ( .A(KEYINPUT93), .B(KEYINPUT6), .ZN(n357) );
  XNOR2_X1 U428 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U429 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U430 ( .A(n362), .B(n361), .ZN(n405) );
  XOR2_X1 U431 ( .A(G92GAT), .B(KEYINPUT95), .Z(n364) );
  NAND2_X1 U432 ( .A1(G226GAT), .A2(G233GAT), .ZN(n363) );
  XNOR2_X1 U433 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U434 ( .A(KEYINPUT96), .B(n365), .Z(n368) );
  XNOR2_X1 U435 ( .A(G36GAT), .B(G190GAT), .ZN(n366) );
  XNOR2_X1 U436 ( .A(n366), .B(G218GAT), .ZN(n410) );
  XNOR2_X1 U437 ( .A(n410), .B(G8GAT), .ZN(n367) );
  XNOR2_X1 U438 ( .A(n368), .B(n367), .ZN(n370) );
  XOR2_X1 U439 ( .A(n370), .B(n369), .Z(n376) );
  XOR2_X1 U440 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n372) );
  XNOR2_X1 U441 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n371) );
  XNOR2_X1 U442 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U443 ( .A(G169GAT), .B(n373), .Z(n394) );
  XNOR2_X1 U444 ( .A(n394), .B(n374), .ZN(n375) );
  XOR2_X1 U445 ( .A(n376), .B(n375), .Z(n519) );
  XOR2_X1 U446 ( .A(n519), .B(KEYINPUT97), .Z(n377) );
  XNOR2_X1 U447 ( .A(n377), .B(KEYINPUT27), .ZN(n401) );
  NOR2_X1 U448 ( .A1(n565), .A2(n401), .ZN(n378) );
  XOR2_X1 U449 ( .A(KEYINPUT98), .B(n378), .Z(n537) );
  INV_X1 U450 ( .A(n514), .ZN(n379) );
  NOR2_X1 U451 ( .A1(n537), .A2(n379), .ZN(n523) );
  AND2_X1 U452 ( .A1(G227GAT), .A2(G233GAT), .ZN(n380) );
  XOR2_X1 U453 ( .A(G43GAT), .B(G134GAT), .Z(n417) );
  XNOR2_X1 U454 ( .A(n383), .B(n417), .ZN(n393) );
  XOR2_X1 U455 ( .A(KEYINPUT79), .B(KEYINPUT80), .Z(n385) );
  XNOR2_X1 U456 ( .A(G99GAT), .B(G190GAT), .ZN(n384) );
  XNOR2_X1 U457 ( .A(n385), .B(n384), .ZN(n387) );
  XOR2_X1 U458 ( .A(n387), .B(n386), .Z(n391) );
  XOR2_X1 U459 ( .A(KEYINPUT81), .B(KEYINPUT82), .Z(n389) );
  XNOR2_X1 U460 ( .A(G15GAT), .B(KEYINPUT20), .ZN(n388) );
  XNOR2_X1 U461 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U462 ( .A(KEYINPUT83), .B(n521), .Z(n396) );
  AND2_X1 U463 ( .A1(n523), .A2(n396), .ZN(n407) );
  XNOR2_X1 U464 ( .A(KEYINPUT99), .B(n397), .ZN(n398) );
  NOR2_X1 U465 ( .A1(n398), .A2(n466), .ZN(n399) );
  XNOR2_X1 U466 ( .A(KEYINPUT25), .B(n289), .ZN(n403) );
  NAND2_X1 U467 ( .A1(n521), .A2(n466), .ZN(n400) );
  XNOR2_X1 U468 ( .A(n400), .B(KEYINPUT26), .ZN(n577) );
  NOR2_X1 U469 ( .A1(n577), .A2(n401), .ZN(n402) );
  NOR2_X1 U470 ( .A1(n403), .A2(n402), .ZN(n404) );
  NOR2_X1 U471 ( .A1(n405), .A2(n404), .ZN(n406) );
  NOR2_X1 U472 ( .A1(n407), .A2(n406), .ZN(n480) );
  XOR2_X1 U473 ( .A(KEYINPUT72), .B(KEYINPUT10), .Z(n409) );
  XNOR2_X1 U474 ( .A(KEYINPUT9), .B(KEYINPUT65), .ZN(n408) );
  XNOR2_X1 U475 ( .A(n409), .B(n408), .ZN(n425) );
  XNOR2_X1 U476 ( .A(n411), .B(n410), .ZN(n416) );
  XNOR2_X1 U477 ( .A(KEYINPUT11), .B(KEYINPUT66), .ZN(n413) );
  AND2_X1 U478 ( .A1(G232GAT), .A2(G233GAT), .ZN(n412) );
  XNOR2_X1 U479 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U480 ( .A(n414), .B(KEYINPUT67), .Z(n415) );
  XNOR2_X1 U481 ( .A(n416), .B(n415), .ZN(n423) );
  XNOR2_X1 U482 ( .A(n418), .B(n417), .ZN(n421) );
  XNOR2_X1 U483 ( .A(n425), .B(n424), .ZN(n551) );
  XNOR2_X1 U484 ( .A(n476), .B(KEYINPUT36), .ZN(n576) );
  XOR2_X1 U485 ( .A(G64GAT), .B(G211GAT), .Z(n427) );
  XNOR2_X1 U486 ( .A(G127GAT), .B(G155GAT), .ZN(n426) );
  XNOR2_X1 U487 ( .A(n427), .B(n426), .ZN(n442) );
  XOR2_X1 U488 ( .A(n428), .B(G71GAT), .Z(n431) );
  XNOR2_X1 U489 ( .A(n429), .B(G183GAT), .ZN(n430) );
  XNOR2_X1 U490 ( .A(n431), .B(n430), .ZN(n435) );
  XOR2_X1 U491 ( .A(KEYINPUT76), .B(KEYINPUT12), .Z(n433) );
  NAND2_X1 U492 ( .A1(G231GAT), .A2(G233GAT), .ZN(n432) );
  XNOR2_X1 U493 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U494 ( .A(n435), .B(n434), .Z(n440) );
  XOR2_X1 U495 ( .A(KEYINPUT75), .B(KEYINPUT74), .Z(n437) );
  XNOR2_X1 U496 ( .A(G57GAT), .B(KEYINPUT15), .ZN(n436) );
  XNOR2_X1 U497 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U498 ( .A(n438), .B(KEYINPUT14), .ZN(n439) );
  XNOR2_X1 U499 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U500 ( .A(n442), .B(n441), .Z(n573) );
  INV_X1 U501 ( .A(n573), .ZN(n547) );
  OR2_X1 U502 ( .A1(n480), .A2(n444), .ZN(n445) );
  XNOR2_X1 U503 ( .A(n446), .B(n445), .ZN(n489) );
  NAND2_X1 U504 ( .A1(n504), .A2(n489), .ZN(n447) );
  XOR2_X1 U505 ( .A(KEYINPUT113), .B(n447), .Z(n518) );
  NOR2_X1 U506 ( .A1(n514), .A2(n518), .ZN(n450) );
  XNOR2_X1 U507 ( .A(n450), .B(n449), .ZN(G1339GAT) );
  NOR2_X1 U508 ( .A1(n576), .A2(n547), .ZN(n451) );
  XNOR2_X1 U509 ( .A(n451), .B(KEYINPUT45), .ZN(n453) );
  INV_X1 U510 ( .A(n570), .ZN(n452) );
  NAND2_X1 U511 ( .A1(n453), .A2(n452), .ZN(n454) );
  XNOR2_X1 U512 ( .A(n454), .B(KEYINPUT115), .ZN(n455) );
  AND2_X1 U513 ( .A1(n455), .A2(n540), .ZN(n456) );
  XNOR2_X1 U514 ( .A(n456), .B(KEYINPUT116), .ZN(n462) );
  NAND2_X1 U515 ( .A1(n551), .A2(n547), .ZN(n459) );
  NOR2_X1 U516 ( .A1(n540), .A2(n544), .ZN(n457) );
  XNOR2_X1 U517 ( .A(n457), .B(KEYINPUT46), .ZN(n458) );
  NOR2_X1 U518 ( .A1(n459), .A2(n458), .ZN(n460) );
  XOR2_X1 U519 ( .A(KEYINPUT47), .B(n460), .Z(n461) );
  NOR2_X1 U520 ( .A1(n462), .A2(n461), .ZN(n463) );
  XNOR2_X1 U521 ( .A(n463), .B(KEYINPUT48), .ZN(n536) );
  XNOR2_X1 U522 ( .A(KEYINPUT122), .B(n519), .ZN(n464) );
  NOR2_X1 U523 ( .A1(n536), .A2(n464), .ZN(n465) );
  XNOR2_X1 U524 ( .A(KEYINPUT54), .B(n465), .ZN(n566) );
  INV_X1 U525 ( .A(n466), .ZN(n467) );
  AND2_X1 U526 ( .A1(n565), .A2(n467), .ZN(n468) );
  AND2_X1 U527 ( .A1(n566), .A2(n468), .ZN(n469) );
  XNOR2_X1 U528 ( .A(n469), .B(KEYINPUT55), .ZN(n470) );
  INV_X1 U529 ( .A(n476), .ZN(n531) );
  NAND2_X1 U530 ( .A1(n560), .A2(n531), .ZN(n472) );
  INV_X1 U531 ( .A(G99GAT), .ZN(n475) );
  NOR2_X1 U532 ( .A1(n521), .A2(n518), .ZN(n473) );
  XNOR2_X1 U533 ( .A(KEYINPUT114), .B(n473), .ZN(n474) );
  XNOR2_X1 U534 ( .A(n475), .B(n474), .ZN(G1338GAT) );
  NOR2_X1 U535 ( .A1(n540), .A2(n570), .ZN(n488) );
  XOR2_X1 U536 ( .A(KEYINPUT16), .B(KEYINPUT77), .Z(n478) );
  NAND2_X1 U537 ( .A1(n573), .A2(n476), .ZN(n477) );
  XNOR2_X1 U538 ( .A(n478), .B(n477), .ZN(n479) );
  NOR2_X1 U539 ( .A1(n480), .A2(n479), .ZN(n505) );
  NAND2_X1 U540 ( .A1(n488), .A2(n505), .ZN(n486) );
  NOR2_X1 U541 ( .A1(n565), .A2(n486), .ZN(n481) );
  XOR2_X1 U542 ( .A(KEYINPUT34), .B(n481), .Z(n482) );
  XNOR2_X1 U543 ( .A(G1GAT), .B(n482), .ZN(G1324GAT) );
  NOR2_X1 U544 ( .A1(n519), .A2(n486), .ZN(n483) );
  XOR2_X1 U545 ( .A(G8GAT), .B(n483), .Z(G1325GAT) );
  NOR2_X1 U546 ( .A1(n521), .A2(n486), .ZN(n485) );
  XNOR2_X1 U547 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n484) );
  XNOR2_X1 U548 ( .A(n485), .B(n484), .ZN(G1326GAT) );
  NOR2_X1 U549 ( .A1(n514), .A2(n486), .ZN(n487) );
  XOR2_X1 U550 ( .A(G22GAT), .B(n487), .Z(G1327GAT) );
  XNOR2_X1 U551 ( .A(KEYINPUT101), .B(KEYINPUT39), .ZN(n492) );
  NAND2_X1 U552 ( .A1(n489), .A2(n488), .ZN(n490) );
  XNOR2_X1 U553 ( .A(n490), .B(KEYINPUT38), .ZN(n499) );
  NOR2_X1 U554 ( .A1(n565), .A2(n499), .ZN(n491) );
  XNOR2_X1 U555 ( .A(n492), .B(n491), .ZN(n493) );
  XOR2_X1 U556 ( .A(G29GAT), .B(n493), .Z(G1328GAT) );
  NOR2_X1 U557 ( .A1(n499), .A2(n519), .ZN(n495) );
  XNOR2_X1 U558 ( .A(G36GAT), .B(KEYINPUT103), .ZN(n494) );
  XNOR2_X1 U559 ( .A(n495), .B(n494), .ZN(G1329GAT) );
  NOR2_X1 U560 ( .A1(n499), .A2(n521), .ZN(n497) );
  XNOR2_X1 U561 ( .A(KEYINPUT104), .B(KEYINPUT40), .ZN(n496) );
  XNOR2_X1 U562 ( .A(n497), .B(n496), .ZN(n498) );
  XOR2_X1 U563 ( .A(G43GAT), .B(n498), .Z(G1330GAT) );
  XNOR2_X1 U564 ( .A(G50GAT), .B(KEYINPUT105), .ZN(n501) );
  NOR2_X1 U565 ( .A1(n514), .A2(n499), .ZN(n500) );
  XNOR2_X1 U566 ( .A(n501), .B(n500), .ZN(G1331GAT) );
  XOR2_X1 U567 ( .A(KEYINPUT109), .B(KEYINPUT110), .Z(n503) );
  XNOR2_X1 U568 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n502) );
  XNOR2_X1 U569 ( .A(n503), .B(n502), .ZN(n507) );
  NAND2_X1 U570 ( .A1(n505), .A2(n504), .ZN(n513) );
  NOR2_X1 U571 ( .A1(n565), .A2(n513), .ZN(n506) );
  XOR2_X1 U572 ( .A(n507), .B(n506), .Z(n508) );
  XNOR2_X1 U573 ( .A(KEYINPUT106), .B(n508), .ZN(G1332GAT) );
  NOR2_X1 U574 ( .A1(n519), .A2(n513), .ZN(n510) );
  XNOR2_X1 U575 ( .A(G64GAT), .B(KEYINPUT111), .ZN(n509) );
  XNOR2_X1 U576 ( .A(n510), .B(n509), .ZN(G1333GAT) );
  NOR2_X1 U577 ( .A1(n521), .A2(n513), .ZN(n511) );
  XOR2_X1 U578 ( .A(KEYINPUT112), .B(n511), .Z(n512) );
  XNOR2_X1 U579 ( .A(G71GAT), .B(n512), .ZN(G1334GAT) );
  NOR2_X1 U580 ( .A1(n514), .A2(n513), .ZN(n516) );
  XNOR2_X1 U581 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n515) );
  XNOR2_X1 U582 ( .A(n516), .B(n515), .ZN(G1335GAT) );
  NOR2_X1 U583 ( .A1(n518), .A2(n565), .ZN(n517) );
  XOR2_X1 U584 ( .A(G85GAT), .B(n517), .Z(G1336GAT) );
  NOR2_X1 U585 ( .A1(n519), .A2(n518), .ZN(n520) );
  XOR2_X1 U586 ( .A(G92GAT), .B(n520), .Z(G1337GAT) );
  INV_X1 U587 ( .A(n540), .ZN(n567) );
  NOR2_X1 U588 ( .A1(n521), .A2(n536), .ZN(n522) );
  NAND2_X1 U589 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U590 ( .A(KEYINPUT117), .B(n524), .ZN(n532) );
  NAND2_X1 U591 ( .A1(n567), .A2(n532), .ZN(n525) );
  XNOR2_X1 U592 ( .A(G113GAT), .B(n525), .ZN(G1340GAT) );
  XOR2_X1 U593 ( .A(KEYINPUT118), .B(KEYINPUT49), .Z(n527) );
  NAND2_X1 U594 ( .A1(n532), .A2(n557), .ZN(n526) );
  XNOR2_X1 U595 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U596 ( .A(G120GAT), .B(n528), .ZN(G1341GAT) );
  NAND2_X1 U597 ( .A1(n532), .A2(n573), .ZN(n529) );
  XNOR2_X1 U598 ( .A(n529), .B(KEYINPUT50), .ZN(n530) );
  XNOR2_X1 U599 ( .A(G127GAT), .B(n530), .ZN(G1342GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT51), .B(KEYINPUT119), .Z(n534) );
  NAND2_X1 U601 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U602 ( .A(n534), .B(n533), .ZN(n535) );
  XOR2_X1 U603 ( .A(G134GAT), .B(n535), .Z(G1343GAT) );
  INV_X1 U604 ( .A(n536), .ZN(n539) );
  NOR2_X1 U605 ( .A1(n577), .A2(n537), .ZN(n538) );
  NAND2_X1 U606 ( .A1(n539), .A2(n538), .ZN(n550) );
  NOR2_X1 U607 ( .A1(n540), .A2(n550), .ZN(n541) );
  XOR2_X1 U608 ( .A(G141GAT), .B(n541), .Z(G1344GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT52), .B(KEYINPUT53), .Z(n543) );
  XNOR2_X1 U610 ( .A(G148GAT), .B(KEYINPUT120), .ZN(n542) );
  XNOR2_X1 U611 ( .A(n543), .B(n542), .ZN(n546) );
  NOR2_X1 U612 ( .A1(n544), .A2(n550), .ZN(n545) );
  XOR2_X1 U613 ( .A(n546), .B(n545), .Z(G1345GAT) );
  NOR2_X1 U614 ( .A1(n547), .A2(n550), .ZN(n549) );
  XNOR2_X1 U615 ( .A(G155GAT), .B(KEYINPUT121), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n549), .B(n548), .ZN(G1346GAT) );
  NOR2_X1 U617 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U618 ( .A(G162GAT), .B(n552), .Z(G1347GAT) );
  NAND2_X1 U619 ( .A1(n567), .A2(n560), .ZN(n553) );
  XNOR2_X1 U620 ( .A(G169GAT), .B(n553), .ZN(G1348GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT57), .B(KEYINPUT124), .Z(n555) );
  XNOR2_X1 U622 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n554) );
  XNOR2_X1 U623 ( .A(n555), .B(n554), .ZN(n556) );
  XOR2_X1 U624 ( .A(KEYINPUT123), .B(n556), .Z(n559) );
  NAND2_X1 U625 ( .A1(n557), .A2(n560), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(G1349GAT) );
  XOR2_X1 U627 ( .A(G183GAT), .B(KEYINPUT125), .Z(n562) );
  NAND2_X1 U628 ( .A1(n560), .A2(n573), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(G1350GAT) );
  XNOR2_X1 U630 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n563), .B(KEYINPUT60), .ZN(n564) );
  XOR2_X1 U632 ( .A(KEYINPUT126), .B(n564), .Z(n569) );
  NAND2_X1 U633 ( .A1(n566), .A2(n565), .ZN(n579) );
  NOR2_X1 U634 ( .A1(n577), .A2(n579), .ZN(n574) );
  NAND2_X1 U635 ( .A1(n574), .A2(n567), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n569), .B(n568), .ZN(G1352GAT) );
  XOR2_X1 U637 ( .A(G204GAT), .B(KEYINPUT61), .Z(n572) );
  NAND2_X1 U638 ( .A1(n574), .A2(n570), .ZN(n571) );
  XNOR2_X1 U639 ( .A(n572), .B(n571), .ZN(G1353GAT) );
  NAND2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n575), .B(G211GAT), .ZN(G1354GAT) );
  OR2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n578) );
  NOR2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n581) );
  XNOR2_X1 U644 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U646 ( .A(n582), .B(G218GAT), .ZN(G1355GAT) );
endmodule

