//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 1 1 1 0 0 1 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 1 0 1 1 0 0 0 1 0 0 0 1 1 1 0 0 1 0 0 0 0 1 0 0 0 1 1 0 1 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n691, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n742, new_n744,
    new_n745, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n778, new_n779, new_n780, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n840, new_n841,
    new_n843, new_n844, new_n845, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n963, new_n964, new_n965, new_n966, new_n967;
  INV_X1    g000(.A(G15gat), .ZN(new_n202));
  INV_X1    g001(.A(G22gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(G15gat), .A2(G22gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT16), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n206), .B1(new_n207), .B2(G1gat), .ZN(new_n208));
  INV_X1    g007(.A(G1gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n204), .A2(new_n209), .A3(new_n205), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G8gat), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT85), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n212), .B1(new_n210), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n211), .A2(new_n214), .ZN(new_n215));
  OAI211_X1 g014(.A(new_n208), .B(new_n210), .C1(new_n213), .C2(new_n212), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  XNOR2_X1  g017(.A(G43gat), .B(G50gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(KEYINPUT15), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  NOR2_X1   g020(.A1(G29gat), .A2(G36gat), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT14), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g023(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n226), .A2(KEYINPUT84), .ZN(new_n227));
  NAND2_X1  g026(.A1(G29gat), .A2(G36gat), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT84), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n228), .B1(new_n224), .B2(new_n229), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n221), .B1(new_n227), .B2(new_n230), .ZN(new_n231));
  OR2_X1    g030(.A1(new_n219), .A2(KEYINPUT15), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n232), .A2(new_n220), .A3(new_n226), .A4(new_n228), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT17), .ZN(new_n234));
  AND3_X1   g033(.A1(new_n231), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n234), .B1(new_n231), .B2(new_n233), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n218), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n231), .A2(new_n233), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n217), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(G229gat), .A2(G233gat), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n237), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT18), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n217), .B(new_n238), .ZN(new_n244));
  XOR2_X1   g043(.A(new_n240), .B(KEYINPUT13), .Z(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n237), .A2(KEYINPUT18), .A3(new_n239), .A4(new_n240), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n243), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(KEYINPUT11), .B(G169gat), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n249), .B(G197gat), .ZN(new_n250));
  XOR2_X1   g049(.A(G113gat), .B(G141gat), .Z(new_n251));
  XNOR2_X1  g050(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n252), .B(KEYINPUT12), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n248), .A2(new_n254), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n243), .A2(new_n253), .A3(new_n246), .A4(new_n247), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(G78gat), .B(G106gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n258), .B(new_n203), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(G197gat), .B(G204gat), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT22), .ZN(new_n262));
  INV_X1    g061(.A(G211gat), .ZN(new_n263));
  INV_X1    g062(.A(G218gat), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n262), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n261), .A2(new_n265), .ZN(new_n266));
  XOR2_X1   g065(.A(G211gat), .B(G218gat), .Z(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT72), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n266), .A2(new_n267), .ZN(new_n271));
  NOR3_X1   g070(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  AND2_X1   g071(.A1(new_n261), .A2(new_n265), .ZN(new_n273));
  INV_X1    g072(.A(new_n267), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(KEYINPUT72), .B1(new_n275), .B2(new_n268), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n272), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(G141gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(G148gat), .ZN(new_n279));
  INV_X1    g078(.A(G148gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(G141gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT2), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT75), .ZN(new_n285));
  INV_X1    g084(.A(G155gat), .ZN(new_n286));
  INV_X1    g085(.A(G162gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(G155gat), .A2(G162gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n284), .A2(new_n285), .A3(new_n291), .ZN(new_n292));
  AOI21_X1  g091(.A(KEYINPUT2), .B1(new_n279), .B2(new_n281), .ZN(new_n293));
  OAI21_X1  g092(.A(KEYINPUT75), .B1(new_n293), .B2(new_n290), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n289), .B1(new_n288), .B2(KEYINPUT2), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n278), .A2(G148gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(KEYINPUT76), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT76), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n281), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n297), .A2(new_n279), .A3(new_n299), .ZN(new_n300));
  AOI22_X1  g099(.A1(new_n292), .A2(new_n294), .B1(new_n295), .B2(new_n300), .ZN(new_n301));
  XOR2_X1   g100(.A(KEYINPUT78), .B(KEYINPUT3), .Z(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  AOI21_X1  g102(.A(KEYINPUT29), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g103(.A(KEYINPUT81), .B1(new_n277), .B2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT81), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n270), .B1(new_n269), .B2(new_n271), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n275), .A2(KEYINPUT72), .A3(new_n268), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n300), .A2(new_n295), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n285), .B1(new_n284), .B2(new_n291), .ZN(new_n311));
  NOR3_X1   g110(.A1(new_n293), .A2(KEYINPUT75), .A3(new_n290), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n310), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n313), .A2(new_n302), .ZN(new_n314));
  OAI211_X1 g113(.A(new_n306), .B(new_n309), .C1(new_n314), .C2(KEYINPUT29), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n313), .A2(KEYINPUT3), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT29), .ZN(new_n317));
  OAI211_X1 g116(.A(new_n313), .B(new_n317), .C1(new_n271), .C2(new_n269), .ZN(new_n318));
  NAND4_X1  g117(.A1(new_n305), .A2(new_n315), .A3(new_n316), .A4(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n319), .A2(G228gat), .A3(G233gat), .ZN(new_n320));
  XNOR2_X1  g119(.A(KEYINPUT31), .B(G50gat), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n309), .B1(new_n314), .B2(KEYINPUT29), .ZN(new_n323));
  NAND2_X1  g122(.A1(G228gat), .A2(G233gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n313), .A2(new_n302), .ZN(new_n325));
  NAND4_X1  g124(.A1(new_n323), .A2(new_n324), .A3(new_n318), .A4(new_n325), .ZN(new_n326));
  AND3_X1   g125(.A1(new_n320), .A2(new_n322), .A3(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n322), .B1(new_n320), .B2(new_n326), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n260), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n320), .A2(new_n326), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(new_n321), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n320), .A2(new_n322), .A3(new_n326), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n331), .A2(new_n259), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n329), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(G227gat), .ZN(new_n335));
  INV_X1    g134(.A(G233gat), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  XOR2_X1   g136(.A(G127gat), .B(G134gat), .Z(new_n338));
  INV_X1    g137(.A(KEYINPUT70), .ZN(new_n339));
  INV_X1    g138(.A(G120gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(G113gat), .ZN(new_n341));
  INV_X1    g140(.A(G113gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(G120gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT1), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n339), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  AOI211_X1 g145(.A(KEYINPUT70), .B(KEYINPUT1), .C1(new_n341), .C2(new_n343), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n338), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n338), .ZN(new_n349));
  AOI21_X1  g148(.A(KEYINPUT1), .B1(new_n341), .B2(new_n343), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n349), .B1(new_n350), .B2(new_n339), .ZN(new_n351));
  XNOR2_X1  g150(.A(KEYINPUT67), .B(G190gat), .ZN(new_n352));
  XNOR2_X1  g151(.A(KEYINPUT27), .B(G183gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(KEYINPUT28), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT28), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n352), .A2(new_n353), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT26), .ZN(new_n359));
  INV_X1    g158(.A(G169gat), .ZN(new_n360));
  INV_X1    g159(.A(G176gat), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n359), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT68), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(G169gat), .A2(G176gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(new_n359), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n360), .A2(new_n361), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n359), .A2(new_n360), .A3(new_n361), .A4(KEYINPUT68), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n364), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(G183gat), .A2(G190gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(KEYINPUT69), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT69), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n370), .A2(new_n374), .A3(new_n371), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n358), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(G183gat), .ZN(new_n377));
  AND2_X1   g176(.A1(KEYINPUT67), .A2(G190gat), .ZN(new_n378));
  NOR2_X1   g177(.A1(KEYINPUT67), .A2(G190gat), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n377), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT24), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n371), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n380), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  AND2_X1   g183(.A1(new_n384), .A2(KEYINPUT25), .ZN(new_n385));
  OAI21_X1  g184(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(KEYINPUT23), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT23), .ZN(new_n388));
  OAI211_X1 g187(.A(new_n388), .B(KEYINPUT66), .C1(G169gat), .C2(G176gat), .ZN(new_n389));
  AND3_X1   g188(.A1(new_n387), .A2(new_n365), .A3(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT65), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n382), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n371), .A2(KEYINPUT65), .A3(new_n381), .ZN(new_n393));
  OR2_X1    g192(.A1(G183gat), .A2(G190gat), .ZN(new_n394));
  NAND4_X1  g193(.A1(new_n392), .A2(new_n393), .A3(new_n394), .A4(new_n383), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(new_n390), .ZN(new_n396));
  XOR2_X1   g195(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n397));
  AOI22_X1  g196(.A1(new_n385), .A2(new_n390), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  OAI211_X1 g197(.A(new_n348), .B(new_n351), .C1(new_n376), .C2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n358), .ZN(new_n400));
  INV_X1    g199(.A(new_n375), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n374), .B1(new_n370), .B2(new_n371), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n400), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n396), .A2(new_n397), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n390), .A2(new_n384), .A3(KEYINPUT25), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n348), .A2(new_n351), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n403), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n337), .B1(new_n399), .B2(new_n408), .ZN(new_n409));
  OR2_X1    g208(.A1(new_n409), .A2(KEYINPUT34), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(KEYINPUT34), .ZN(new_n411));
  AND2_X1   g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n399), .A2(new_n337), .A3(new_n408), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT33), .ZN(new_n414));
  XNOR2_X1  g213(.A(G15gat), .B(G43gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(G71gat), .B(G99gat), .ZN(new_n416));
  XOR2_X1   g215(.A(new_n415), .B(new_n416), .Z(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  OAI211_X1 g217(.A(new_n413), .B(KEYINPUT32), .C1(new_n414), .C2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n413), .A2(KEYINPUT32), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n413), .A2(new_n414), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n420), .A2(new_n421), .A3(new_n417), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n412), .A2(new_n419), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n419), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n410), .A2(new_n411), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n423), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT35), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n334), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  XOR2_X1   g228(.A(G8gat), .B(G36gat), .Z(new_n430));
  XNOR2_X1  g229(.A(new_n430), .B(G64gat), .ZN(new_n431));
  INV_X1    g230(.A(G92gat), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n431), .B(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(G226gat), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n435), .A2(new_n336), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n436), .A2(KEYINPUT29), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n438), .B1(new_n376), .B2(new_n398), .ZN(new_n439));
  INV_X1    g238(.A(new_n436), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n403), .A2(new_n406), .A3(new_n440), .ZN(new_n441));
  AND3_X1   g240(.A1(new_n439), .A2(new_n309), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n309), .B1(new_n439), .B2(new_n441), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n434), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT30), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n445), .A2(KEYINPUT74), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n445), .A2(KEYINPUT74), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n444), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT5), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n407), .A2(new_n313), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n292), .A2(new_n294), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n452), .A2(new_n348), .A3(new_n310), .A4(new_n351), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(G225gat), .A2(G233gat), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n450), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT77), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT3), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n458), .B1(new_n301), .B2(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n313), .A2(KEYINPUT77), .A3(KEYINPUT3), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n301), .A2(new_n303), .ZN(new_n462));
  AND4_X1   g261(.A1(new_n460), .A2(new_n461), .A3(new_n407), .A4(new_n462), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n301), .A2(KEYINPUT4), .A3(new_n348), .A4(new_n351), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n407), .A2(new_n313), .ZN(new_n465));
  XOR2_X1   g264(.A(KEYINPUT79), .B(KEYINPUT4), .Z(new_n466));
  OAI211_X1 g265(.A(new_n455), .B(new_n464), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n457), .B1(new_n463), .B2(new_n467), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n460), .A2(new_n461), .A3(new_n407), .A4(new_n462), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n456), .A2(KEYINPUT5), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT4), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n453), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n465), .A2(new_n466), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n469), .A2(new_n470), .A3(new_n472), .A4(new_n473), .ZN(new_n474));
  XNOR2_X1  g273(.A(KEYINPUT0), .B(G57gat), .ZN(new_n475));
  XNOR2_X1  g274(.A(new_n475), .B(G85gat), .ZN(new_n476));
  XNOR2_X1  g275(.A(G1gat), .B(G29gat), .ZN(new_n477));
  XOR2_X1   g276(.A(new_n476), .B(new_n477), .Z(new_n478));
  NAND3_X1  g277(.A1(new_n468), .A2(new_n474), .A3(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT6), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n478), .B1(new_n468), .B2(new_n474), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n468), .A2(new_n474), .ZN(new_n484));
  INV_X1    g283(.A(new_n478), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n484), .A2(KEYINPUT6), .A3(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n449), .B1(new_n483), .B2(new_n487), .ZN(new_n488));
  OAI211_X1 g287(.A(KEYINPUT30), .B(new_n434), .C1(new_n442), .C2(new_n443), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n439), .A2(new_n441), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(new_n277), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n439), .A2(new_n441), .A3(new_n309), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n491), .A2(new_n433), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  NOR3_X1   g293(.A1(new_n429), .A2(new_n488), .A3(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT80), .ZN(new_n496));
  AND3_X1   g295(.A1(new_n489), .A2(KEYINPUT73), .A3(new_n493), .ZN(new_n497));
  AOI21_X1  g296(.A(KEYINPUT73), .B1(new_n489), .B2(new_n493), .ZN(new_n498));
  OR2_X1    g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n496), .B1(new_n488), .B2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(new_n449), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n484), .A2(new_n485), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n502), .A2(new_n480), .A3(new_n479), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n501), .B1(new_n503), .B2(new_n486), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n497), .A2(new_n498), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n504), .A2(KEYINPUT80), .A3(new_n505), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n412), .A2(KEYINPUT71), .A3(new_n419), .A4(new_n422), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT71), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n424), .B1(new_n508), .B2(new_n425), .ZN(new_n509));
  AOI22_X1  g308(.A1(new_n333), .A2(new_n329), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n500), .A2(new_n506), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n495), .B1(KEYINPUT35), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n334), .ZN(new_n513));
  AND3_X1   g312(.A1(new_n504), .A2(KEYINPUT80), .A3(new_n505), .ZN(new_n514));
  AOI21_X1  g313(.A(KEYINPUT80), .B1(new_n504), .B2(new_n505), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT36), .ZN(new_n517));
  AND3_X1   g316(.A1(new_n423), .A2(new_n426), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n517), .B1(new_n507), .B2(new_n509), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(KEYINPUT83), .B(KEYINPUT38), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  NOR3_X1   g322(.A1(new_n442), .A2(new_n443), .A3(KEYINPUT37), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT37), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n525), .B1(new_n491), .B2(new_n492), .ZN(new_n526));
  OAI211_X1 g325(.A(new_n433), .B(new_n523), .C1(new_n524), .C2(new_n526), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n503), .A2(new_n527), .A3(new_n486), .A4(new_n444), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n433), .B1(new_n524), .B2(new_n526), .ZN(new_n529));
  AND2_X1   g328(.A1(new_n529), .A2(new_n522), .ZN(new_n530));
  OR2_X1    g329(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n494), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(new_n449), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT82), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n534), .A2(KEYINPUT40), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n469), .A2(new_n472), .A3(new_n473), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(new_n456), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n451), .A2(new_n455), .A3(new_n453), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n537), .A2(KEYINPUT39), .A3(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n478), .B1(new_n537), .B2(KEYINPUT39), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n535), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  OR2_X1    g341(.A1(new_n537), .A2(KEYINPUT39), .ZN(new_n543));
  INV_X1    g342(.A(new_n535), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n543), .A2(new_n478), .A3(new_n544), .A4(new_n539), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n533), .A2(new_n542), .A3(new_n502), .A4(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n531), .A2(new_n334), .A3(new_n546), .ZN(new_n547));
  AND3_X1   g346(.A1(new_n516), .A2(new_n521), .A3(new_n547), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n257), .B1(new_n512), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(KEYINPUT86), .ZN(new_n550));
  NAND2_X1  g349(.A1(G230gat), .A2(G233gat), .ZN(new_n551));
  INV_X1    g350(.A(G85gat), .ZN(new_n552));
  OAI21_X1  g351(.A(KEYINPUT91), .B1(new_n552), .B2(new_n432), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT91), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n554), .A2(G85gat), .A3(G92gat), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n553), .A2(new_n555), .A3(KEYINPUT7), .ZN(new_n556));
  NAND2_X1  g355(.A1(G99gat), .A2(G106gat), .ZN(new_n557));
  AOI22_X1  g356(.A1(KEYINPUT8), .A2(new_n557), .B1(new_n552), .B2(new_n432), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT7), .ZN(new_n559));
  OAI211_X1 g358(.A(KEYINPUT91), .B(new_n559), .C1(new_n552), .C2(new_n432), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n556), .A2(new_n558), .A3(new_n560), .ZN(new_n561));
  XOR2_X1   g360(.A(G99gat), .B(G106gat), .Z(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n562), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n564), .A2(new_n558), .A3(new_n556), .A4(new_n560), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(G57gat), .B(G64gat), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  OR2_X1    g367(.A1(G71gat), .A2(G78gat), .ZN(new_n569));
  NAND2_X1  g368(.A1(G71gat), .A2(G78gat), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT9), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n568), .A2(new_n571), .A3(new_n573), .ZN(new_n574));
  OAI211_X1 g373(.A(new_n570), .B(new_n569), .C1(new_n567), .C2(new_n572), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n566), .A2(new_n576), .ZN(new_n577));
  AND2_X1   g376(.A1(new_n574), .A2(new_n575), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n578), .A2(new_n563), .A3(new_n565), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n551), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(G176gat), .B(G204gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(G148gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(KEYINPUT95), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(G120gat), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT10), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n577), .A2(new_n586), .A3(new_n579), .ZN(new_n587));
  NAND4_X1  g386(.A1(new_n578), .A2(new_n563), .A3(KEYINPUT10), .A4(new_n565), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(KEYINPUT94), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT94), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n587), .A2(new_n588), .A3(new_n591), .ZN(new_n592));
  AND2_X1   g391(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n551), .ZN(new_n594));
  OAI211_X1 g393(.A(new_n581), .B(new_n585), .C1(new_n593), .C2(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n594), .B1(new_n587), .B2(new_n588), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n596), .A2(new_n580), .ZN(new_n597));
  OR2_X1    g396(.A1(new_n597), .A2(new_n585), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT86), .ZN(new_n601));
  OAI211_X1 g400(.A(new_n601), .B(new_n257), .C1(new_n512), .C2(new_n548), .ZN(new_n602));
  AND3_X1   g401(.A1(new_n550), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G134gat), .B(G162gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(KEYINPUT90), .ZN(new_n605));
  AOI21_X1  g404(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n606));
  XOR2_X1   g405(.A(new_n606), .B(KEYINPUT89), .Z(new_n607));
  XNOR2_X1  g406(.A(new_n605), .B(new_n607), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n566), .B1(new_n235), .B2(new_n236), .ZN(new_n609));
  NAND3_X1  g408(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n610));
  INV_X1    g409(.A(new_n238), .ZN(new_n611));
  OAI211_X1 g410(.A(new_n609), .B(new_n610), .C1(new_n566), .C2(new_n611), .ZN(new_n612));
  XOR2_X1   g411(.A(G190gat), .B(G218gat), .Z(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(KEYINPUT92), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n608), .B1(new_n615), .B2(KEYINPUT93), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n612), .B(new_n614), .ZN(new_n617));
  OR2_X1    g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n616), .A2(new_n617), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n217), .B1(KEYINPUT21), .B2(new_n578), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(new_n263), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n578), .A2(KEYINPUT21), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(G127gat), .B(G155gat), .ZN(new_n626));
  XOR2_X1   g425(.A(new_n626), .B(KEYINPUT20), .Z(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  OR2_X1    g427(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(G231gat), .A2(G233gat), .ZN(new_n630));
  XOR2_X1   g429(.A(new_n630), .B(KEYINPUT87), .Z(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(KEYINPUT19), .ZN(new_n632));
  XOR2_X1   g431(.A(KEYINPUT88), .B(G183gat), .Z(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n625), .A2(new_n628), .ZN(new_n635));
  AND3_X1   g434(.A1(new_n629), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n634), .B1(new_n629), .B2(new_n635), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n621), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n603), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n483), .A2(new_n487), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(KEYINPUT96), .B(G1gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(G1324gat));
  INV_X1    g444(.A(new_n640), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n646), .A2(new_n533), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT97), .ZN(new_n648));
  XNOR2_X1  g447(.A(KEYINPUT16), .B(G8gat), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n647), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n649), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n651), .B1(KEYINPUT97), .B2(KEYINPUT42), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT42), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n653), .B1(new_n647), .B2(G8gat), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n646), .A2(new_n533), .A3(new_n651), .ZN(new_n655));
  AOI22_X1  g454(.A1(new_n650), .A2(new_n652), .B1(new_n654), .B2(new_n655), .ZN(G1325gat));
  NOR3_X1   g455(.A1(new_n640), .A2(new_n202), .A3(new_n521), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n646), .A2(new_n427), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n657), .B1(new_n202), .B2(new_n658), .ZN(G1326gat));
  NOR2_X1   g458(.A1(new_n640), .A2(new_n334), .ZN(new_n660));
  XOR2_X1   g459(.A(KEYINPUT43), .B(G22gat), .Z(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT98), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n660), .B(new_n662), .ZN(G1327gat));
  OAI211_X1 g462(.A(KEYINPUT44), .B(new_n620), .C1(new_n512), .C2(new_n548), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n636), .A2(new_n637), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n257), .ZN(new_n667));
  NOR3_X1   g466(.A1(new_n666), .A2(new_n599), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n516), .A2(KEYINPUT99), .ZN(new_n669));
  AND2_X1   g468(.A1(new_n546), .A2(new_n334), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n520), .B1(new_n531), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n500), .A2(new_n506), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT99), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n672), .A2(new_n673), .A3(new_n513), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n669), .A2(new_n671), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n511), .A2(KEYINPUT35), .ZN(new_n676));
  OR2_X1    g475(.A1(new_n429), .A2(new_n488), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n676), .B1(new_n494), .B2(new_n677), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n621), .B1(new_n675), .B2(new_n678), .ZN(new_n679));
  OAI211_X1 g478(.A(new_n664), .B(new_n668), .C1(new_n679), .C2(KEYINPUT44), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT100), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n680), .B(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(G29gat), .B1(new_n682), .B2(new_n642), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n666), .A2(new_n599), .ZN(new_n684));
  NAND4_X1  g483(.A1(new_n550), .A2(new_n602), .A3(new_n620), .A4(new_n684), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n685), .A2(G29gat), .A3(new_n642), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT45), .ZN(new_n687));
  AND2_X1   g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n686), .A2(new_n687), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n683), .B1(new_n688), .B2(new_n689), .ZN(G1328gat));
  INV_X1    g489(.A(new_n533), .ZN(new_n691));
  NOR3_X1   g490(.A1(new_n685), .A2(G36gat), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(KEYINPUT46), .ZN(new_n693));
  OAI21_X1  g492(.A(G36gat), .B1(new_n682), .B2(new_n691), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(G1329gat));
  INV_X1    g494(.A(KEYINPUT101), .ZN(new_n696));
  OAI211_X1 g495(.A(new_n696), .B(G43gat), .C1(new_n682), .C2(new_n521), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n673), .B1(new_n672), .B2(new_n513), .ZN(new_n699));
  AOI211_X1 g498(.A(KEYINPUT99), .B(new_n334), .C1(new_n500), .C2(new_n506), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n512), .B1(new_n701), .B2(new_n671), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n698), .B1(new_n702), .B2(new_n621), .ZN(new_n703));
  NAND4_X1  g502(.A1(new_n703), .A2(new_n681), .A3(new_n664), .A4(new_n668), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n680), .A2(KEYINPUT100), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n521), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(G43gat), .ZN(new_n707));
  OAI21_X1  g506(.A(KEYINPUT101), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(new_n427), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n709), .A2(G43gat), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  OR3_X1    g510(.A1(new_n685), .A2(KEYINPUT102), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(KEYINPUT102), .B1(new_n685), .B2(new_n711), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n697), .A2(new_n708), .A3(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT47), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(G43gat), .B1(new_n680), .B2(new_n521), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n714), .A2(KEYINPUT47), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n717), .A2(new_n719), .ZN(G1330gat));
  NOR3_X1   g519(.A1(new_n685), .A2(G50gat), .A3(new_n334), .ZN(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  OAI21_X1  g521(.A(G50gat), .B1(new_n680), .B2(new_n334), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n722), .A2(KEYINPUT48), .A3(new_n723), .ZN(new_n724));
  OR2_X1    g523(.A1(new_n682), .A2(new_n334), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n721), .B1(new_n725), .B2(G50gat), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n724), .B1(new_n726), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR3_X1   g526(.A1(new_n702), .A2(new_n638), .A3(new_n257), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(new_n599), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(new_n641), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g531(.A(new_n533), .B(KEYINPUT103), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n729), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g534(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n736));
  AND2_X1   g535(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n735), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n738), .B1(new_n735), .B2(new_n736), .ZN(G1333gat));
  NAND3_X1  g538(.A1(new_n730), .A2(G71gat), .A3(new_n520), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n729), .A2(new_n709), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n740), .B1(G71gat), .B2(new_n741), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g542(.A1(new_n729), .A2(new_n334), .ZN(new_n744));
  XOR2_X1   g543(.A(KEYINPUT104), .B(G78gat), .Z(new_n745));
  XNOR2_X1  g544(.A(new_n744), .B(new_n745), .ZN(G1335gat));
  NOR2_X1   g545(.A1(new_n666), .A2(new_n257), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n703), .A2(new_n599), .A3(new_n664), .A4(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(G85gat), .B1(new_n748), .B2(new_n642), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n675), .A2(new_n678), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n750), .A2(new_n620), .A3(new_n747), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT51), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n679), .A2(KEYINPUT51), .A3(new_n747), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n641), .A2(new_n552), .A3(new_n599), .ZN(new_n757));
  XOR2_X1   g556(.A(new_n757), .B(KEYINPUT105), .Z(new_n758));
  OAI21_X1  g557(.A(new_n749), .B1(new_n756), .B2(new_n758), .ZN(G1336gat));
  OR3_X1    g558(.A1(new_n748), .A2(KEYINPUT108), .A3(new_n734), .ZN(new_n760));
  OAI21_X1  g559(.A(KEYINPUT108), .B1(new_n748), .B2(new_n734), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n760), .A2(G92gat), .A3(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT52), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n734), .A2(G92gat), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n751), .A2(new_n752), .ZN(new_n765));
  AOI21_X1  g564(.A(KEYINPUT51), .B1(new_n679), .B2(new_n747), .ZN(new_n766));
  OAI211_X1 g565(.A(new_n599), .B(new_n764), .C1(new_n765), .C2(new_n766), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n762), .A2(new_n763), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(KEYINPUT106), .ZN(new_n769));
  OAI21_X1  g568(.A(G92gat), .B1(new_n748), .B2(new_n691), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT106), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n755), .A2(new_n771), .A3(new_n599), .A4(new_n764), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n769), .A2(new_n770), .A3(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT107), .ZN(new_n774));
  AND3_X1   g573(.A1(new_n773), .A2(new_n774), .A3(KEYINPUT52), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n774), .B1(new_n773), .B2(KEYINPUT52), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n768), .B1(new_n775), .B2(new_n776), .ZN(G1337gat));
  INV_X1    g576(.A(G99gat), .ZN(new_n778));
  NOR3_X1   g577(.A1(new_n748), .A2(new_n778), .A3(new_n521), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n755), .A2(new_n599), .A3(new_n427), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n779), .B1(new_n778), .B2(new_n780), .ZN(G1338gat));
  INV_X1    g580(.A(KEYINPUT110), .ZN(new_n782));
  OAI21_X1  g581(.A(G106gat), .B1(new_n748), .B2(new_n334), .ZN(new_n783));
  INV_X1    g582(.A(G106gat), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n755), .A2(new_n784), .A3(new_n599), .A4(new_n513), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n782), .B1(new_n783), .B2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n785), .A2(KEYINPUT109), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n783), .A2(new_n785), .A3(new_n782), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n787), .A2(KEYINPUT53), .A3(new_n788), .A4(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n788), .A2(KEYINPUT53), .ZN(new_n791));
  INV_X1    g590(.A(new_n789), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n791), .B1(new_n792), .B2(new_n786), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n790), .A2(new_n793), .ZN(G1339gat));
  INV_X1    g593(.A(KEYINPUT54), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n585), .B1(new_n596), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n594), .B1(new_n590), .B2(new_n592), .ZN(new_n797));
  OAI21_X1  g596(.A(KEYINPUT54), .B1(new_n589), .B2(new_n551), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n796), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT55), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  OAI211_X1 g600(.A(new_n796), .B(KEYINPUT55), .C1(new_n797), .C2(new_n798), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n801), .A2(new_n257), .A3(new_n595), .A4(new_n802), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n244), .A2(new_n245), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n240), .B1(new_n237), .B2(new_n239), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n252), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n256), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n599), .A2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT111), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n803), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n809), .B1(new_n803), .B2(new_n808), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n811), .A2(new_n812), .A3(new_n620), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n801), .A2(new_n802), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n814), .A2(new_n620), .A3(new_n595), .A4(new_n807), .ZN(new_n815));
  INV_X1    g614(.A(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n665), .B1(new_n813), .B2(new_n816), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n638), .A2(new_n599), .A3(new_n257), .ZN(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n817), .A2(KEYINPUT112), .A3(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT112), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n803), .A2(new_n808), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(KEYINPUT111), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n823), .A2(new_n621), .A3(new_n810), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n666), .B1(new_n824), .B2(new_n815), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n821), .B1(new_n825), .B2(new_n818), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n820), .A2(new_n826), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n827), .A2(new_n641), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n828), .A2(new_n510), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n829), .A2(new_n734), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n257), .A2(new_n342), .ZN(new_n831));
  XNOR2_X1  g630(.A(new_n831), .B(KEYINPUT113), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n513), .A2(new_n709), .ZN(new_n834));
  AND2_X1   g633(.A1(new_n827), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n733), .A2(new_n642), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(G113gat), .B1(new_n837), .B2(new_n667), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n833), .A2(new_n838), .ZN(G1340gat));
  NAND3_X1  g638(.A1(new_n830), .A2(new_n340), .A3(new_n599), .ZN(new_n840));
  OAI21_X1  g639(.A(G120gat), .B1(new_n837), .B2(new_n600), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(G1341gat));
  AOI21_X1  g641(.A(G127gat), .B1(new_n830), .B2(new_n666), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n835), .A2(G127gat), .A3(new_n666), .A4(new_n836), .ZN(new_n844));
  XNOR2_X1  g643(.A(new_n844), .B(KEYINPUT114), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n843), .A2(new_n845), .ZN(G1342gat));
  INV_X1    g645(.A(G134gat), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n620), .A2(new_n691), .ZN(new_n848));
  XNOR2_X1  g647(.A(new_n848), .B(KEYINPUT115), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n829), .A2(new_n847), .A3(new_n849), .ZN(new_n850));
  OR2_X1    g649(.A1(new_n850), .A2(KEYINPUT56), .ZN(new_n851));
  OAI21_X1  g650(.A(G134gat), .B1(new_n837), .B2(new_n621), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n850), .A2(KEYINPUT56), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(G1343gat));
  NAND3_X1  g653(.A1(new_n820), .A2(new_n826), .A3(new_n513), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT57), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT116), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n855), .A2(KEYINPUT116), .A3(new_n856), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n822), .A2(new_n621), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n815), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n862), .A2(new_n665), .ZN(new_n863));
  OAI211_X1 g662(.A(KEYINPUT57), .B(new_n513), .C1(new_n863), .C2(new_n818), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n859), .A2(new_n860), .A3(new_n864), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n520), .A2(new_n733), .A3(new_n642), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n865), .A2(new_n257), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(G141gat), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n520), .A2(new_n334), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n828), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n870), .A2(new_n733), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n871), .A2(new_n278), .A3(new_n257), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n868), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(KEYINPUT58), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT58), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n868), .A2(new_n872), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n874), .A2(new_n876), .ZN(G1344gat));
  INV_X1    g676(.A(KEYINPUT59), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n865), .A2(new_n866), .ZN(new_n879));
  OAI211_X1 g678(.A(new_n878), .B(G148gat), .C1(new_n879), .C2(new_n600), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n855), .A2(KEYINPUT57), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n862), .A2(KEYINPUT118), .ZN(new_n882));
  OR2_X1    g681(.A1(new_n862), .A2(KEYINPUT118), .ZN(new_n883));
  AND3_X1   g682(.A1(new_n882), .A2(new_n665), .A3(new_n883), .ZN(new_n884));
  OAI211_X1 g683(.A(new_n856), .B(new_n513), .C1(new_n884), .C2(new_n818), .ZN(new_n885));
  AND3_X1   g684(.A1(new_n881), .A2(new_n599), .A3(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT117), .ZN(new_n887));
  OR2_X1    g686(.A1(new_n866), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n866), .A2(new_n887), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n886), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n890), .A2(G148gat), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n880), .B1(new_n891), .B2(new_n878), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n871), .A2(new_n280), .A3(new_n599), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(G1345gat));
  NOR3_X1   g693(.A1(new_n879), .A2(new_n286), .A3(new_n665), .ZN(new_n895));
  AOI21_X1  g694(.A(G155gat), .B1(new_n871), .B2(new_n666), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n895), .A2(new_n896), .ZN(G1346gat));
  INV_X1    g696(.A(KEYINPUT119), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n898), .B1(new_n879), .B2(new_n621), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n865), .A2(KEYINPUT119), .A3(new_n620), .A4(new_n866), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n899), .A2(G162gat), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n849), .A2(new_n287), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n901), .B1(new_n870), .B2(new_n902), .ZN(G1347gat));
  AND2_X1   g702(.A1(new_n827), .A2(new_n642), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n733), .A2(new_n510), .ZN(new_n905));
  XNOR2_X1  g704(.A(new_n905), .B(KEYINPUT120), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n907), .A2(new_n360), .A3(new_n257), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n641), .A2(new_n691), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n827), .A2(new_n834), .A3(new_n909), .ZN(new_n910));
  OAI21_X1  g709(.A(G169gat), .B1(new_n910), .B2(new_n667), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n908), .A2(new_n911), .ZN(G1348gat));
  NOR3_X1   g711(.A1(new_n910), .A2(new_n361), .A3(new_n600), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n907), .A2(new_n599), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n913), .B1(new_n914), .B2(new_n361), .ZN(G1349gat));
  NOR2_X1   g714(.A1(KEYINPUT122), .A2(KEYINPUT60), .ZN(new_n916));
  AND2_X1   g715(.A1(KEYINPUT122), .A2(KEYINPUT60), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n907), .A2(new_n666), .A3(new_n353), .ZN(new_n918));
  NAND4_X1  g717(.A1(new_n835), .A2(KEYINPUT121), .A3(new_n666), .A4(new_n909), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT121), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n920), .B1(new_n910), .B2(new_n665), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n919), .A2(G183gat), .A3(new_n921), .ZN(new_n922));
  AOI211_X1 g721(.A(new_n916), .B(new_n917), .C1(new_n918), .C2(new_n922), .ZN(new_n923));
  AND4_X1   g722(.A1(KEYINPUT122), .A2(new_n918), .A3(new_n922), .A4(KEYINPUT60), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n923), .A2(new_n924), .ZN(G1350gat));
  NAND3_X1  g724(.A1(new_n907), .A2(new_n620), .A3(new_n352), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT123), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n926), .B(new_n927), .ZN(new_n928));
  OAI21_X1  g727(.A(G190gat), .B1(new_n910), .B2(new_n621), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n929), .B(KEYINPUT61), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n928), .A2(new_n930), .ZN(G1351gat));
  AND2_X1   g730(.A1(new_n904), .A2(new_n733), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n932), .A2(new_n869), .ZN(new_n933));
  INV_X1    g732(.A(G197gat), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n933), .A2(new_n934), .A3(new_n257), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n521), .A2(new_n909), .ZN(new_n936));
  INV_X1    g735(.A(new_n936), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n881), .A2(new_n885), .A3(new_n937), .ZN(new_n938));
  OAI21_X1  g737(.A(G197gat), .B1(new_n938), .B2(new_n667), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n935), .A2(new_n939), .ZN(G1352gat));
  INV_X1    g739(.A(G204gat), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n933), .A2(new_n941), .A3(new_n599), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(KEYINPUT62), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT62), .ZN(new_n944));
  NAND4_X1  g743(.A1(new_n933), .A2(new_n944), .A3(new_n941), .A4(new_n599), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n886), .A2(new_n937), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(G204gat), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n943), .A2(new_n945), .A3(new_n947), .ZN(G1353gat));
  NAND4_X1  g747(.A1(new_n881), .A2(new_n885), .A3(new_n666), .A4(new_n937), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT125), .ZN(new_n950));
  OR2_X1    g749(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n949), .A2(new_n950), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n951), .A2(G211gat), .A3(new_n952), .ZN(new_n953));
  OR2_X1    g752(.A1(new_n953), .A2(KEYINPUT63), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(KEYINPUT63), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n665), .A2(G211gat), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n932), .A2(new_n869), .A3(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT124), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND4_X1  g758(.A1(new_n932), .A2(KEYINPUT124), .A3(new_n869), .A4(new_n956), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n954), .A2(new_n955), .A3(new_n961), .ZN(G1354gat));
  NAND3_X1  g761(.A1(new_n933), .A2(new_n264), .A3(new_n620), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT126), .ZN(new_n964));
  AND2_X1   g763(.A1(new_n938), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n620), .B1(new_n938), .B2(new_n964), .ZN(new_n966));
  OAI21_X1  g765(.A(G218gat), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n963), .A2(new_n967), .ZN(G1355gat));
endmodule


