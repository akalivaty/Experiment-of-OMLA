//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 1 0 0 0 1 1 1 0 0 0 1 1 0 1 0 1 0 1 0 1 1 0 1 1 0 0 0 1 0 0 1 1 0 0 0 0 1 0 1 1 0 0 1 0 0 0 0 0 0 1 0 1 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:06 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1290, new_n1291, new_n1292, new_n1293, new_n1294,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1315, new_n1316, new_n1317, new_n1318, new_n1319,
    new_n1320, new_n1321, new_n1322, new_n1323, new_n1325, new_n1326,
    new_n1327, new_n1328, new_n1330, new_n1331, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1379, new_n1380, new_n1381, new_n1382, new_n1383,
    new_n1384, new_n1385, new_n1386;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n208), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  OR2_X1    g0018(.A1(new_n218), .A2(KEYINPUT1), .ZN(new_n219));
  OR2_X1    g0019(.A1(new_n202), .A2(KEYINPUT64), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n202), .A2(KEYINPUT64), .ZN(new_n221));
  NAND3_X1  g0021(.A1(new_n220), .A2(G50), .A3(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n224), .A2(new_n206), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  NAND3_X1  g0026(.A1(new_n211), .A2(new_n219), .A3(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n218), .ZN(G361));
  XOR2_X1   g0028(.A(G238), .B(G244), .Z(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G226), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n233), .B(new_n236), .Z(G358));
  XNOR2_X1  g0037(.A(G50), .B(G68), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G58), .B(G77), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n238), .B(new_n239), .Z(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XOR2_X1   g0041(.A(G107), .B(G116), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G351));
  NAND3_X1  g0044(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n245), .A2(new_n224), .ZN(new_n246));
  INV_X1    g0046(.A(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(KEYINPUT8), .B(G58), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n206), .A2(G33), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  NOR2_X1   g0051(.A1(G20), .A2(G33), .ZN(new_n252));
  AOI22_X1  g0052(.A1(new_n249), .A2(new_n251), .B1(G150), .B2(new_n252), .ZN(new_n253));
  OAI21_X1  g0053(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n247), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  OR2_X1    g0055(.A1(new_n255), .A2(KEYINPUT67), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(KEYINPUT67), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n259), .A2(new_n246), .ZN(new_n260));
  INV_X1    g0060(.A(G50), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n261), .B1(new_n205), .B2(G20), .ZN(new_n262));
  AOI22_X1  g0062(.A1(new_n260), .A2(new_n262), .B1(new_n261), .B2(new_n259), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n256), .A2(new_n257), .A3(new_n263), .ZN(new_n264));
  XNOR2_X1  g0064(.A(new_n264), .B(KEYINPUT9), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT3), .ZN(new_n266));
  INV_X1    g0066(.A(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(KEYINPUT3), .A2(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G1698), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n270), .A2(G222), .A3(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G77), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n270), .A2(G1698), .ZN(new_n274));
  INV_X1    g0074(.A(G223), .ZN(new_n275));
  OAI221_X1 g0075(.A(new_n272), .B1(new_n273), .B2(new_n270), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(G33), .A2(G41), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n277), .A2(G1), .A3(G13), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G41), .ZN(new_n281));
  INV_X1    g0081(.A(G45), .ZN(new_n282));
  AOI21_X1  g0082(.A(G1), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n283), .A2(new_n278), .A3(G274), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n279), .A2(new_n283), .ZN(new_n286));
  XNOR2_X1  g0086(.A(KEYINPUT66), .B(G226), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n285), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n280), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G200), .ZN(new_n290));
  INV_X1    g0090(.A(G190), .ZN(new_n291));
  OAI211_X1 g0091(.A(new_n265), .B(new_n290), .C1(new_n291), .C2(new_n289), .ZN(new_n292));
  XNOR2_X1  g0092(.A(new_n292), .B(KEYINPUT10), .ZN(new_n293));
  INV_X1    g0093(.A(G179), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n280), .A2(new_n294), .A3(new_n288), .ZN(new_n295));
  INV_X1    g0095(.A(G169), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n289), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n264), .A2(new_n295), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n293), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n275), .A2(new_n271), .ZN(new_n300));
  INV_X1    g0100(.A(G226), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G1698), .ZN(new_n302));
  AND2_X1   g0102(.A1(KEYINPUT3), .A2(G33), .ZN(new_n303));
  NOR2_X1   g0103(.A1(KEYINPUT3), .A2(G33), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n300), .B(new_n302), .C1(new_n303), .C2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(G33), .A2(G87), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n278), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n278), .A2(G232), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n284), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n308), .A2(new_n312), .A3(new_n294), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n296), .B1(new_n307), .B2(new_n311), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n303), .A2(new_n304), .ZN(new_n316));
  AOI21_X1  g0116(.A(KEYINPUT7), .B1(new_n316), .B2(new_n206), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n268), .A2(KEYINPUT7), .A3(new_n206), .A4(new_n269), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(G68), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  AND2_X1   g0120(.A1(G58), .A2(G68), .ZN(new_n321));
  OAI21_X1  g0121(.A(G20), .B1(new_n321), .B2(new_n201), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n252), .A2(G159), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n322), .A2(KEYINPUT16), .A3(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n247), .B1(new_n320), .B2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT16), .ZN(new_n327));
  INV_X1    g0127(.A(G68), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n268), .A2(new_n206), .A3(new_n269), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT7), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n328), .B1(new_n331), .B2(new_n318), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n322), .A2(new_n323), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n327), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n326), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n248), .B1(new_n205), .B2(G20), .ZN(new_n336));
  AOI22_X1  g0136(.A1(new_n336), .A2(new_n260), .B1(new_n259), .B2(new_n248), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n315), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  XNOR2_X1  g0138(.A(new_n338), .B(KEYINPUT18), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT73), .ZN(new_n340));
  INV_X1    g0140(.A(new_n333), .ZN(new_n341));
  AOI21_X1  g0141(.A(KEYINPUT16), .B1(new_n320), .B2(new_n341), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n246), .B1(new_n332), .B2(new_n324), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n337), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n308), .A2(new_n312), .A3(new_n291), .ZN(new_n345));
  INV_X1    g0145(.A(G200), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n346), .B1(new_n307), .B2(new_n311), .ZN(new_n347));
  AND2_X1   g0147(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n340), .B1(new_n344), .B2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n337), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n350), .B1(new_n326), .B2(new_n334), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n345), .A2(new_n347), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n351), .A2(KEYINPUT73), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n349), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(KEYINPUT17), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n344), .A2(new_n348), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n356), .A2(KEYINPUT17), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n339), .A2(new_n355), .A3(new_n358), .ZN(new_n359));
  OAI211_X1 g0159(.A(G232), .B(G1698), .C1(new_n303), .C2(new_n304), .ZN(new_n360));
  OAI211_X1 g0160(.A(G226), .B(new_n271), .C1(new_n303), .C2(new_n304), .ZN(new_n361));
  NAND2_X1  g0161(.A1(G33), .A2(G97), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n360), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n279), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n278), .A2(G238), .A3(new_n309), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n284), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n368), .A2(KEYINPUT69), .A3(KEYINPUT13), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT69), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n366), .B1(new_n279), .B2(new_n363), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT13), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n370), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n294), .B1(new_n371), .B2(new_n372), .ZN(new_n374));
  AND3_X1   g0174(.A1(new_n369), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  AND3_X1   g0175(.A1(new_n364), .A2(new_n372), .A3(new_n367), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n372), .B1(new_n364), .B2(new_n367), .ZN(new_n377));
  OAI21_X1  g0177(.A(G169), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT72), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(KEYINPUT14), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n380), .ZN(new_n382));
  OAI211_X1 g0182(.A(G169), .B(new_n382), .C1(new_n376), .C2(new_n377), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n375), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT71), .ZN(new_n385));
  OAI22_X1  g0185(.A1(new_n250), .A2(new_n273), .B1(new_n206), .B2(G68), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT70), .ZN(new_n387));
  INV_X1    g0187(.A(new_n252), .ZN(new_n388));
  OAI22_X1  g0188(.A1(new_n386), .A2(new_n387), .B1(new_n261), .B2(new_n388), .ZN(new_n389));
  AND2_X1   g0189(.A1(new_n386), .A2(new_n387), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n385), .B(new_n246), .C1(new_n389), .C2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n386), .A2(new_n387), .ZN(new_n393));
  OAI221_X1 g0193(.A(KEYINPUT70), .B1(new_n206), .B2(G68), .C1(new_n250), .C2(new_n273), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n393), .B(new_n394), .C1(new_n261), .C2(new_n388), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n385), .B1(new_n395), .B2(new_n246), .ZN(new_n396));
  OAI21_X1  g0196(.A(KEYINPUT11), .B1(new_n392), .B2(new_n396), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n246), .B1(new_n389), .B2(new_n390), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(KEYINPUT71), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT11), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n399), .A2(new_n400), .A3(new_n391), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT12), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n402), .B1(new_n259), .B2(new_n328), .ZN(new_n403));
  NOR3_X1   g0203(.A1(new_n258), .A2(KEYINPUT12), .A3(G68), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n328), .B1(new_n205), .B2(G20), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n405), .B1(new_n260), .B2(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n397), .A2(new_n401), .A3(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n384), .A2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n407), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n399), .A2(new_n391), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n412), .B1(new_n413), .B2(KEYINPUT11), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n368), .A2(KEYINPUT13), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n371), .A2(new_n372), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(G200), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n369), .A2(new_n373), .A3(G190), .A4(new_n416), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n414), .A2(new_n418), .A3(new_n419), .A4(new_n401), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n411), .A2(new_n420), .ZN(new_n421));
  XOR2_X1   g0221(.A(KEYINPUT15), .B(G87), .Z(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n423), .A2(new_n250), .ZN(new_n424));
  OAI22_X1  g0224(.A1(new_n248), .A2(new_n388), .B1(new_n206), .B2(new_n273), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n246), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n260), .ZN(new_n427));
  OAI21_X1  g0227(.A(G77), .B1(new_n206), .B2(G1), .ZN(new_n428));
  OAI221_X1 g0228(.A(new_n426), .B1(G77), .B2(new_n258), .C1(new_n427), .C2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n270), .A2(G232), .A3(new_n271), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n316), .A2(G107), .ZN(new_n431));
  INV_X1    g0231(.A(G238), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n430), .B(new_n431), .C1(new_n274), .C2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(new_n279), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT68), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n285), .B1(G244), .B2(new_n286), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n434), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n435), .B1(new_n434), .B2(new_n436), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n429), .B1(new_n440), .B2(G200), .ZN(new_n441));
  OAI21_X1  g0241(.A(G190), .B1(new_n438), .B2(new_n439), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n440), .A2(new_n296), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n294), .B1(new_n438), .B2(new_n439), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n444), .A2(new_n429), .A3(new_n445), .ZN(new_n446));
  AND2_X1   g0246(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  NOR4_X1   g0248(.A1(new_n299), .A2(new_n359), .A3(new_n421), .A4(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  XNOR2_X1  g0250(.A(KEYINPUT77), .B(KEYINPUT19), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n251), .A2(G97), .ZN(new_n452));
  AOI21_X1  g0252(.A(G20), .B1(new_n268), .B2(new_n269), .ZN(new_n453));
  AOI22_X1  g0253(.A1(new_n451), .A2(new_n452), .B1(new_n453), .B2(G68), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT78), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n455), .B(new_n206), .C1(new_n451), .C2(new_n362), .ZN(new_n456));
  NOR3_X1   g0256(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n362), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT77), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n461), .A2(KEYINPUT19), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT19), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n463), .A2(KEYINPUT77), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n460), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n455), .B1(new_n465), .B2(new_n206), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n454), .B1(new_n459), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(new_n246), .ZN(new_n468));
  OAI211_X1 g0268(.A(G244), .B(G1698), .C1(new_n303), .C2(new_n304), .ZN(new_n469));
  OAI211_X1 g0269(.A(G238), .B(new_n271), .C1(new_n303), .C2(new_n304), .ZN(new_n470));
  NAND2_X1  g0270(.A1(G33), .A2(G116), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(new_n279), .ZN(new_n473));
  INV_X1    g0273(.A(G274), .ZN(new_n474));
  AND2_X1   g0274(.A1(G1), .A2(G13), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n474), .B1(new_n475), .B2(new_n277), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n282), .A2(G1), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n205), .A2(G45), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n278), .A2(G250), .A3(new_n479), .ZN(new_n480));
  AND2_X1   g0280(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n473), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(G200), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n422), .A2(new_n258), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n205), .A2(G33), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n258), .A2(new_n486), .A3(new_n224), .A4(new_n245), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(G87), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n468), .A2(new_n483), .A3(new_n485), .A4(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(KEYINPUT80), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n484), .B1(new_n467), .B2(new_n246), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT80), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n492), .A2(new_n493), .A3(new_n483), .A4(new_n489), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n478), .A2(new_n480), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n495), .B1(new_n279), .B2(new_n472), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(G190), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n491), .A2(new_n494), .A3(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(G97), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n259), .A2(new_n499), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n500), .B1(new_n487), .B2(new_n499), .ZN(new_n501));
  XNOR2_X1  g0301(.A(G97), .B(G107), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT6), .ZN(new_n503));
  INV_X1    g0303(.A(G107), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n503), .A2(new_n499), .ZN(new_n505));
  AOI22_X1  g0305(.A1(new_n502), .A2(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  OAI22_X1  g0306(.A1(new_n506), .A2(new_n206), .B1(new_n273), .B2(new_n388), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n504), .B1(new_n331), .B2(new_n318), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n246), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(KEYINPUT74), .ZN(new_n510));
  OAI21_X1  g0310(.A(G107), .B1(new_n317), .B2(new_n319), .ZN(new_n511));
  AND2_X1   g0311(.A1(G97), .A2(G107), .ZN(new_n512));
  NOR2_X1   g0312(.A1(G97), .A2(G107), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n503), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n504), .A2(KEYINPUT6), .A3(G97), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n516), .A2(G20), .B1(G77), .B2(new_n252), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n511), .A2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT74), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n518), .A2(new_n519), .A3(new_n246), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n501), .B1(new_n510), .B2(new_n520), .ZN(new_n521));
  XNOR2_X1  g0321(.A(KEYINPUT5), .B(G41), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n522), .A2(new_n477), .B1(new_n475), .B2(new_n277), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(G257), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n476), .A2(new_n477), .A3(new_n522), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  OAI211_X1 g0326(.A(G244), .B(new_n271), .C1(new_n303), .C2(new_n304), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT4), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT75), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n527), .A2(KEYINPUT75), .A3(new_n528), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n270), .A2(KEYINPUT4), .A3(G244), .A4(new_n271), .ZN(new_n533));
  OAI211_X1 g0333(.A(G250), .B(G1698), .C1(new_n303), .C2(new_n304), .ZN(new_n534));
  NAND2_X1  g0334(.A1(G33), .A2(G283), .ZN(new_n535));
  AND2_X1   g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n531), .A2(new_n532), .A3(new_n533), .A4(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n526), .B1(new_n537), .B2(new_n279), .ZN(new_n538));
  OAI21_X1  g0338(.A(KEYINPUT76), .B1(new_n538), .B2(new_n346), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT76), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n534), .B(new_n535), .C1(new_n527), .C2(new_n528), .ZN(new_n541));
  AOI21_X1  g0341(.A(KEYINPUT75), .B1(new_n527), .B2(new_n528), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n278), .B1(new_n543), .B2(new_n532), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n540), .B(G200), .C1(new_n544), .C2(new_n526), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n538), .A2(G190), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n521), .A2(new_n539), .A3(new_n545), .A4(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n488), .A2(new_n422), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n452), .A2(new_n451), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n453), .A2(G68), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n463), .A2(KEYINPUT77), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n461), .A2(KEYINPUT19), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(G20), .B1(new_n554), .B2(new_n460), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n457), .B1(new_n555), .B2(new_n455), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n465), .A2(new_n206), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(KEYINPUT78), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n551), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n485), .B(new_n548), .C1(new_n559), .C2(new_n247), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT79), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n492), .A2(KEYINPUT79), .A3(new_n548), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n496), .A2(G179), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n482), .A2(G169), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n562), .A2(new_n563), .A3(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n501), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n519), .B1(new_n518), .B2(new_n246), .ZN(new_n569));
  AOI211_X1 g0369(.A(KEYINPUT74), .B(new_n247), .C1(new_n511), .C2(new_n517), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n537), .A2(new_n279), .ZN(new_n572));
  INV_X1    g0372(.A(new_n526), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n296), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n538), .A2(new_n294), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n571), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n498), .A2(new_n547), .A3(new_n567), .A4(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n523), .A2(KEYINPUT81), .A3(G270), .ZN(new_n579));
  AND2_X1   g0379(.A1(KEYINPUT5), .A2(G41), .ZN(new_n580));
  NOR2_X1   g0380(.A1(KEYINPUT5), .A2(G41), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n477), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n582), .A2(G270), .A3(new_n278), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT81), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  OAI211_X1 g0385(.A(G264), .B(G1698), .C1(new_n303), .C2(new_n304), .ZN(new_n586));
  OAI211_X1 g0386(.A(G257), .B(new_n271), .C1(new_n303), .C2(new_n304), .ZN(new_n587));
  XOR2_X1   g0387(.A(KEYINPUT82), .B(G303), .Z(new_n588));
  OAI211_X1 g0388(.A(new_n586), .B(new_n587), .C1(new_n588), .C2(new_n270), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n579), .A2(new_n585), .B1(new_n279), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n590), .A2(G179), .A3(new_n525), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n589), .A2(new_n279), .ZN(new_n592));
  AOI21_X1  g0392(.A(KEYINPUT81), .B1(new_n523), .B2(G270), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n583), .A2(new_n584), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n592), .B(new_n525), .C1(new_n593), .C2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(G169), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT21), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n591), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT83), .ZN(new_n599));
  INV_X1    g0399(.A(G116), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n245), .A2(new_n224), .B1(G20), .B2(new_n600), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n535), .B(new_n206), .C1(G33), .C2(new_n499), .ZN(new_n602));
  AND3_X1   g0402(.A1(new_n601), .A2(KEYINPUT20), .A3(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(KEYINPUT20), .B1(new_n601), .B2(new_n602), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(G13), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n606), .A2(G1), .ZN(new_n607));
  AOI21_X1  g0407(.A(G116), .B1(new_n607), .B2(G20), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n608), .B1(G116), .B2(new_n487), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n599), .B1(new_n605), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n600), .A2(G20), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n602), .A2(new_n246), .A3(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT20), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n601), .A2(KEYINPUT20), .A3(new_n602), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n258), .A2(new_n600), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n617), .B1(new_n488), .B2(new_n600), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n616), .A2(new_n618), .A3(KEYINPUT83), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n610), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n598), .A2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n620), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n595), .A2(G200), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n622), .B(new_n623), .C1(new_n291), .C2(new_n595), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n296), .B1(new_n590), .B2(new_n525), .ZN(new_n625));
  AOI211_X1 g0425(.A(KEYINPUT84), .B(KEYINPUT21), .C1(new_n625), .C2(new_n620), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT84), .ZN(new_n627));
  NOR3_X1   g0427(.A1(new_n605), .A2(new_n599), .A3(new_n609), .ZN(new_n628));
  AOI21_X1  g0428(.A(KEYINPUT83), .B1(new_n616), .B2(new_n618), .ZN(new_n629));
  OAI211_X1 g0429(.A(G169), .B(new_n595), .C1(new_n628), .C2(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n627), .B1(new_n630), .B2(new_n597), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n621), .B(new_n624), .C1(new_n626), .C2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT23), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n633), .B1(new_n206), .B2(G107), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n504), .A2(KEYINPUT23), .A3(G20), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n206), .A2(G33), .A3(G116), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT22), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n640), .B1(new_n453), .B2(G87), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n206), .B(G87), .C1(new_n303), .C2(new_n304), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n642), .A2(KEYINPUT22), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n639), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  XNOR2_X1  g0444(.A(KEYINPUT85), .B(KEYINPUT24), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n644), .A2(KEYINPUT86), .A3(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n645), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n642), .A2(KEYINPUT22), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n270), .A2(new_n640), .A3(new_n206), .A4(G87), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n638), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT86), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n647), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  AOI211_X1 g0452(.A(KEYINPUT86), .B(new_n638), .C1(new_n648), .C2(new_n649), .ZN(new_n653));
  OAI211_X1 g0453(.A(new_n646), .B(new_n246), .C1(new_n652), .C2(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n259), .A2(KEYINPUT25), .A3(new_n504), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT25), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n656), .B1(new_n258), .B2(G107), .ZN(new_n657));
  AOI22_X1  g0457(.A1(G107), .A2(new_n488), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n654), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n582), .A2(G264), .A3(new_n278), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n660), .A2(new_n525), .ZN(new_n661));
  OAI211_X1 g0461(.A(G257), .B(G1698), .C1(new_n303), .C2(new_n304), .ZN(new_n662));
  OAI211_X1 g0462(.A(G250), .B(new_n271), .C1(new_n303), .C2(new_n304), .ZN(new_n663));
  INV_X1    g0463(.A(G294), .ZN(new_n664));
  OAI211_X1 g0464(.A(new_n662), .B(new_n663), .C1(new_n267), .C2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(new_n279), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n661), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n667), .A2(G179), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n668), .B1(new_n296), .B2(new_n667), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n659), .A2(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(G200), .B1(new_n661), .B2(new_n666), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT87), .ZN(new_n672));
  OAI22_X1  g0472(.A1(new_n671), .A2(new_n672), .B1(new_n667), .B2(G190), .ZN(new_n673));
  AOI211_X1 g0473(.A(KEYINPUT87), .B(G200), .C1(new_n661), .C2(new_n666), .ZN(new_n674));
  OAI211_X1 g0474(.A(new_n654), .B(new_n658), .C1(new_n673), .C2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n670), .A2(new_n675), .ZN(new_n676));
  NOR4_X1   g0476(.A1(new_n450), .A2(new_n578), .A3(new_n632), .A4(new_n676), .ZN(G372));
  INV_X1    g0477(.A(new_n298), .ZN(new_n678));
  INV_X1    g0478(.A(new_n446), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n410), .B1(new_n420), .B2(new_n679), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n357), .B1(KEYINPUT17), .B2(new_n354), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n339), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n678), .B1(new_n293), .B2(new_n683), .ZN(new_n684));
  AND2_X1   g0484(.A1(new_n547), .A2(new_n577), .ZN(new_n685));
  OAI211_X1 g0485(.A(new_n621), .B(new_n670), .C1(new_n626), .C2(new_n631), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n560), .A2(new_n566), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n492), .A2(new_n483), .A3(new_n489), .A4(new_n497), .ZN(new_n688));
  AND3_X1   g0488(.A1(new_n675), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n685), .A2(new_n686), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n687), .A2(new_n688), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n691), .B1(new_n577), .B2(KEYINPUT88), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT88), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n571), .A2(new_n575), .A3(new_n693), .A4(new_n576), .ZN(new_n694));
  AOI21_X1  g0494(.A(KEYINPUT26), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n538), .A2(G169), .ZN(new_n696));
  NOR3_X1   g0496(.A1(new_n544), .A2(G179), .A3(new_n526), .ZN(new_n697));
  NOR3_X1   g0497(.A1(new_n521), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  AND4_X1   g0498(.A1(KEYINPUT26), .A2(new_n498), .A3(new_n698), .A4(new_n567), .ZN(new_n699));
  OAI211_X1 g0499(.A(new_n690), .B(new_n687), .C1(new_n695), .C2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n684), .B1(new_n450), .B2(new_n701), .ZN(G369));
  NAND2_X1  g0502(.A1(new_n607), .A2(new_n206), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(KEYINPUT27), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT89), .ZN(new_n705));
  XNOR2_X1  g0505(.A(new_n704), .B(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(G213), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n707), .B1(new_n703), .B2(KEYINPUT27), .ZN(new_n708));
  AND3_X1   g0508(.A1(new_n706), .A2(G343), .A3(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n622), .A2(new_n710), .ZN(new_n711));
  OR2_X1    g0511(.A1(new_n632), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n621), .B1(new_n626), .B2(new_n631), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(new_n711), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(G330), .ZN(new_n716));
  XNOR2_X1  g0516(.A(new_n716), .B(KEYINPUT90), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n670), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(new_n709), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n659), .A2(new_n709), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n670), .A2(new_n721), .A3(new_n675), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n718), .A2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n670), .A2(new_n675), .A3(new_n710), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(new_n713), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n729), .B1(new_n670), .B2(new_n709), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n726), .A2(new_n731), .ZN(G399));
  INV_X1    g0532(.A(new_n209), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n733), .A2(G41), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n458), .A2(G116), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n735), .A2(G1), .A3(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n737), .B1(new_n222), .B2(new_n735), .ZN(new_n738));
  XNOR2_X1  g0538(.A(new_n738), .B(KEYINPUT28), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n701), .A2(new_n709), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT29), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n577), .A2(KEYINPUT88), .ZN(new_n743));
  INV_X1    g0543(.A(new_n691), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n743), .A2(new_n744), .A3(new_n694), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(KEYINPUT26), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT26), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n498), .A2(new_n698), .A3(new_n747), .A4(new_n567), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n746), .A2(new_n690), .A3(new_n687), .A4(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(new_n710), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(KEYINPUT29), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n742), .A2(new_n751), .ZN(new_n752));
  NOR3_X1   g0552(.A1(new_n578), .A2(new_n632), .A3(new_n727), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT30), .ZN(new_n754));
  AND3_X1   g0554(.A1(new_n473), .A2(new_n481), .A3(G179), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n755), .A2(new_n590), .A3(new_n666), .A4(new_n661), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n754), .B1(new_n756), .B2(new_n574), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n496), .A2(G179), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n574), .A2(new_n595), .A3(new_n667), .A4(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n579), .A2(new_n585), .ZN(new_n760));
  AND4_X1   g0560(.A1(new_n760), .A2(new_n592), .A3(new_n666), .A4(new_n661), .ZN(new_n761));
  NAND4_X1  g0561(.A1(new_n761), .A2(KEYINPUT30), .A3(new_n538), .A4(new_n755), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n757), .A2(new_n759), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(new_n709), .ZN(new_n764));
  INV_X1    g0564(.A(KEYINPUT31), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n763), .A2(KEYINPUT31), .A3(new_n709), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(G330), .B1(new_n753), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(KEYINPUT91), .ZN(new_n770));
  INV_X1    g0570(.A(new_n578), .ZN(new_n771));
  INV_X1    g0571(.A(new_n632), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n771), .A2(new_n772), .A3(new_n728), .ZN(new_n773));
  INV_X1    g0573(.A(new_n767), .ZN(new_n774));
  AOI21_X1  g0574(.A(KEYINPUT31), .B1(new_n763), .B2(new_n709), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n773), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(KEYINPUT91), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n777), .A2(new_n778), .A3(G330), .ZN(new_n779));
  AND2_X1   g0579(.A1(new_n770), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n752), .A2(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n739), .B1(new_n781), .B2(G1), .ZN(G364));
  NOR2_X1   g0582(.A1(new_n606), .A2(G20), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n205), .B1(new_n783), .B2(G45), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n734), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  OAI211_X1 g0587(.A(new_n718), .B(new_n787), .C1(G330), .C2(new_n715), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n209), .A2(new_n270), .ZN(new_n789));
  INV_X1    g0589(.A(G355), .ZN(new_n790));
  OAI22_X1  g0590(.A1(new_n789), .A2(new_n790), .B1(G116), .B2(new_n209), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n733), .A2(new_n270), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n793), .B1(new_n223), .B2(new_n282), .ZN(new_n794));
  OR2_X1    g0594(.A1(new_n240), .A2(new_n282), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n791), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(G13), .A2(G33), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(G20), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n224), .B1(G20), .B2(new_n296), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n786), .B1(new_n796), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n294), .A2(new_n346), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n804), .B(KEYINPUT93), .ZN(new_n805));
  OAI21_X1  g0605(.A(KEYINPUT92), .B1(new_n206), .B2(G190), .ZN(new_n806));
  OR3_X1    g0606(.A1(new_n206), .A2(KEYINPUT92), .A3(G190), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n805), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  OR2_X1    g0609(.A1(new_n809), .A2(KEYINPUT95), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n809), .A2(KEYINPUT95), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(G329), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n206), .A2(new_n294), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(G200), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n816), .A2(new_n291), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(G326), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n816), .A2(G190), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  XOR2_X1   g0620(.A(KEYINPUT33), .B(G317), .Z(new_n821));
  OAI21_X1  g0621(.A(new_n818), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n815), .A2(new_n291), .A3(new_n346), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n346), .A2(G179), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n825), .A2(G20), .A3(G190), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  AOI22_X1  g0627(.A1(G311), .A2(new_n824), .B1(new_n827), .B2(G303), .ZN(new_n828));
  INV_X1    g0628(.A(G322), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n815), .A2(G190), .A3(new_n346), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n828), .B(new_n316), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n807), .A2(new_n806), .A3(new_n825), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n822), .B(new_n831), .C1(G283), .C2(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n805), .A2(G190), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(G20), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  OAI211_X1 g0637(.A(new_n814), .B(new_n834), .C1(new_n664), .C2(new_n837), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n836), .A2(G97), .B1(G68), .B2(new_n819), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n839), .B(KEYINPUT94), .ZN(new_n840));
  INV_X1    g0640(.A(G159), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n808), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n842), .B(KEYINPUT32), .ZN(new_n843));
  INV_X1    g0643(.A(new_n830), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n316), .B1(new_n844), .B2(G58), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n827), .A2(G87), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n845), .B(new_n846), .C1(new_n273), .C2(new_n823), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n847), .B1(G50), .B2(new_n817), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n843), .B(new_n848), .C1(new_n504), .C2(new_n832), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n838), .B1(new_n840), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n803), .B1(new_n850), .B2(new_n800), .ZN(new_n851));
  INV_X1    g0651(.A(new_n799), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n851), .B1(new_n715), .B2(new_n852), .ZN(new_n853));
  AND2_X1   g0653(.A1(new_n788), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(G396));
  INV_X1    g0655(.A(new_n780), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n447), .A2(new_n710), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n700), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n444), .A2(new_n445), .A3(new_n429), .A4(new_n710), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  AOI22_X1  g0661(.A1(new_n441), .A2(new_n442), .B1(new_n429), .B2(new_n709), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n861), .B1(new_n863), .B2(new_n446), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n859), .B1(new_n740), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n786), .B1(new_n856), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n866), .B1(new_n856), .B2(new_n865), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n800), .A2(new_n797), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n787), .B1(new_n273), .B2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n800), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n817), .A2(G303), .ZN(new_n871));
  INV_X1    g0671(.A(G283), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n871), .B1(new_n820), .B2(new_n872), .ZN(new_n873));
  AOI22_X1  g0673(.A1(G116), .A2(new_n824), .B1(new_n827), .B2(G107), .ZN(new_n874));
  OAI211_X1 g0674(.A(new_n874), .B(new_n316), .C1(new_n664), .C2(new_n830), .ZN(new_n875));
  AOI211_X1 g0675(.A(new_n873), .B(new_n875), .C1(G87), .C2(new_n833), .ZN(new_n876));
  INV_X1    g0676(.A(G311), .ZN(new_n877));
  OAI221_X1 g0677(.A(new_n876), .B1(new_n499), .B2(new_n837), .C1(new_n877), .C2(new_n812), .ZN(new_n878));
  AOI22_X1  g0678(.A1(G143), .A2(new_n844), .B1(new_n824), .B2(G159), .ZN(new_n879));
  INV_X1    g0679(.A(G137), .ZN(new_n880));
  INV_X1    g0680(.A(new_n817), .ZN(new_n881));
  INV_X1    g0681(.A(G150), .ZN(new_n882));
  OAI221_X1 g0682(.A(new_n879), .B1(new_n880), .B2(new_n881), .C1(new_n882), .C2(new_n820), .ZN(new_n883));
  XNOR2_X1  g0683(.A(new_n883), .B(KEYINPUT34), .ZN(new_n884));
  OAI221_X1 g0684(.A(new_n270), .B1(new_n826), .B2(new_n261), .C1(new_n832), .C2(new_n328), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n885), .B1(G58), .B2(new_n836), .ZN(new_n886));
  INV_X1    g0686(.A(G132), .ZN(new_n887));
  OAI211_X1 g0687(.A(new_n884), .B(new_n886), .C1(new_n887), .C2(new_n812), .ZN(new_n888));
  AND2_X1   g0688(.A1(new_n878), .A2(new_n888), .ZN(new_n889));
  OAI221_X1 g0689(.A(new_n869), .B1(new_n870), .B2(new_n889), .C1(new_n864), .C2(new_n798), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n867), .A2(new_n890), .ZN(G384));
  NOR2_X1   g0691(.A1(new_n783), .A2(new_n205), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT38), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n706), .A2(new_n708), .ZN(new_n894));
  AOI22_X1  g0694(.A1(new_n335), .A2(new_n337), .B1(new_n315), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(KEYINPUT37), .B1(new_n354), .B2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n315), .ZN(new_n897));
  INV_X1    g0697(.A(new_n894), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n344), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT37), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n349), .A2(new_n899), .A3(new_n353), .A4(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n896), .A2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n344), .A2(new_n898), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n904), .B1(new_n681), .B2(new_n339), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n893), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n904), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n359), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n908), .A2(KEYINPUT38), .A3(new_n902), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n906), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n408), .A2(new_n709), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n420), .B(new_n911), .C1(new_n384), .C2(new_n409), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT97), .ZN(new_n913));
  NOR3_X1   g0713(.A1(new_n384), .A2(new_n911), .A3(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n373), .A2(new_n369), .A3(new_n374), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n382), .B1(new_n417), .B2(G169), .ZN(new_n916));
  INV_X1    g0716(.A(new_n383), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n915), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n710), .B1(new_n414), .B2(new_n401), .ZN(new_n919));
  AOI21_X1  g0719(.A(KEYINPUT97), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n912), .B1(new_n914), .B2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT98), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n913), .B1(new_n384), .B2(new_n911), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n918), .A2(KEYINPUT97), .A3(new_n919), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n926), .A2(KEYINPUT98), .A3(new_n912), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n923), .A2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT96), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n929), .B1(new_n859), .B2(new_n860), .ZN(new_n930));
  AOI211_X1 g0730(.A(KEYINPUT96), .B(new_n861), .C1(new_n700), .C2(new_n858), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n910), .B(new_n928), .C1(new_n930), .C2(new_n931), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n339), .A2(new_n898), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT39), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n910), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n901), .A2(KEYINPUT100), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n895), .A2(KEYINPUT37), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT100), .ZN(new_n940));
  NAND4_X1  g0740(.A1(new_n939), .A2(new_n940), .A3(new_n349), .A4(new_n353), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n938), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n344), .A2(new_n897), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n351), .A2(new_n352), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT99), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n904), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n945), .B1(new_n943), .B2(new_n944), .ZN(new_n948));
  OAI21_X1  g0748(.A(KEYINPUT37), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT101), .ZN(new_n950));
  AND3_X1   g0750(.A1(new_n942), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n950), .B1(new_n942), .B2(new_n949), .ZN(new_n952));
  NOR3_X1   g0752(.A1(new_n951), .A2(new_n952), .A3(new_n905), .ZN(new_n953));
  OAI21_X1  g0753(.A(KEYINPUT102), .B1(new_n953), .B2(KEYINPUT38), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT102), .ZN(new_n955));
  OAI21_X1  g0755(.A(KEYINPUT99), .B1(new_n356), .B2(new_n338), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n956), .A2(new_n904), .A3(new_n946), .ZN(new_n957));
  AOI22_X1  g0757(.A1(new_n938), .A2(new_n941), .B1(new_n957), .B2(KEYINPUT37), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n908), .B1(new_n958), .B2(new_n950), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n955), .B(new_n893), .C1(new_n959), .C2(new_n951), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n954), .A2(new_n909), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n937), .B1(new_n961), .B2(new_n936), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n411), .A2(new_n709), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n935), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n752), .A2(new_n449), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n684), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n964), .B(new_n966), .Z(new_n967));
  OAI21_X1  g0767(.A(new_n860), .B1(new_n862), .B2(new_n679), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n968), .B1(new_n773), .B2(new_n776), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n910), .A2(new_n928), .A3(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT40), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT103), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n970), .A2(KEYINPUT103), .A3(new_n971), .ZN(new_n975));
  AND4_X1   g0775(.A1(KEYINPUT40), .A2(new_n928), .A3(new_n777), .A4(new_n864), .ZN(new_n976));
  AOI22_X1  g0776(.A1(new_n974), .A2(new_n975), .B1(new_n961), .B2(new_n976), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n977), .A2(new_n449), .A3(new_n777), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(G330), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n977), .B1(new_n449), .B2(new_n777), .ZN(new_n980));
  OR2_X1    g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n892), .B1(new_n967), .B2(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n967), .B2(new_n981), .ZN(new_n983));
  OR2_X1    g0783(.A1(new_n516), .A2(KEYINPUT35), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n516), .A2(KEYINPUT35), .ZN(new_n985));
  NAND4_X1  g0785(.A1(new_n984), .A2(new_n985), .A3(G116), .A4(new_n225), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT36), .ZN(new_n987));
  NOR3_X1   g0787(.A1(new_n222), .A2(new_n273), .A3(new_n321), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n328), .A2(G50), .ZN(new_n989));
  OAI211_X1 g0789(.A(G1), .B(new_n606), .C1(new_n988), .C2(new_n989), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n983), .A2(new_n987), .A3(new_n990), .ZN(G367));
  NAND2_X1  g0791(.A1(new_n547), .A2(new_n577), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n521), .A2(new_n710), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n992), .A2(new_n993), .B1(new_n577), .B2(new_n710), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT104), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n994), .B(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n729), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n998), .B(KEYINPUT42), .Z(new_n999));
  AND2_X1   g0799(.A1(new_n996), .A2(new_n719), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n710), .B1(new_n1000), .B2(new_n698), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n492), .A2(new_n489), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(new_n709), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n744), .A2(new_n1003), .ZN(new_n1004));
  OR2_X1    g0804(.A1(new_n1003), .A2(new_n687), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n999), .A2(new_n1001), .B1(KEYINPUT43), .B2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1007), .B1(KEYINPUT43), .B2(new_n1006), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT43), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1006), .ZN(new_n1010));
  NAND4_X1  g0810(.A1(new_n999), .A2(new_n1009), .A3(new_n1010), .A4(new_n1001), .ZN(new_n1011));
  AND4_X1   g0811(.A1(new_n725), .A2(new_n1008), .A3(new_n996), .A4(new_n1011), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n1008), .A2(new_n1011), .B1(new_n725), .B2(new_n996), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n734), .B(KEYINPUT41), .Z(new_n1015));
  NAND2_X1  g0815(.A1(new_n996), .A2(new_n731), .ZN(new_n1016));
  XOR2_X1   g0816(.A(new_n1016), .B(KEYINPUT45), .Z(new_n1017));
  NOR2_X1   g0817(.A1(new_n996), .A2(new_n731), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT44), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(KEYINPUT105), .B1(new_n1020), .B2(new_n725), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n725), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n729), .A2(KEYINPUT106), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n713), .A2(new_n710), .ZN(new_n1025));
  AOI21_X1  g0825(.A(KEYINPUT106), .B1(new_n724), .B2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1024), .B1(new_n1026), .B2(new_n997), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n718), .A2(new_n1027), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n717), .B(new_n1024), .C1(new_n997), .C2(new_n1026), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n781), .ZN(new_n1031));
  OAI21_X1  g0831(.A(KEYINPUT107), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  AND2_X1   g0832(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT107), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1033), .A2(new_n1034), .A3(new_n781), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1020), .A2(KEYINPUT105), .A3(new_n725), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1023), .A2(new_n1032), .A3(new_n1035), .A4(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1015), .B1(new_n1037), .B2(new_n781), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1014), .B1(new_n1038), .B2(new_n785), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n792), .A2(new_n236), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1040), .B(new_n801), .C1(new_n209), .C2(new_n423), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n832), .A2(new_n499), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n270), .B1(new_n824), .B2(G283), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n1043), .B1(new_n588), .B2(new_n830), .C1(new_n877), .C2(new_n881), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n1042), .B(new_n1044), .C1(G317), .C2(new_n809), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n827), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT46), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n826), .B2(new_n600), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1046), .B(new_n1048), .C1(new_n820), .C2(new_n664), .ZN(new_n1049));
  XOR2_X1   g0849(.A(new_n1049), .B(KEYINPUT108), .Z(new_n1050));
  OAI211_X1 g0850(.A(new_n1045), .B(new_n1050), .C1(new_n504), .C2(new_n837), .ZN(new_n1051));
  XOR2_X1   g0851(.A(new_n1051), .B(KEYINPUT109), .Z(new_n1052));
  NOR2_X1   g0852(.A1(new_n832), .A2(new_n273), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n270), .B1(new_n261), .B2(new_n823), .C1(new_n820), .C2(new_n841), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n809), .A2(G137), .B1(G58), .B2(new_n827), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT111), .ZN(new_n1056));
  AOI211_X1 g0856(.A(new_n1053), .B(new_n1054), .C1(new_n1055), .C2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n1056), .B2(new_n1055), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n836), .A2(G68), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(G143), .A2(new_n817), .B1(new_n844), .B2(G150), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT110), .Z(new_n1062));
  OAI21_X1  g0862(.A(new_n1052), .B1(new_n1058), .B2(new_n1062), .ZN(new_n1063));
  XOR2_X1   g0863(.A(new_n1063), .B(KEYINPUT47), .Z(new_n1064));
  OAI211_X1 g0864(.A(new_n786), .B(new_n1041), .C1(new_n1064), .C2(new_n870), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1065), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n1066), .A2(KEYINPUT112), .B1(new_n799), .B2(new_n1010), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1067), .B1(KEYINPUT112), .B2(new_n1066), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1039), .A2(new_n1068), .ZN(G387));
  AND2_X1   g0869(.A1(new_n1035), .A2(new_n1032), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n734), .B1(new_n1033), .B2(new_n781), .ZN(new_n1071));
  OR2_X1    g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n789), .A2(new_n736), .B1(G107), .B2(new_n209), .ZN(new_n1073));
  OR2_X1    g0873(.A1(new_n233), .A2(new_n282), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n736), .ZN(new_n1075));
  AOI211_X1 g0875(.A(G45), .B(new_n1075), .C1(G68), .C2(G77), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n248), .A2(G50), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1077), .B(KEYINPUT50), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n793), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1073), .B1(new_n1074), .B2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n786), .B1(new_n1080), .B2(new_n802), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n836), .A2(new_n422), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1082), .B1(new_n261), .B2(new_n830), .ZN(new_n1083));
  XOR2_X1   g0883(.A(new_n1083), .B(KEYINPUT113), .Z(new_n1084));
  AOI22_X1  g0884(.A1(G159), .A2(new_n817), .B1(new_n819), .B2(new_n249), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n316), .B1(new_n824), .B2(G68), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1085), .B(new_n1086), .C1(new_n273), .C2(new_n826), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n808), .A2(new_n882), .ZN(new_n1088));
  OR4_X1    g0888(.A1(new_n1042), .A2(new_n1084), .A3(new_n1087), .A4(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n270), .B1(new_n809), .B2(G326), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n837), .A2(new_n872), .B1(new_n664), .B2(new_n826), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT48), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n588), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n1093), .A2(new_n824), .B1(new_n844), .B2(G317), .ZN(new_n1094));
  OAI221_X1 g0894(.A(new_n1094), .B1(new_n877), .B2(new_n820), .C1(new_n829), .C2(new_n881), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1091), .B1(new_n1092), .B2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1096), .B1(new_n1092), .B2(new_n1095), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT49), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n1090), .B1(new_n600), .B2(new_n832), .C1(new_n1097), .C2(new_n1098), .ZN(new_n1099));
  AND2_X1   g0899(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1089), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1081), .B1(new_n1101), .B2(new_n800), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1102), .B1(new_n723), .B2(new_n852), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(new_n1103), .B(KEYINPUT114), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(new_n1033), .B2(new_n785), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1072), .A2(new_n1105), .ZN(G393));
  XNOR2_X1  g0906(.A(new_n726), .B(new_n1020), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n785), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n792), .A2(new_n243), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n802), .B1(G97), .B2(new_n733), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n787), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n881), .A2(new_n882), .B1(new_n841), .B2(new_n830), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT51), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n826), .A2(new_n328), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n270), .B1(new_n823), .B2(new_n248), .ZN(new_n1115));
  AOI211_X1 g0915(.A(new_n1114), .B(new_n1115), .C1(G50), .C2(new_n819), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n836), .A2(G77), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n809), .A2(G143), .B1(G87), .B2(new_n833), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n1113), .A2(new_n1116), .A3(new_n1117), .A4(new_n1118), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n808), .A2(new_n829), .B1(new_n872), .B2(new_n826), .ZN(new_n1120));
  XOR2_X1   g0920(.A(new_n1120), .B(KEYINPUT115), .Z(new_n1121));
  AOI22_X1  g0921(.A1(G317), .A2(new_n817), .B1(new_n844), .B2(G311), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n1122), .B(KEYINPUT52), .ZN(new_n1123));
  OAI221_X1 g0923(.A(new_n316), .B1(new_n823), .B2(new_n664), .C1(new_n832), .C2(new_n504), .ZN(new_n1124));
  OR3_X1    g0924(.A1(new_n1121), .A2(new_n1123), .A3(new_n1124), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n836), .A2(G116), .B1(new_n1093), .B2(new_n819), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(new_n1126), .B(KEYINPUT116), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1119), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(new_n1128), .B(KEYINPUT117), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n1111), .B1(new_n996), .B2(new_n852), .C1(new_n870), .C2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1037), .A2(new_n734), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n1070), .A2(new_n1107), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n1108), .B(new_n1130), .C1(new_n1131), .C2(new_n1132), .ZN(G390));
  NAND3_X1  g0933(.A1(new_n770), .A2(new_n779), .A3(new_n864), .ZN(new_n1134));
  AND3_X1   g0934(.A1(new_n926), .A2(KEYINPUT98), .A3(new_n912), .ZN(new_n1135));
  AOI21_X1  g0935(.A(KEYINPUT98), .B1(new_n926), .B2(new_n912), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1134), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(G330), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n1139), .B(new_n968), .C1(new_n773), .C2(new_n776), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n928), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n859), .A2(new_n929), .A3(new_n860), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n745), .A2(new_n747), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n498), .A2(new_n698), .A3(new_n567), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1143), .B1(new_n1144), .B2(new_n747), .ZN(new_n1145));
  AND4_X1   g0945(.A1(new_n577), .A2(new_n744), .A3(new_n547), .A4(new_n675), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n1146), .A2(new_n686), .B1(new_n560), .B2(new_n566), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n857), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(KEYINPUT96), .B1(new_n1148), .B2(new_n861), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n1138), .A2(new_n1141), .B1(new_n1142), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n770), .A2(new_n779), .A3(new_n864), .A4(new_n928), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n863), .A2(new_n446), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n749), .A2(new_n710), .A3(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1154), .A2(new_n860), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  AND2_X1   g0956(.A1(new_n1152), .A2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g0957(.A(KEYINPUT118), .B1(new_n1140), .B2(new_n928), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT118), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n864), .B(G330), .C1(new_n753), .C2(new_n768), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1137), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1158), .A2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(KEYINPUT119), .B1(new_n1157), .B2(new_n1162), .ZN(new_n1163));
  AND3_X1   g0963(.A1(new_n1137), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1159), .B1(new_n1137), .B2(new_n1160), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n1152), .B(new_n1156), .C1(new_n1164), .C2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT119), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1151), .B1(new_n1163), .B2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n449), .A2(G330), .A3(new_n777), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n965), .A2(new_n684), .A3(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1169), .A2(KEYINPUT120), .A3(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1141), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n960), .A2(new_n909), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n942), .A2(new_n949), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(KEYINPUT101), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n958), .A2(new_n950), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1177), .A2(new_n1178), .A3(new_n908), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n955), .B1(new_n1179), .B2(new_n893), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n936), .B1(new_n1175), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n937), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n928), .B1(new_n930), .B2(new_n931), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n963), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n1181), .A2(new_n1182), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1155), .A2(new_n928), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1186), .B(new_n1184), .C1(new_n1175), .C2(new_n1180), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1174), .B1(new_n1185), .B2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1149), .A2(new_n1142), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n963), .B1(new_n1190), .B2(new_n928), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n1152), .B(new_n1187), .C1(new_n962), .C2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1189), .A2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT120), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1162), .A2(KEYINPUT119), .A3(new_n1152), .A4(new_n1156), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1150), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1194), .B1(new_n1197), .B2(new_n1171), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1173), .A2(new_n1193), .A3(new_n1198), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1197), .A2(new_n1171), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1200), .A2(new_n1192), .A3(new_n1189), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1199), .A2(new_n734), .A3(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n813), .A2(G125), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n836), .A2(G159), .ZN(new_n1204));
  XNOR2_X1  g1004(.A(KEYINPUT54), .B(G143), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n270), .B1(new_n823), .B2(new_n1205), .C1(new_n887), .C2(new_n830), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n820), .A2(new_n880), .ZN(new_n1207));
  AOI211_X1 g1007(.A(new_n1206), .B(new_n1207), .C1(G128), .C2(new_n817), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n827), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT53), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1210), .B1(new_n826), .B2(new_n882), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n1209), .A2(new_n1211), .B1(new_n833), .B2(G50), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1203), .A2(new_n1204), .A3(new_n1208), .A4(new_n1212), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(G97), .A2(new_n824), .B1(new_n844), .B2(G116), .ZN(new_n1214));
  OAI221_X1 g1014(.A(new_n1214), .B1(new_n504), .B2(new_n820), .C1(new_n872), .C2(new_n881), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(G77), .B2(new_n836), .ZN(new_n1216));
  AOI21_X1  g1016(.A(KEYINPUT122), .B1(new_n846), .B2(new_n316), .ZN(new_n1217));
  AND3_X1   g1017(.A1(new_n846), .A2(KEYINPUT122), .A3(new_n316), .ZN(new_n1218));
  AOI211_X1 g1018(.A(new_n1217), .B(new_n1218), .C1(G68), .C2(new_n833), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1216), .B(new_n1219), .C1(new_n664), .C2(new_n812), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n870), .B1(new_n1213), .B2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n868), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n786), .B1(new_n249), .B2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1224));
  AOI211_X1 g1024(.A(new_n1221), .B(new_n1223), .C1(new_n1224), .C2(new_n797), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1189), .A2(new_n785), .A3(new_n1192), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1226), .A2(KEYINPUT121), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT121), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1189), .A2(new_n1192), .A3(new_n1228), .A4(new_n785), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1225), .B1(new_n1227), .B2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1202), .A2(new_n1230), .ZN(G378));
  AND2_X1   g1031(.A1(new_n1189), .A2(new_n1192), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1171), .B1(new_n1232), .B2(new_n1200), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n976), .B1(new_n1175), .B2(new_n1180), .ZN(new_n1234));
  AND3_X1   g1034(.A1(new_n970), .A2(KEYINPUT103), .A3(new_n971), .ZN(new_n1235));
  AOI21_X1  g1035(.A(KEYINPUT103), .B1(new_n970), .B2(new_n971), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n1234), .B(G330), .C1(new_n1235), .C2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n264), .A2(new_n898), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n299), .A2(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n293), .A2(new_n298), .A3(new_n1238), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  XNOR2_X1  g1042(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1242), .A2(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1240), .A2(new_n1241), .A3(new_n1243), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1237), .A2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n974), .A2(new_n975), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1250), .A2(new_n1247), .A3(G330), .A4(new_n1234), .ZN(new_n1251));
  AND3_X1   g1051(.A1(new_n1249), .A2(new_n964), .A3(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n964), .B1(new_n1249), .B2(new_n1251), .ZN(new_n1253));
  OAI21_X1  g1053(.A(KEYINPUT57), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n734), .B1(new_n1233), .B2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1249), .A2(new_n1251), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n964), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1249), .A2(new_n964), .A3(new_n1251), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1172), .B1(new_n1193), .B2(new_n1197), .ZN(new_n1261));
  AOI21_X1  g1061(.A(KEYINPUT57), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  OR2_X1    g1062(.A1(new_n1255), .A2(new_n1262), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n785), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n786), .B1(G50), .B2(new_n1222), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n261), .B1(G33), .B2(G41), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1266), .B1(new_n316), .B2(new_n281), .ZN(new_n1267));
  AOI22_X1  g1067(.A1(new_n422), .A2(new_n824), .B1(new_n827), .B2(G77), .ZN(new_n1268));
  AOI211_X1 g1068(.A(G41), .B(new_n270), .C1(new_n844), .C2(G107), .ZN(new_n1269));
  AOI22_X1  g1069(.A1(new_n819), .A2(G97), .B1(new_n817), .B2(G116), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1059), .A2(new_n1268), .A3(new_n1269), .A4(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n833), .A2(G58), .ZN(new_n1272));
  XOR2_X1   g1072(.A(new_n1272), .B(KEYINPUT123), .Z(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  AOI211_X1 g1074(.A(new_n1271), .B(new_n1274), .C1(G283), .C2(new_n813), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1267), .B1(new_n1275), .B2(KEYINPUT58), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n809), .A2(G124), .ZN(new_n1277));
  AOI211_X1 g1077(.A(G33), .B(G41), .C1(new_n833), .C2(G159), .ZN(new_n1278));
  OR2_X1    g1078(.A1(new_n826), .A2(new_n1205), .ZN(new_n1279));
  AOI22_X1  g1079(.A1(new_n1279), .A2(KEYINPUT124), .B1(new_n819), .B2(G132), .ZN(new_n1280));
  AOI22_X1  g1080(.A1(G128), .A2(new_n844), .B1(new_n824), .B2(G137), .ZN(new_n1281));
  OAI211_X1 g1081(.A(new_n1280), .B(new_n1281), .C1(KEYINPUT124), .C2(new_n1279), .ZN(new_n1282));
  AOI22_X1  g1082(.A1(new_n836), .A2(G150), .B1(G125), .B2(new_n817), .ZN(new_n1283));
  OR2_X1    g1083(.A1(new_n1283), .A2(KEYINPUT125), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(KEYINPUT125), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1282), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT59), .ZN(new_n1287));
  OAI211_X1 g1087(.A(new_n1277), .B(new_n1278), .C1(new_n1286), .C2(new_n1287), .ZN(new_n1288));
  AND2_X1   g1088(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1289));
  OAI221_X1 g1089(.A(new_n1276), .B1(KEYINPUT58), .B2(new_n1275), .C1(new_n1288), .C2(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1265), .B1(new_n1290), .B2(new_n800), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1291), .B1(new_n1247), .B2(new_n798), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1264), .A2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1263), .A2(new_n1294), .ZN(G375));
  OAI21_X1  g1095(.A(new_n786), .B1(G68), .B2(new_n1222), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n813), .A2(G128), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n836), .A2(G50), .ZN(new_n1298));
  OAI22_X1  g1098(.A1(new_n887), .A2(new_n881), .B1(new_n820), .B2(new_n1205), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n270), .B1(new_n830), .B2(new_n880), .ZN(new_n1300));
  OAI22_X1  g1100(.A1(new_n823), .A2(new_n882), .B1(new_n826), .B2(new_n841), .ZN(new_n1301));
  NOR3_X1   g1101(.A1(new_n1299), .A2(new_n1300), .A3(new_n1301), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1297), .A2(new_n1273), .A3(new_n1298), .A4(new_n1302), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1082), .B1(new_n872), .B2(new_n830), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT126), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  OAI22_X1  g1106(.A1(new_n600), .A2(new_n820), .B1(new_n881), .B2(new_n664), .ZN(new_n1307));
  OAI221_X1 g1107(.A(new_n316), .B1(new_n826), .B2(new_n499), .C1(new_n504), .C2(new_n823), .ZN(new_n1308));
  NOR3_X1   g1108(.A1(new_n1307), .A2(new_n1053), .A3(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(G303), .ZN(new_n1310));
  OAI211_X1 g1110(.A(new_n1306), .B(new_n1309), .C1(new_n1310), .C2(new_n812), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1303), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1296), .B1(new_n1313), .B2(new_n800), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1314), .B1(new_n928), .B2(new_n798), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1315), .B1(new_n1197), .B2(new_n784), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(KEYINPUT127), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT127), .ZN(new_n1318));
  OAI211_X1 g1118(.A(new_n1318), .B(new_n1315), .C1(new_n1197), .C2(new_n784), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1317), .A2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1015), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1197), .A2(new_n1171), .ZN(new_n1322));
  NAND4_X1  g1122(.A1(new_n1173), .A2(new_n1198), .A3(new_n1321), .A4(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1320), .A2(new_n1323), .ZN(G381));
  INV_X1    g1124(.A(G384), .ZN(new_n1325));
  NAND4_X1  g1125(.A1(new_n1072), .A2(new_n854), .A3(new_n1325), .A4(new_n1105), .ZN(new_n1326));
  NOR4_X1   g1126(.A1(G387), .A2(G390), .A3(G381), .A4(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(G378), .ZN(new_n1328));
  NAND4_X1  g1128(.A1(new_n1327), .A2(new_n1328), .A3(new_n1263), .A4(new_n1294), .ZN(G407));
  NOR2_X1   g1129(.A1(new_n707), .A2(G343), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1328), .A2(new_n1330), .ZN(new_n1331));
  OAI211_X1 g1131(.A(G407), .B(G213), .C1(G375), .C2(new_n1331), .ZN(G409));
  XNOR2_X1  g1132(.A(G393), .B(G396), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1039), .A2(G390), .A3(new_n1068), .ZN(new_n1334));
  INV_X1    g1134(.A(new_n1334), .ZN(new_n1335));
  AOI21_X1  g1135(.A(G390), .B1(new_n1039), .B2(new_n1068), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1333), .B1(new_n1335), .B2(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(G390), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(G387), .A2(new_n1338), .ZN(new_n1339));
  XNOR2_X1  g1139(.A(G393), .B(new_n854), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1339), .A2(new_n1340), .A3(new_n1334), .ZN(new_n1341));
  AND2_X1   g1141(.A1(new_n1337), .A2(new_n1341), .ZN(new_n1342));
  INV_X1    g1142(.A(KEYINPUT63), .ZN(new_n1343));
  OAI211_X1 g1143(.A(G378), .B(new_n1294), .C1(new_n1255), .C2(new_n1262), .ZN(new_n1344));
  AND3_X1   g1144(.A1(new_n1260), .A2(new_n1261), .A3(new_n1321), .ZN(new_n1345));
  OAI211_X1 g1145(.A(new_n1202), .B(new_n1230), .C1(new_n1345), .C2(new_n1293), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1344), .A2(new_n1346), .ZN(new_n1347));
  INV_X1    g1147(.A(new_n1330), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1347), .A2(new_n1348), .ZN(new_n1349));
  OAI21_X1  g1149(.A(KEYINPUT60), .B1(new_n1197), .B2(new_n1171), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1350), .A2(new_n1322), .ZN(new_n1351));
  NAND3_X1  g1151(.A1(new_n1197), .A2(KEYINPUT60), .A3(new_n1171), .ZN(new_n1352));
  NAND3_X1  g1152(.A1(new_n1351), .A2(new_n734), .A3(new_n1352), .ZN(new_n1353));
  AND3_X1   g1153(.A1(new_n1353), .A2(G384), .A3(new_n1320), .ZN(new_n1354));
  AOI21_X1  g1154(.A(G384), .B1(new_n1353), .B2(new_n1320), .ZN(new_n1355));
  NOR2_X1   g1155(.A1(new_n1354), .A2(new_n1355), .ZN(new_n1356));
  INV_X1    g1156(.A(new_n1356), .ZN(new_n1357));
  OAI21_X1  g1157(.A(new_n1343), .B1(new_n1349), .B2(new_n1357), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1330), .A2(G2897), .ZN(new_n1359));
  INV_X1    g1159(.A(new_n1359), .ZN(new_n1360));
  OAI21_X1  g1160(.A(new_n1360), .B1(new_n1354), .B2(new_n1355), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1353), .A2(new_n1320), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1362), .A2(new_n1325), .ZN(new_n1363));
  NAND3_X1  g1163(.A1(new_n1353), .A2(G384), .A3(new_n1320), .ZN(new_n1364));
  NAND3_X1  g1164(.A1(new_n1363), .A2(new_n1364), .A3(new_n1359), .ZN(new_n1365));
  AND2_X1   g1165(.A1(new_n1361), .A2(new_n1365), .ZN(new_n1366));
  AOI21_X1  g1166(.A(KEYINPUT61), .B1(new_n1349), .B2(new_n1366), .ZN(new_n1367));
  AOI21_X1  g1167(.A(new_n1330), .B1(new_n1344), .B2(new_n1346), .ZN(new_n1368));
  NAND3_X1  g1168(.A1(new_n1368), .A2(KEYINPUT63), .A3(new_n1356), .ZN(new_n1369));
  NAND4_X1  g1169(.A1(new_n1342), .A2(new_n1358), .A3(new_n1367), .A4(new_n1369), .ZN(new_n1370));
  INV_X1    g1170(.A(KEYINPUT62), .ZN(new_n1371));
  AND3_X1   g1171(.A1(new_n1368), .A2(new_n1371), .A3(new_n1356), .ZN(new_n1372));
  INV_X1    g1172(.A(KEYINPUT61), .ZN(new_n1373));
  NAND2_X1  g1173(.A1(new_n1361), .A2(new_n1365), .ZN(new_n1374));
  OAI21_X1  g1174(.A(new_n1373), .B1(new_n1368), .B2(new_n1374), .ZN(new_n1375));
  AOI21_X1  g1175(.A(new_n1371), .B1(new_n1368), .B2(new_n1356), .ZN(new_n1376));
  NOR3_X1   g1176(.A1(new_n1372), .A2(new_n1375), .A3(new_n1376), .ZN(new_n1377));
  OAI21_X1  g1177(.A(new_n1370), .B1(new_n1377), .B2(new_n1342), .ZN(G405));
  NAND2_X1  g1178(.A1(new_n1337), .A2(new_n1341), .ZN(new_n1379));
  NAND2_X1  g1179(.A1(G375), .A2(new_n1328), .ZN(new_n1380));
  NAND3_X1  g1180(.A1(new_n1380), .A2(new_n1357), .A3(new_n1344), .ZN(new_n1381));
  INV_X1    g1181(.A(new_n1381), .ZN(new_n1382));
  AOI21_X1  g1182(.A(new_n1357), .B1(new_n1380), .B2(new_n1344), .ZN(new_n1383));
  OAI21_X1  g1183(.A(new_n1379), .B1(new_n1382), .B2(new_n1383), .ZN(new_n1384));
  INV_X1    g1184(.A(new_n1383), .ZN(new_n1385));
  NAND3_X1  g1185(.A1(new_n1385), .A2(new_n1342), .A3(new_n1381), .ZN(new_n1386));
  NAND2_X1  g1186(.A1(new_n1384), .A2(new_n1386), .ZN(G402));
endmodule


