//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 0 1 1 0 1 0 0 1 0 0 0 0 0 1 0 0 0 1 0 0 1 0 1 1 1 1 1 1 0 0 0 0 1 0 0 0 1 0 1 1 1 1 1 1 0 1 1 0 1 0 1 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n763, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n857, new_n859, new_n860, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n927, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n939, new_n940, new_n941,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n982, new_n983;
  INV_X1    g000(.A(KEYINPUT82), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT4), .ZN(new_n203));
  AND2_X1   g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(G155gat), .A2(G162gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G155gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT76), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT76), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G155gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n208), .A2(new_n210), .A3(G162gat), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n206), .B1(new_n211), .B2(KEYINPUT2), .ZN(new_n212));
  INV_X1    g011(.A(G148gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(G141gat), .ZN(new_n214));
  INV_X1    g013(.A(G141gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(G148gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT2), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n204), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n205), .B(KEYINPUT75), .ZN(new_n220));
  AOI22_X1  g019(.A1(new_n212), .A2(new_n217), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT70), .ZN(new_n222));
  INV_X1    g021(.A(G113gat), .ZN(new_n223));
  OR2_X1    g022(.A1(KEYINPUT69), .A2(G120gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(KEYINPUT69), .A2(G120gat), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n223), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(G120gat), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n227), .A2(G113gat), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n222), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT1), .ZN(new_n230));
  XNOR2_X1  g029(.A(G127gat), .B(G134gat), .ZN(new_n231));
  AND2_X1   g030(.A1(KEYINPUT69), .A2(G120gat), .ZN(new_n232));
  NOR2_X1   g031(.A1(KEYINPUT69), .A2(G120gat), .ZN(new_n233));
  OAI21_X1  g032(.A(G113gat), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n228), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n234), .A2(KEYINPUT70), .A3(new_n235), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n229), .A2(new_n230), .A3(new_n231), .A4(new_n236), .ZN(new_n237));
  XOR2_X1   g036(.A(G113gat), .B(G120gat), .Z(new_n238));
  AOI21_X1  g037(.A(new_n231), .B1(new_n238), .B2(new_n230), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n221), .A2(new_n237), .A3(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT79), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(KEYINPUT69), .B(G120gat), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n228), .B1(new_n244), .B2(G113gat), .ZN(new_n245));
  AOI21_X1  g044(.A(KEYINPUT1), .B1(new_n245), .B2(KEYINPUT70), .ZN(new_n246));
  INV_X1    g045(.A(new_n231), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n234), .A2(new_n235), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n247), .B1(new_n248), .B2(new_n222), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n239), .B1(new_n246), .B2(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n250), .A2(KEYINPUT79), .A3(new_n221), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n203), .B1(new_n243), .B2(new_n251), .ZN(new_n252));
  XOR2_X1   g051(.A(KEYINPUT78), .B(KEYINPUT4), .Z(new_n253));
  NOR2_X1   g052(.A1(new_n241), .A2(new_n253), .ZN(new_n254));
  OAI21_X1  g053(.A(KEYINPUT81), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  AOI21_X1  g054(.A(KEYINPUT79), .B1(new_n250), .B2(new_n221), .ZN(new_n256));
  AND4_X1   g055(.A1(KEYINPUT79), .A2(new_n221), .A3(new_n237), .A4(new_n240), .ZN(new_n257));
  OAI21_X1  g056(.A(KEYINPUT4), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT81), .ZN(new_n259));
  INV_X1    g058(.A(new_n254), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n258), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(G225gat), .A2(G233gat), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n263), .A2(KEYINPUT5), .ZN(new_n264));
  AND2_X1   g063(.A1(new_n219), .A2(new_n220), .ZN(new_n265));
  XNOR2_X1  g064(.A(G141gat), .B(G148gat), .ZN(new_n266));
  AOI211_X1 g065(.A(new_n266), .B(new_n206), .C1(KEYINPUT2), .C2(new_n211), .ZN(new_n267));
  OAI21_X1  g066(.A(KEYINPUT3), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT3), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n221), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n237), .A2(new_n240), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n268), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT77), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n268), .A2(new_n270), .A3(new_n271), .A4(KEYINPUT77), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n255), .A2(new_n261), .A3(new_n264), .A4(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n243), .A2(new_n203), .A3(new_n251), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n241), .A2(new_n262), .A3(new_n253), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(new_n276), .ZN(new_n281));
  OAI22_X1  g080(.A1(new_n256), .A2(new_n257), .B1(new_n221), .B2(new_n250), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(new_n263), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n281), .A2(KEYINPUT5), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n277), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(G57gat), .B(G85gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(G1gat), .B(G29gat), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n286), .B(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n289));
  XOR2_X1   g088(.A(new_n288), .B(new_n289), .Z(new_n290));
  NAND2_X1  g089(.A1(new_n285), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT6), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n202), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n290), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n277), .A2(new_n284), .A3(new_n294), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n291), .A2(new_n292), .A3(new_n295), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n294), .B1(new_n277), .B2(new_n284), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n297), .A2(KEYINPUT82), .A3(KEYINPUT6), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n293), .A2(new_n296), .A3(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(G197gat), .B(G204gat), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT22), .ZN(new_n301));
  INV_X1    g100(.A(G211gat), .ZN(new_n302));
  INV_X1    g101(.A(G218gat), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n300), .A2(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(G211gat), .B(G218gat), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n305), .B(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT26), .ZN(new_n308));
  INV_X1    g107(.A(G169gat), .ZN(new_n309));
  INV_X1    g108(.A(G176gat), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(G169gat), .A2(G176gat), .ZN(new_n312));
  OAI21_X1  g111(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n311), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(G183gat), .A2(G190gat), .ZN(new_n315));
  OR2_X1    g114(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n317));
  AOI21_X1  g116(.A(G190gat), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT28), .ZN(new_n319));
  OAI211_X1 g118(.A(new_n314), .B(new_n315), .C1(new_n318), .C2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n318), .A2(new_n319), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT67), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT23), .ZN(new_n324));
  NOR3_X1   g123(.A1(new_n324), .A2(G169gat), .A3(G176gat), .ZN(new_n325));
  INV_X1    g124(.A(new_n312), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n323), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT66), .ZN(new_n328));
  NOR2_X1   g127(.A1(G169gat), .A2(G176gat), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n328), .B1(new_n329), .B2(KEYINPUT23), .ZN(new_n330));
  OAI211_X1 g129(.A(new_n324), .B(KEYINPUT66), .C1(G169gat), .C2(G176gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT24), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n315), .A2(new_n333), .ZN(new_n334));
  OAI22_X1  g133(.A1(new_n334), .A2(KEYINPUT68), .B1(G183gat), .B2(G190gat), .ZN(new_n335));
  NAND3_X1  g134(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n336));
  AOI21_X1  g135(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT68), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n336), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  OAI211_X1 g138(.A(new_n327), .B(new_n332), .C1(new_n335), .C2(new_n339), .ZN(new_n340));
  AOI22_X1  g139(.A1(new_n321), .A2(new_n322), .B1(new_n340), .B2(KEYINPUT25), .ZN(new_n341));
  INV_X1    g140(.A(G183gat), .ZN(new_n342));
  INV_X1    g141(.A(G190gat), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n342), .A2(new_n343), .A3(KEYINPUT65), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT65), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n345), .B1(G183gat), .B2(G190gat), .ZN(new_n346));
  NAND4_X1  g145(.A1(new_n344), .A2(new_n334), .A3(new_n346), .A4(new_n336), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT25), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n332), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(KEYINPUT67), .A2(KEYINPUT25), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n325), .A2(new_n326), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n341), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT29), .ZN(new_n355));
  AOI22_X1  g154(.A1(new_n354), .A2(new_n355), .B1(G226gat), .B2(G233gat), .ZN(new_n356));
  INV_X1    g155(.A(G226gat), .ZN(new_n357));
  INV_X1    g156(.A(G233gat), .ZN(new_n358));
  AOI211_X1 g157(.A(new_n357), .B(new_n358), .C1(new_n341), .C2(new_n353), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n307), .B1(new_n356), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n340), .A2(KEYINPUT25), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n316), .A2(new_n317), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(new_n343), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT28), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n364), .A2(new_n315), .A3(new_n322), .A4(new_n314), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n361), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n352), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n367), .B1(new_n349), .B2(new_n350), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  OAI22_X1  g168(.A1(new_n369), .A2(KEYINPUT29), .B1(new_n357), .B2(new_n358), .ZN(new_n370));
  INV_X1    g169(.A(new_n307), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n354), .A2(G226gat), .A3(G233gat), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n360), .A2(new_n373), .ZN(new_n374));
  XOR2_X1   g173(.A(G8gat), .B(G36gat), .Z(new_n375));
  XNOR2_X1  g174(.A(new_n375), .B(G64gat), .ZN(new_n376));
  INV_X1    g175(.A(G92gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n376), .B(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n374), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n378), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n360), .A2(new_n373), .A3(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n379), .A2(KEYINPUT30), .A3(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT30), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n360), .A2(new_n373), .A3(new_n383), .A4(new_n380), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n299), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n307), .A2(KEYINPUT29), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT84), .ZN(new_n389));
  AOI21_X1  g188(.A(KEYINPUT3), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g189(.A(KEYINPUT84), .B1(new_n307), .B2(KEYINPUT29), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n221), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n371), .B1(new_n270), .B2(new_n355), .ZN(new_n393));
  INV_X1    g192(.A(G228gat), .ZN(new_n394));
  OAI22_X1  g193(.A1(new_n392), .A2(new_n393), .B1(new_n394), .B2(new_n358), .ZN(new_n395));
  INV_X1    g194(.A(new_n221), .ZN(new_n396));
  AOI211_X1 g195(.A(new_n394), .B(new_n358), .C1(new_n388), .C2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n393), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n397), .A2(new_n268), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n395), .A2(new_n399), .ZN(new_n400));
  XOR2_X1   g199(.A(KEYINPUT85), .B(G22gat), .Z(new_n401));
  NOR2_X1   g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(KEYINPUT86), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT86), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n404), .B1(new_n400), .B2(new_n401), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n400), .A2(G22gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(G78gat), .B(G106gat), .ZN(new_n407));
  INV_X1    g206(.A(G50gat), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n407), .B(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n409), .B(KEYINPUT83), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n410), .B(KEYINPUT31), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n403), .A2(new_n405), .A3(new_n406), .A4(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n411), .ZN(new_n413));
  AND2_X1   g212(.A1(new_n400), .A2(new_n401), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n413), .B1(new_n414), .B2(new_n402), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n250), .B1(new_n366), .B2(new_n368), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n341), .A2(new_n271), .A3(new_n353), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT34), .ZN(new_n420));
  NAND2_X1  g219(.A1(G227gat), .A2(G233gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n421), .B(KEYINPUT64), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n419), .A2(new_n420), .A3(new_n422), .ZN(new_n423));
  NOR3_X1   g222(.A1(new_n366), .A2(new_n250), .A3(new_n368), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n271), .B1(new_n341), .B2(new_n353), .ZN(new_n425));
  OAI21_X1  g224(.A(KEYINPUT72), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT72), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n417), .A2(new_n418), .A3(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n426), .A2(new_n421), .A3(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT73), .ZN(new_n430));
  XOR2_X1   g229(.A(KEYINPUT71), .B(KEYINPUT34), .Z(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  AND3_X1   g231(.A1(new_n429), .A2(new_n430), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n430), .B1(new_n429), .B2(new_n432), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n423), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  OR2_X1    g234(.A1(new_n419), .A2(new_n422), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(KEYINPUT32), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n435), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT33), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n436), .A2(new_n440), .ZN(new_n441));
  XNOR2_X1  g240(.A(G15gat), .B(G43gat), .ZN(new_n442));
  INV_X1    g241(.A(G71gat), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n442), .B(new_n443), .ZN(new_n444));
  XNOR2_X1  g243(.A(new_n444), .B(G99gat), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n441), .A2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  OAI211_X1 g246(.A(new_n437), .B(new_n423), .C1(new_n433), .C2(new_n434), .ZN(new_n448));
  AND3_X1   g247(.A1(new_n439), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n447), .B1(new_n439), .B2(new_n448), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT89), .ZN(new_n451));
  NOR3_X1   g250(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n429), .A2(new_n432), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT73), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n429), .A2(new_n430), .A3(new_n432), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n437), .B1(new_n456), .B2(new_n423), .ZN(new_n457));
  INV_X1    g256(.A(new_n448), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n446), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n439), .A2(new_n447), .A3(new_n448), .ZN(new_n460));
  AOI21_X1  g259(.A(KEYINPUT89), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n387), .B(new_n416), .C1(new_n452), .C2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT35), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n416), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n386), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT40), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT39), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n282), .A2(new_n263), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n255), .A2(new_n261), .A3(new_n276), .ZN(new_n470));
  AOI211_X1 g269(.A(new_n468), .B(new_n469), .C1(new_n470), .C2(new_n263), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n470), .A2(new_n468), .A3(new_n263), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(new_n294), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n467), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n469), .B1(new_n470), .B2(new_n263), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(KEYINPUT39), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n476), .A2(KEYINPUT40), .A3(new_n294), .A4(new_n472), .ZN(new_n477));
  INV_X1    g276(.A(new_n385), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n474), .A2(new_n477), .A3(new_n291), .A4(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT37), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n480), .B1(new_n360), .B2(new_n373), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  OR2_X1    g281(.A1(new_n482), .A2(KEYINPUT87), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n380), .B1(new_n482), .B2(KEYINPUT87), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT38), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n360), .A2(new_n373), .A3(new_n480), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n483), .A2(new_n484), .A3(new_n485), .A4(new_n486), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n487), .A2(new_n293), .A3(new_n298), .A4(new_n296), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT88), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n489), .B1(new_n481), .B2(new_n380), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(new_n486), .ZN(new_n491));
  NOR3_X1   g290(.A1(new_n481), .A2(new_n489), .A3(new_n380), .ZN(new_n492));
  OAI21_X1  g291(.A(KEYINPUT38), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(new_n381), .ZN(new_n494));
  OAI211_X1 g293(.A(new_n479), .B(new_n416), .C1(new_n488), .C2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT36), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n459), .A2(new_n460), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT74), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  AOI211_X1 g298(.A(KEYINPUT74), .B(KEYINPUT36), .C1(new_n459), .C2(new_n460), .ZN(new_n500));
  OAI211_X1 g299(.A(new_n466), .B(new_n495), .C1(new_n499), .C2(new_n500), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n497), .A2(new_n465), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n502), .A2(KEYINPUT35), .A3(new_n387), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n464), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(G8gat), .ZN(new_n505));
  XNOR2_X1  g304(.A(G15gat), .B(G22gat), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT16), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n506), .B1(new_n507), .B2(G1gat), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT94), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n505), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n508), .B1(G1gat), .B2(new_n506), .ZN(new_n511));
  XOR2_X1   g310(.A(new_n510), .B(new_n511), .Z(new_n512));
  INV_X1    g311(.A(KEYINPUT15), .ZN(new_n513));
  OR2_X1    g312(.A1(G43gat), .A2(G50gat), .ZN(new_n514));
  NAND2_X1  g313(.A1(G43gat), .A2(G50gat), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  XOR2_X1   g315(.A(KEYINPUT92), .B(G43gat), .Z(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(new_n408), .ZN(new_n518));
  AOI21_X1  g317(.A(KEYINPUT15), .B1(G43gat), .B2(G50gat), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n516), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(G29gat), .ZN(new_n521));
  INV_X1    g320(.A(G36gat), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n521), .A2(new_n522), .A3(KEYINPUT90), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT90), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n524), .B1(G29gat), .B2(G36gat), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n523), .A2(new_n525), .A3(KEYINPUT14), .ZN(new_n526));
  XOR2_X1   g325(.A(KEYINPUT91), .B(G36gat), .Z(new_n527));
  OAI221_X1 g326(.A(new_n526), .B1(KEYINPUT14), .B2(new_n525), .C1(new_n527), .C2(new_n521), .ZN(new_n528));
  OR2_X1    g327(.A1(new_n520), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(new_n516), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n512), .A2(new_n532), .ZN(new_n533));
  AND2_X1   g332(.A1(new_n529), .A2(new_n531), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n534), .A2(KEYINPUT93), .A3(KEYINPUT17), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT17), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT93), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n536), .B1(new_n532), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n535), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n533), .B1(new_n539), .B2(new_n512), .ZN(new_n540));
  NAND2_X1  g339(.A1(G229gat), .A2(G233gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n542), .B(KEYINPUT18), .ZN(new_n543));
  XNOR2_X1  g342(.A(G113gat), .B(G141gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n544), .B(G197gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n545), .B(KEYINPUT11), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n546), .B(new_n309), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(KEYINPUT12), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n534), .B(new_n512), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n541), .B(KEYINPUT13), .ZN(new_n550));
  OR2_X1    g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AND3_X1   g350(.A1(new_n543), .A2(new_n548), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n548), .B1(new_n543), .B2(new_n551), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n504), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT95), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n556), .B(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n512), .ZN(new_n559));
  XNOR2_X1  g358(.A(G57gat), .B(G64gat), .ZN(new_n560));
  AOI21_X1  g359(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n560), .B1(KEYINPUT96), .B2(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(G71gat), .B(G78gat), .ZN(new_n563));
  OAI211_X1 g362(.A(new_n562), .B(new_n563), .C1(KEYINPUT96), .C2(new_n561), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT9), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n560), .A2(new_n565), .ZN(new_n566));
  OR2_X1    g365(.A1(new_n566), .A2(new_n563), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(KEYINPUT97), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n559), .B1(new_n569), .B2(KEYINPUT21), .ZN(new_n570));
  AOI21_X1  g369(.A(KEYINPUT21), .B1(new_n564), .B2(new_n567), .ZN(new_n571));
  INV_X1    g370(.A(G127gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n570), .B(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n575));
  XNOR2_X1  g374(.A(G155gat), .B(G183gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n574), .B(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(G231gat), .A2(G233gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(new_n302), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n578), .B(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(G85gat), .A2(G92gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(KEYINPUT7), .ZN(new_n583));
  NAND2_X1  g382(.A1(G99gat), .A2(G106gat), .ZN(new_n584));
  INV_X1    g383(.A(G85gat), .ZN(new_n585));
  AOI22_X1  g384(.A1(KEYINPUT8), .A2(new_n584), .B1(new_n585), .B2(new_n377), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G99gat), .B(G106gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n589), .B1(new_n535), .B2(new_n538), .ZN(new_n590));
  INV_X1    g389(.A(G232gat), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n591), .A2(new_n358), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT41), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n590), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n589), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n532), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n343), .B1(new_n596), .B2(new_n599), .ZN(new_n600));
  NOR4_X1   g399(.A1(new_n590), .A2(G190gat), .A3(new_n598), .A4(new_n595), .ZN(new_n601));
  NOR3_X1   g400(.A1(new_n600), .A2(new_n601), .A3(new_n303), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n539), .A2(new_n597), .ZN(new_n603));
  INV_X1    g402(.A(new_n595), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n603), .A2(new_n599), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(G190gat), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n596), .A2(new_n343), .A3(new_n599), .ZN(new_n607));
  AOI21_X1  g406(.A(G218gat), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  OAI21_X1  g407(.A(KEYINPUT98), .B1(new_n602), .B2(new_n608), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n303), .B1(new_n600), .B2(new_n601), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n606), .A2(G218gat), .A3(new_n607), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT98), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n592), .A2(KEYINPUT41), .ZN(new_n614));
  XNOR2_X1  g413(.A(G134gat), .B(G162gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n609), .A2(new_n613), .A3(new_n617), .ZN(new_n618));
  OR2_X1    g417(.A1(new_n613), .A2(new_n617), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n581), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT100), .ZN(new_n621));
  NAND2_X1  g420(.A1(G230gat), .A2(G233gat), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n569), .A2(KEYINPUT10), .A3(new_n589), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n589), .B(new_n568), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT10), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n623), .B1(new_n624), .B2(new_n627), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n625), .A2(new_n622), .ZN(new_n629));
  XNOR2_X1  g428(.A(G120gat), .B(G148gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(new_n310), .ZN(new_n631));
  INV_X1    g430(.A(G204gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NOR3_X1   g432(.A1(new_n628), .A2(new_n629), .A3(new_n633), .ZN(new_n634));
  OR2_X1    g433(.A1(new_n634), .A2(KEYINPUT99), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(KEYINPUT99), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n633), .B1(new_n628), .B2(new_n629), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  AND3_X1   g439(.A1(new_n620), .A2(new_n621), .A3(new_n640), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n621), .B1(new_n620), .B2(new_n640), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  AND2_X1   g443(.A1(new_n558), .A2(new_n644), .ZN(new_n645));
  AND3_X1   g444(.A1(new_n293), .A2(new_n296), .A3(new_n298), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(G1gat), .ZN(G1324gat));
  NAND3_X1  g447(.A1(new_n558), .A2(new_n478), .A3(new_n644), .ZN(new_n649));
  NOR2_X1   g448(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n507), .A2(new_n505), .ZN(new_n651));
  NOR3_X1   g450(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  AND2_X1   g451(.A1(new_n649), .A2(G8gat), .ZN(new_n653));
  OAI21_X1  g452(.A(KEYINPUT42), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n654), .B1(KEYINPUT42), .B2(new_n652), .ZN(G1325gat));
  OR2_X1    g454(.A1(new_n452), .A2(new_n461), .ZN(new_n656));
  AOI21_X1  g455(.A(G15gat), .B1(new_n645), .B2(new_n656), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n499), .A2(new_n500), .ZN(new_n658));
  AND2_X1   g457(.A1(new_n658), .A2(G15gat), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n657), .B1(new_n645), .B2(new_n659), .ZN(G1326gat));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n465), .ZN(new_n661));
  XNOR2_X1  g460(.A(KEYINPUT43), .B(G22gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(G1327gat));
  NAND2_X1  g462(.A1(new_n618), .A2(new_n619), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n581), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n666), .A2(new_n639), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g467(.A(new_n668), .B(KEYINPUT101), .Z(new_n669));
  NAND3_X1  g468(.A1(new_n558), .A2(new_n646), .A3(new_n669), .ZN(new_n670));
  OR3_X1    g469(.A1(new_n670), .A2(KEYINPUT45), .A3(G29gat), .ZN(new_n671));
  OAI21_X1  g470(.A(KEYINPUT45), .B1(new_n670), .B2(G29gat), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AND2_X1   g472(.A1(new_n504), .A2(new_n665), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT44), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n464), .A2(new_n503), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT103), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n495), .B1(new_n499), .B2(new_n500), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n466), .A2(KEYINPUT102), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT102), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n386), .A2(new_n680), .A3(new_n465), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n677), .B1(new_n678), .B2(new_n682), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n498), .B1(new_n449), .B2(new_n450), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(KEYINPUT36), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n497), .A2(new_n498), .A3(new_n496), .ZN(new_n686));
  AND2_X1   g485(.A1(new_n479), .A2(new_n416), .ZN(new_n687));
  NAND4_X1  g486(.A1(new_n646), .A2(new_n381), .A3(new_n493), .A4(new_n487), .ZN(new_n688));
  AOI22_X1  g487(.A1(new_n685), .A2(new_n686), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  AOI211_X1 g488(.A(KEYINPUT102), .B(new_n416), .C1(new_n299), .C2(new_n385), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n680), .B1(new_n386), .B2(new_n465), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n689), .A2(KEYINPUT103), .A3(new_n692), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n676), .B1(new_n683), .B2(new_n693), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n618), .A2(new_n619), .A3(KEYINPUT104), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  AOI21_X1  g495(.A(KEYINPUT104), .B1(new_n618), .B2(new_n619), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n699), .A2(KEYINPUT44), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  OAI22_X1  g500(.A1(new_n674), .A2(new_n675), .B1(new_n694), .B2(new_n701), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n702), .A2(new_n555), .A3(new_n667), .ZN(new_n703));
  OAI21_X1  g502(.A(G29gat), .B1(new_n703), .B2(new_n299), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n673), .A2(new_n704), .ZN(G1328gat));
  NAND3_X1  g504(.A1(new_n558), .A2(new_n478), .A3(new_n669), .ZN(new_n706));
  INV_X1    g505(.A(new_n527), .ZN(new_n707));
  OR3_X1    g506(.A1(new_n706), .A2(KEYINPUT46), .A3(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n707), .B1(new_n703), .B2(new_n385), .ZN(new_n709));
  OAI21_X1  g508(.A(KEYINPUT46), .B1(new_n706), .B2(new_n707), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n708), .A2(new_n709), .A3(new_n710), .ZN(G1329gat));
  AOI21_X1  g510(.A(new_n675), .B1(new_n504), .B2(new_n665), .ZN(new_n712));
  AND2_X1   g511(.A1(new_n464), .A2(new_n503), .ZN(new_n713));
  NOR3_X1   g512(.A1(new_n678), .A2(new_n682), .A3(new_n677), .ZN(new_n714));
  AOI21_X1  g513(.A(KEYINPUT103), .B1(new_n689), .B2(new_n692), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n713), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n712), .B1(new_n716), .B2(new_n700), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n717), .A2(new_n554), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT106), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n718), .A2(new_n719), .A3(new_n658), .A4(new_n667), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n702), .A2(new_n555), .A3(new_n658), .A4(new_n667), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(KEYINPUT106), .ZN(new_n722));
  INV_X1    g521(.A(new_n517), .ZN(new_n723));
  AND3_X1   g522(.A1(new_n720), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n558), .A2(new_n517), .A3(new_n656), .A4(new_n669), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(KEYINPUT47), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n721), .A2(new_n723), .ZN(new_n727));
  AND2_X1   g526(.A1(new_n727), .A2(new_n725), .ZN(new_n728));
  XNOR2_X1  g527(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n729));
  OAI22_X1  g528(.A1(new_n724), .A2(new_n726), .B1(new_n728), .B2(new_n729), .ZN(G1330gat));
  OAI21_X1  g529(.A(G50gat), .B1(new_n703), .B2(new_n416), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n558), .A2(new_n669), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n465), .A2(new_n408), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(KEYINPUT107), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n731), .B1(new_n732), .B2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT48), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  OAI211_X1 g536(.A(new_n731), .B(KEYINPUT48), .C1(new_n732), .C2(new_n734), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(G1331gat));
  NOR2_X1   g538(.A1(new_n694), .A2(new_n555), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n646), .B(KEYINPUT108), .ZN(new_n741));
  INV_X1    g540(.A(new_n620), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n742), .A2(new_n640), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n740), .A2(new_n741), .A3(new_n743), .ZN(new_n744));
  XNOR2_X1  g543(.A(KEYINPUT109), .B(G57gat), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n744), .B(new_n745), .ZN(G1332gat));
  AOI21_X1  g545(.A(KEYINPUT110), .B1(new_n740), .B2(new_n743), .ZN(new_n747));
  AND4_X1   g546(.A1(KEYINPUT110), .A2(new_n716), .A3(new_n554), .A4(new_n743), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n749), .A2(new_n385), .ZN(new_n750));
  NOR2_X1   g549(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n751));
  AND2_X1   g550(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n750), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n753), .B1(new_n750), .B2(new_n751), .ZN(G1333gat));
  XNOR2_X1  g553(.A(new_n656), .B(KEYINPUT111), .ZN(new_n755));
  AND4_X1   g554(.A1(new_n443), .A2(new_n740), .A3(new_n743), .A4(new_n755), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n658), .B1(new_n747), .B2(new_n748), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n756), .B1(new_n757), .B2(G71gat), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT50), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  AOI211_X1 g559(.A(KEYINPUT50), .B(new_n756), .C1(new_n757), .C2(G71gat), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n760), .A2(new_n761), .ZN(G1334gat));
  OAI21_X1  g561(.A(new_n465), .B1(new_n747), .B2(new_n748), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(G78gat), .ZN(G1335gat));
  INV_X1    g563(.A(KEYINPUT112), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n555), .A2(new_n666), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n767), .A2(new_n640), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n765), .B1(new_n717), .B2(new_n769), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n694), .A2(new_n701), .ZN(new_n771));
  OAI211_X1 g570(.A(KEYINPUT112), .B(new_n768), .C1(new_n771), .C2(new_n712), .ZN(new_n772));
  AND2_X1   g571(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n773), .A2(new_n585), .A3(new_n299), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n683), .A2(new_n693), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n767), .B1(new_n775), .B2(new_n713), .ZN(new_n776));
  AOI21_X1  g575(.A(KEYINPUT51), .B1(new_n776), .B2(new_n665), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT51), .ZN(new_n778));
  NOR4_X1   g577(.A1(new_n694), .A2(new_n778), .A3(new_n664), .A4(new_n767), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n780), .A2(new_n640), .ZN(new_n781));
  AOI21_X1  g580(.A(G85gat), .B1(new_n781), .B2(new_n646), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n774), .A2(new_n782), .ZN(G1336gat));
  OAI211_X1 g582(.A(KEYINPUT52), .B(G92gat), .C1(new_n773), .C2(new_n385), .ZN(new_n784));
  NOR2_X1   g583(.A1(KEYINPUT113), .A2(KEYINPUT52), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n385), .A2(G92gat), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n785), .B1(new_n781), .B2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT52), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n702), .A2(new_n768), .ZN(new_n789));
  OAI21_X1  g588(.A(G92gat), .B1(new_n789), .B2(new_n385), .ZN(new_n790));
  OAI211_X1 g589(.A(new_n639), .B(new_n786), .C1(new_n777), .C2(new_n779), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n790), .B1(new_n791), .B2(KEYINPUT113), .ZN(new_n792));
  AOI22_X1  g591(.A1(new_n784), .A2(new_n787), .B1(new_n788), .B2(new_n792), .ZN(G1337gat));
  AOI21_X1  g592(.A(G99gat), .B1(new_n781), .B2(new_n656), .ZN(new_n794));
  INV_X1    g593(.A(new_n658), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n773), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n794), .B1(new_n796), .B2(G99gat), .ZN(G1338gat));
  XNOR2_X1  g596(.A(KEYINPUT114), .B(G106gat), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n770), .A2(new_n772), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n799), .B1(new_n800), .B2(new_n465), .ZN(new_n801));
  OAI211_X1 g600(.A(new_n465), .B(new_n639), .C1(new_n777), .C2(new_n779), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n802), .A2(G106gat), .ZN(new_n803));
  OAI21_X1  g602(.A(KEYINPUT53), .B1(new_n801), .B2(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n798), .B1(new_n789), .B2(new_n416), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT53), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n805), .B(new_n806), .C1(new_n802), .C2(G106gat), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n804), .A2(new_n807), .ZN(G1339gat));
  NAND3_X1  g607(.A1(new_n543), .A2(new_n548), .A3(new_n551), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n549), .A2(new_n550), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n810), .B1(new_n540), .B2(new_n541), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(new_n547), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n639), .A2(new_n809), .A3(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(new_n633), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT115), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n628), .B1(new_n815), .B2(KEYINPUT54), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n624), .A2(new_n627), .A3(new_n623), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(KEYINPUT54), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  OAI211_X1 g618(.A(KEYINPUT54), .B(new_n817), .C1(new_n628), .C2(new_n815), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n814), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  AOI22_X1  g620(.A1(new_n821), .A2(KEYINPUT55), .B1(new_n635), .B2(new_n636), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n819), .A2(new_n820), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(new_n633), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT55), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n822), .A2(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n813), .B1(new_n554), .B2(new_n827), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n828), .B1(new_n696), .B2(new_n697), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT104), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n664), .A2(new_n830), .ZN(new_n831));
  AND4_X1   g630(.A1(new_n809), .A2(new_n822), .A3(new_n826), .A4(new_n812), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n831), .A2(new_n695), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n666), .B1(new_n829), .B2(new_n833), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n742), .A2(new_n555), .A3(new_n639), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n837), .A2(new_n741), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n838), .A2(KEYINPUT116), .A3(new_n385), .A4(new_n502), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT116), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n837), .A2(new_n385), .A3(new_n741), .ZN(new_n841));
  INV_X1    g640(.A(new_n502), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n840), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n554), .A2(G113gat), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n839), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n836), .A2(new_n465), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n299), .A2(new_n478), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n846), .A2(new_n656), .A3(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(G113gat), .B1(new_n848), .B2(new_n554), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n845), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(KEYINPUT117), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT117), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n845), .A2(new_n852), .A3(new_n849), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n851), .A2(new_n853), .ZN(G1340gat));
  OAI21_X1  g653(.A(G120gat), .B1(new_n848), .B2(new_n640), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n843), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n639), .A2(new_n244), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n855), .B1(new_n856), .B2(new_n857), .ZN(G1341gat));
  NOR3_X1   g657(.A1(new_n848), .A2(new_n572), .A3(new_n581), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n838), .A2(new_n385), .A3(new_n502), .A4(new_n666), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n859), .B1(new_n572), .B2(new_n860), .ZN(G1342gat));
  NOR4_X1   g660(.A1(new_n841), .A2(G134gat), .A3(new_n842), .A4(new_n664), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT56), .ZN(new_n863));
  OR2_X1    g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  OAI21_X1  g663(.A(G134gat), .B1(new_n848), .B2(new_n664), .ZN(new_n865));
  AND3_X1   g664(.A1(new_n862), .A2(KEYINPUT118), .A3(new_n863), .ZN(new_n866));
  AOI21_X1  g665(.A(KEYINPUT118), .B1(new_n862), .B2(new_n863), .ZN(new_n867));
  OAI211_X1 g666(.A(new_n864), .B(new_n865), .C1(new_n866), .C2(new_n867), .ZN(G1343gat));
  NOR2_X1   g667(.A1(new_n658), .A2(new_n416), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  NOR4_X1   g669(.A1(new_n841), .A2(G141gat), .A3(new_n554), .A4(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  AND2_X1   g671(.A1(new_n821), .A2(KEYINPUT119), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n825), .B1(new_n821), .B2(KEYINPUT119), .ZN(new_n874));
  OAI22_X1  g673(.A1(new_n873), .A2(new_n874), .B1(new_n552), .B2(new_n553), .ZN(new_n875));
  INV_X1    g674(.A(new_n822), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n813), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(new_n664), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n666), .B1(new_n878), .B2(new_n833), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n465), .B1(new_n879), .B2(new_n835), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(KEYINPUT57), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n795), .A2(new_n847), .ZN(new_n882));
  INV_X1    g681(.A(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT57), .ZN(new_n884));
  OAI211_X1 g683(.A(new_n884), .B(new_n465), .C1(new_n834), .C2(new_n835), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n881), .A2(new_n883), .A3(new_n885), .ZN(new_n886));
  OAI21_X1  g685(.A(G141gat), .B1(new_n886), .B2(new_n554), .ZN(new_n887));
  XOR2_X1   g686(.A(KEYINPUT121), .B(KEYINPUT58), .Z(new_n888));
  NAND3_X1  g687(.A1(new_n872), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n882), .B1(new_n880), .B2(KEYINPUT57), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT120), .ZN(new_n891));
  AND3_X1   g690(.A1(new_n890), .A2(new_n891), .A3(new_n885), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n891), .B1(new_n890), .B2(new_n885), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n555), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n871), .B1(new_n894), .B2(G141gat), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT58), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n889), .B1(new_n895), .B2(new_n896), .ZN(G1344gat));
  NOR2_X1   g696(.A1(new_n841), .A2(new_n870), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n898), .A2(new_n213), .A3(new_n639), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n886), .A2(KEYINPUT120), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n890), .A2(new_n891), .A3(new_n885), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n640), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n902), .A2(KEYINPUT59), .A3(new_n213), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT59), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n554), .B1(new_n641), .B2(new_n642), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(KEYINPUT122), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n877), .A2(new_n664), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n665), .A2(new_n832), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n581), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT122), .ZN(new_n910));
  OAI211_X1 g709(.A(new_n910), .B(new_n554), .C1(new_n641), .C2(new_n642), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n906), .A2(new_n909), .A3(new_n911), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n912), .A2(new_n884), .A3(new_n465), .ZN(new_n913));
  OAI21_X1  g712(.A(KEYINPUT57), .B1(new_n836), .B2(new_n416), .ZN(new_n914));
  AND3_X1   g713(.A1(new_n913), .A2(new_n639), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(new_n883), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n904), .B1(new_n916), .B2(G148gat), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n899), .B1(new_n903), .B2(new_n917), .ZN(G1345gat));
  NOR2_X1   g717(.A1(new_n892), .A2(new_n893), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n208), .A2(new_n210), .ZN(new_n920));
  NOR3_X1   g719(.A1(new_n919), .A2(new_n920), .A3(new_n581), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n898), .A2(new_n666), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n921), .B1(new_n920), .B2(new_n922), .ZN(G1346gat));
  INV_X1    g722(.A(G162gat), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n898), .A2(new_n924), .A3(new_n665), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(KEYINPUT123), .ZN(new_n926));
  OAI21_X1  g725(.A(G162gat), .B1(new_n919), .B2(new_n699), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(G1347gat));
  NOR2_X1   g727(.A1(new_n741), .A2(new_n385), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n846), .A2(new_n755), .A3(new_n929), .ZN(new_n930));
  OAI21_X1  g729(.A(G169gat), .B1(new_n930), .B2(new_n554), .ZN(new_n931));
  NOR4_X1   g730(.A1(new_n836), .A2(new_n646), .A3(new_n385), .A4(new_n842), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n932), .A2(new_n309), .A3(new_n555), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n931), .A2(new_n933), .ZN(G1348gat));
  AOI21_X1  g733(.A(G176gat), .B1(new_n932), .B2(new_n639), .ZN(new_n935));
  INV_X1    g734(.A(new_n930), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n640), .A2(new_n310), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n935), .B1(new_n936), .B2(new_n937), .ZN(G1349gat));
  OAI21_X1  g737(.A(G183gat), .B1(new_n930), .B2(new_n581), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n932), .A2(new_n362), .A3(new_n666), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n941), .B(KEYINPUT60), .ZN(G1350gat));
  NAND2_X1  g741(.A1(new_n936), .A2(new_n665), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT124), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(KEYINPUT61), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n943), .A2(G190gat), .A3(new_n945), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n944), .A2(KEYINPUT61), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n932), .A2(new_n343), .A3(new_n698), .ZN(new_n949));
  INV_X1    g748(.A(new_n947), .ZN(new_n950));
  NAND4_X1  g749(.A1(new_n943), .A2(G190gat), .A3(new_n945), .A4(new_n950), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n948), .A2(new_n949), .A3(new_n951), .ZN(G1351gat));
  NOR3_X1   g751(.A1(new_n658), .A2(new_n385), .A3(new_n741), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n913), .A2(new_n914), .A3(new_n953), .ZN(new_n954));
  OAI21_X1  g753(.A(G197gat), .B1(new_n954), .B2(new_n554), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n836), .A2(new_n646), .ZN(new_n956));
  OAI21_X1  g755(.A(KEYINPUT125), .B1(new_n870), .B2(new_n385), .ZN(new_n957));
  OR3_X1    g756(.A1(new_n870), .A2(KEYINPUT125), .A3(new_n385), .ZN(new_n958));
  AND3_X1   g757(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  INV_X1    g758(.A(G197gat), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n959), .A2(new_n960), .A3(new_n555), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n955), .A2(new_n961), .ZN(G1352gat));
  INV_X1    g761(.A(KEYINPUT126), .ZN(new_n963));
  NAND4_X1  g762(.A1(new_n959), .A2(new_n963), .A3(new_n632), .A4(new_n639), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT62), .ZN(new_n965));
  NAND4_X1  g764(.A1(new_n956), .A2(new_n632), .A3(new_n957), .A4(new_n958), .ZN(new_n966));
  OAI21_X1  g765(.A(KEYINPUT126), .B1(new_n966), .B2(new_n640), .ZN(new_n967));
  AND3_X1   g766(.A1(new_n964), .A2(new_n965), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n965), .B1(new_n964), .B2(new_n967), .ZN(new_n969));
  AND2_X1   g768(.A1(new_n915), .A2(new_n953), .ZN(new_n970));
  OAI22_X1  g769(.A1(new_n968), .A2(new_n969), .B1(new_n632), .B2(new_n970), .ZN(G1353gat));
  NAND4_X1  g770(.A1(new_n913), .A2(new_n914), .A3(new_n666), .A4(new_n953), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n972), .A2(G211gat), .ZN(new_n973));
  INV_X1    g772(.A(KEYINPUT63), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n972), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n975), .A2(KEYINPUT127), .A3(new_n976), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n959), .A2(new_n302), .A3(new_n666), .ZN(new_n978));
  INV_X1    g777(.A(KEYINPUT127), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n973), .A2(new_n979), .A3(new_n974), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n977), .A2(new_n978), .A3(new_n980), .ZN(G1354gat));
  NOR3_X1   g780(.A1(new_n954), .A2(new_n303), .A3(new_n664), .ZN(new_n982));
  AOI21_X1  g781(.A(G218gat), .B1(new_n959), .B2(new_n698), .ZN(new_n983));
  NOR2_X1   g782(.A1(new_n982), .A2(new_n983), .ZN(G1355gat));
endmodule


