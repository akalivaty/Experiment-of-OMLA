//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 1 0 1 0 0 1 0 1 1 0 1 1 1 1 0 0 1 1 0 1 1 0 1 1 1 1 0 0 0 1 1 0 0 1 0 1 0 1 1 0 1 0 1 0 1 0 1 1 0 0 0 0 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n736, new_n737, new_n739, new_n740, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n807, new_n808, new_n809, new_n811, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n908, new_n910, new_n911, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n968, new_n969, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n982, new_n983,
    new_n984, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1030, new_n1031, new_n1032;
  INV_X1    g000(.A(KEYINPUT76), .ZN(new_n202));
  NAND2_X1  g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203));
  INV_X1    g002(.A(G155gat), .ZN(new_n204));
  INV_X1    g003(.A(G162gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n203), .B1(new_n206), .B2(KEYINPUT2), .ZN(new_n207));
  XOR2_X1   g006(.A(G141gat), .B(G148gat), .Z(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G141gat), .ZN(new_n210));
  INV_X1    g009(.A(G148gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT2), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(KEYINPUT75), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT75), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(KEYINPUT2), .ZN(new_n216));
  NAND2_X1  g015(.A1(G141gat), .A2(G148gat), .ZN(new_n217));
  NAND4_X1  g016(.A1(new_n212), .A2(new_n214), .A3(new_n216), .A4(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n203), .A2(KEYINPUT74), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(new_n206), .ZN(new_n221));
  NOR2_X1   g020(.A1(G155gat), .A2(G162gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(KEYINPUT74), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n209), .B1(new_n219), .B2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(G197gat), .ZN(new_n226));
  INV_X1    g025(.A(G204gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(G197gat), .A2(G204gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(G211gat), .A2(G218gat), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT22), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n230), .A2(new_n233), .ZN(new_n234));
  AND2_X1   g033(.A1(G211gat), .A2(G218gat), .ZN(new_n235));
  NOR2_X1   g034(.A1(G211gat), .A2(G218gat), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT69), .ZN(new_n237));
  NOR3_X1   g036(.A1(new_n235), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n234), .A2(new_n238), .ZN(new_n239));
  AOI22_X1  g038(.A1(new_n228), .A2(new_n229), .B1(new_n232), .B2(new_n231), .ZN(new_n240));
  INV_X1    g039(.A(new_n236), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n241), .A2(KEYINPUT69), .A3(new_n231), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  AOI21_X1  g042(.A(KEYINPUT29), .B1(new_n239), .B2(new_n243), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n225), .B1(new_n244), .B2(KEYINPUT3), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT74), .ZN(new_n246));
  NOR3_X1   g045(.A1(new_n246), .A2(G155gat), .A3(G162gat), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n247), .B1(new_n206), .B2(new_n220), .ZN(new_n248));
  AOI22_X1  g047(.A1(new_n248), .A2(new_n218), .B1(new_n207), .B2(new_n208), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT3), .ZN(new_n250));
  AOI21_X1  g049(.A(KEYINPUT29), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n239), .A2(new_n243), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n245), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(G228gat), .ZN(new_n254));
  INV_X1    g053(.A(G233gat), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT29), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n257), .B1(new_n225), .B2(KEYINPUT3), .ZN(new_n258));
  INV_X1    g057(.A(new_n252), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n235), .A2(new_n236), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n240), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n257), .B1(new_n240), .B2(new_n261), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n250), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n256), .B1(new_n265), .B2(new_n225), .ZN(new_n266));
  AOI22_X1  g065(.A1(new_n253), .A2(new_n256), .B1(new_n260), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(G22gat), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n202), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(G78gat), .ZN(new_n270));
  INV_X1    g069(.A(new_n256), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n271), .B1(new_n260), .B2(new_n245), .ZN(new_n272));
  INV_X1    g071(.A(new_n261), .ZN(new_n273));
  AOI21_X1  g072(.A(KEYINPUT29), .B1(new_n234), .B2(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(KEYINPUT3), .B1(new_n274), .B2(new_n262), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n271), .B1(new_n275), .B2(new_n249), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n248), .A2(new_n218), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n277), .A2(new_n250), .A3(new_n209), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n252), .B1(new_n278), .B2(new_n257), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  OAI21_X1  g079(.A(G22gat), .B1(new_n272), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n269), .A2(new_n270), .A3(new_n281), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n234), .A2(new_n238), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n240), .A2(new_n242), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n257), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n249), .B1(new_n285), .B2(new_n250), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n256), .B1(new_n286), .B2(new_n279), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n260), .A2(new_n266), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n287), .A2(new_n268), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(KEYINPUT76), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n268), .B1(new_n287), .B2(new_n288), .ZN(new_n291));
  OAI21_X1  g090(.A(G78gat), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(KEYINPUT31), .B(G50gat), .ZN(new_n293));
  INV_X1    g092(.A(G106gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n293), .B(new_n294), .ZN(new_n295));
  AND3_X1   g094(.A1(new_n282), .A2(new_n292), .A3(new_n295), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n295), .B1(new_n282), .B2(new_n292), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  XOR2_X1   g097(.A(G8gat), .B(G36gat), .Z(new_n299));
  XNOR2_X1  g098(.A(new_n299), .B(KEYINPUT71), .ZN(new_n300));
  XNOR2_X1  g099(.A(G64gat), .B(G92gat), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n300), .B(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(G226gat), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n304), .A2(new_n255), .ZN(new_n305));
  INV_X1    g104(.A(G183gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(KEYINPUT27), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT27), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(G183gat), .ZN(new_n309));
  INV_X1    g108(.A(G190gat), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n307), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT28), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  XNOR2_X1  g112(.A(KEYINPUT27), .B(G183gat), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n314), .A2(KEYINPUT28), .A3(new_n310), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(G169gat), .ZN(new_n317));
  INV_X1    g116(.A(G176gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT26), .ZN(new_n320));
  NAND2_X1  g119(.A1(G169gat), .A2(G176gat), .ZN(new_n321));
  AND3_X1   g120(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(G183gat), .A2(G190gat), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n323), .B1(new_n319), .B2(new_n320), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n316), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT23), .ZN(new_n327));
  NOR3_X1   g126(.A1(new_n327), .A2(G169gat), .A3(G176gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n321), .A2(KEYINPUT23), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n328), .B1(new_n319), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT24), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n323), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n306), .A2(new_n310), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(KEYINPUT25), .B1(new_n330), .B2(new_n335), .ZN(new_n336));
  NOR2_X1   g135(.A1(G169gat), .A2(G176gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(KEYINPUT23), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n327), .B1(G169gat), .B2(G176gat), .ZN(new_n339));
  OAI211_X1 g138(.A(KEYINPUT25), .B(new_n338), .C1(new_n339), .C2(new_n337), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT65), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n323), .A2(new_n341), .A3(new_n331), .ZN(new_n342));
  OAI211_X1 g141(.A(G183gat), .B(G190gat), .C1(KEYINPUT65), .C2(KEYINPUT24), .ZN(new_n343));
  AND3_X1   g142(.A1(new_n342), .A2(new_n334), .A3(new_n343), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n340), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n326), .B1(new_n336), .B2(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n305), .B1(new_n346), .B2(new_n257), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT25), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n338), .B1(new_n339), .B2(new_n337), .ZN(new_n349));
  AND3_X1   g148(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n348), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n342), .A2(new_n334), .A3(new_n343), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n330), .A2(new_n352), .A3(KEYINPUT25), .ZN(new_n353));
  AOI22_X1  g152(.A1(new_n351), .A2(new_n353), .B1(new_n316), .B2(new_n325), .ZN(new_n354));
  INV_X1    g153(.A(new_n305), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NOR3_X1   g155(.A1(new_n347), .A2(new_n356), .A3(new_n259), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n355), .B1(new_n354), .B2(KEYINPUT29), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n346), .A2(new_n305), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n252), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT70), .ZN(new_n361));
  NOR3_X1   g160(.A1(new_n357), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n259), .B1(new_n347), .B2(new_n356), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n358), .A2(new_n359), .A3(new_n252), .ZN(new_n364));
  AOI21_X1  g163(.A(KEYINPUT70), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n303), .B1(new_n362), .B2(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n363), .A2(new_n302), .A3(new_n364), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT30), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n367), .A2(KEYINPUT73), .A3(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(KEYINPUT73), .B1(new_n367), .B2(new_n368), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n366), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n363), .A2(KEYINPUT30), .A3(new_n364), .A4(new_n302), .ZN(new_n373));
  XNOR2_X1  g172(.A(new_n373), .B(KEYINPUT72), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(G113gat), .ZN(new_n376));
  INV_X1    g175(.A(G120gat), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT1), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n379), .B1(G113gat), .B2(G120gat), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(G127gat), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n382), .A2(G134gat), .ZN(new_n383));
  INV_X1    g182(.A(G134gat), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n384), .A2(G127gat), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n381), .A2(new_n386), .ZN(new_n387));
  OAI22_X1  g186(.A1(new_n378), .A2(new_n380), .B1(new_n383), .B2(new_n385), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n249), .B(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(G225gat), .A2(G233gat), .ZN(new_n391));
  OAI21_X1  g190(.A(KEYINPUT5), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n225), .A2(KEYINPUT3), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n393), .A2(new_n278), .A3(new_n389), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n225), .A2(new_n389), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(KEYINPUT4), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT4), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n397), .B1(new_n225), .B2(new_n389), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n394), .A2(new_n396), .A3(new_n391), .A4(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n392), .A2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n389), .ZN(new_n401));
  AOI21_X1  g200(.A(KEYINPUT4), .B1(new_n401), .B2(new_n249), .ZN(new_n402));
  NOR3_X1   g201(.A1(new_n225), .A2(new_n389), .A3(new_n397), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n404), .A2(KEYINPUT5), .A3(new_n391), .A4(new_n394), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n400), .A2(new_n405), .ZN(new_n406));
  XNOR2_X1  g205(.A(G1gat), .B(G29gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(new_n407), .B(KEYINPUT0), .ZN(new_n408));
  XNOR2_X1  g207(.A(G57gat), .B(G85gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n408), .B(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n406), .A2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT6), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n400), .A2(new_n410), .A3(new_n405), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n400), .A2(KEYINPUT6), .A3(new_n405), .A4(new_n410), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n298), .A2(new_n375), .A3(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT72), .ZN(new_n419));
  AND2_X1   g218(.A1(new_n373), .A2(new_n419), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n373), .A2(new_n419), .ZN(new_n421));
  OAI221_X1 g220(.A(new_n366), .B1(new_n420), .B2(new_n421), .C1(new_n371), .C2(new_n370), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT40), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n394), .A2(new_n396), .A3(new_n398), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT39), .ZN(new_n425));
  INV_X1    g224(.A(new_n391), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n424), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(new_n411), .ZN(new_n428));
  XNOR2_X1  g227(.A(new_n225), .B(new_n389), .ZN(new_n429));
  OAI21_X1  g228(.A(KEYINPUT39), .B1(new_n429), .B2(new_n426), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n430), .B1(new_n426), .B2(new_n424), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n423), .B1(new_n428), .B2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n430), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n424), .A2(new_n426), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n435), .A2(KEYINPUT40), .A3(new_n411), .A4(new_n427), .ZN(new_n436));
  AND3_X1   g235(.A1(new_n432), .A2(new_n414), .A3(new_n436), .ZN(new_n437));
  AND3_X1   g236(.A1(new_n415), .A2(new_n416), .A3(new_n367), .ZN(new_n438));
  OAI21_X1  g237(.A(KEYINPUT37), .B1(new_n357), .B2(new_n360), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT37), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n363), .A2(new_n440), .A3(new_n364), .ZN(new_n441));
  AND3_X1   g240(.A1(new_n439), .A2(new_n303), .A3(new_n441), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n361), .B1(new_n357), .B2(new_n360), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n363), .A2(KEYINPUT70), .A3(new_n364), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n440), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n441), .A2(KEYINPUT38), .A3(new_n303), .ZN(new_n446));
  OAI22_X1  g245(.A1(new_n442), .A2(KEYINPUT38), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  AOI22_X1  g246(.A1(new_n422), .A2(new_n437), .B1(new_n438), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n418), .B1(new_n448), .B2(new_n298), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n346), .A2(new_n389), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n354), .A2(new_n401), .ZN(new_n451));
  NAND2_X1  g250(.A1(G227gat), .A2(G233gat), .ZN(new_n452));
  XNOR2_X1  g251(.A(new_n452), .B(KEYINPUT64), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n450), .A2(new_n451), .A3(new_n454), .ZN(new_n455));
  OAI21_X1  g254(.A(KEYINPUT34), .B1(new_n453), .B2(KEYINPUT67), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n450), .A2(new_n451), .A3(new_n454), .A4(new_n456), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  XNOR2_X1  g259(.A(G15gat), .B(G43gat), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT66), .ZN(new_n462));
  XNOR2_X1  g261(.A(new_n461), .B(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(G71gat), .ZN(new_n464));
  XNOR2_X1  g263(.A(new_n461), .B(KEYINPUT66), .ZN(new_n465));
  INV_X1    g264(.A(G71gat), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(G99gat), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n464), .A2(new_n467), .A3(G99gat), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n346), .A2(new_n389), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n354), .A2(new_n401), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n453), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT33), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n472), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n460), .A2(new_n477), .ZN(new_n478));
  AND2_X1   g277(.A1(new_n470), .A2(new_n471), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n454), .B1(new_n450), .B2(new_n451), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n479), .B1(new_n480), .B2(KEYINPUT33), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n481), .A2(new_n459), .A3(new_n458), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n475), .A2(KEYINPUT32), .ZN(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  AND3_X1   g283(.A1(new_n478), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n484), .B1(new_n478), .B2(new_n482), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT36), .ZN(new_n488));
  AND2_X1   g287(.A1(new_n488), .A2(KEYINPUT68), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n488), .A2(KEYINPUT68), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n487), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n478), .A2(new_n482), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(new_n483), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n478), .A2(new_n482), .A3(new_n484), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n495), .B1(KEYINPUT68), .B2(new_n488), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n491), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n282), .A2(new_n292), .A3(new_n295), .ZN(new_n498));
  INV_X1    g297(.A(new_n295), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n270), .B1(new_n269), .B2(new_n281), .ZN(new_n500));
  AND4_X1   g299(.A1(KEYINPUT76), .A2(new_n281), .A3(new_n270), .A4(new_n289), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n495), .B1(new_n498), .B2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT35), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n503), .A2(new_n504), .A3(new_n417), .A4(new_n375), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n502), .A2(new_n498), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n375), .A2(new_n506), .A3(new_n417), .A4(new_n487), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(KEYINPUT35), .ZN(new_n508));
  AOI22_X1  g307(.A1(new_n449), .A2(new_n497), .B1(new_n505), .B2(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(G15gat), .B(G22gat), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT16), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n510), .B1(new_n511), .B2(G1gat), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n512), .B1(G1gat), .B2(new_n510), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n513), .B(G8gat), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT14), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n515), .B1(G29gat), .B2(G36gat), .ZN(new_n516));
  INV_X1    g315(.A(G29gat), .ZN(new_n517));
  INV_X1    g316(.A(G36gat), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n517), .A2(new_n518), .A3(KEYINPUT14), .ZN(new_n519));
  XNOR2_X1  g318(.A(G43gat), .B(G50gat), .ZN(new_n520));
  XNOR2_X1  g319(.A(KEYINPUT79), .B(KEYINPUT15), .ZN(new_n521));
  OAI211_X1 g320(.A(new_n516), .B(new_n519), .C1(new_n520), .C2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(G50gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(G43gat), .ZN(new_n524));
  INV_X1    g323(.A(G43gat), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(G50gat), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n524), .A2(new_n526), .A3(KEYINPUT15), .ZN(new_n527));
  XNOR2_X1  g326(.A(KEYINPUT78), .B(G29gat), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n527), .B1(new_n528), .B2(new_n518), .ZN(new_n529));
  OAI21_X1  g328(.A(KEYINPUT80), .B1(new_n522), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n519), .A2(new_n516), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n524), .A2(new_n526), .ZN(new_n532));
  XOR2_X1   g331(.A(KEYINPUT79), .B(KEYINPUT15), .Z(new_n533));
  AOI21_X1  g332(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n517), .A2(KEYINPUT78), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT78), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(G29gat), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  AOI22_X1  g337(.A1(G36gat), .A2(new_n538), .B1(new_n520), .B2(KEYINPUT15), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT80), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n534), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n527), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n531), .A2(KEYINPUT77), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n538), .A2(G36gat), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT77), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n519), .A2(new_n516), .A3(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n543), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  AOI22_X1  g346(.A1(new_n530), .A2(new_n541), .B1(new_n542), .B2(new_n547), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n514), .B1(new_n548), .B2(KEYINPUT17), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT81), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n530), .A2(new_n541), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n547), .A2(new_n542), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT17), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n550), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NOR3_X1   g354(.A1(new_n548), .A2(KEYINPUT81), .A3(KEYINPUT17), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n549), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(G229gat), .A2(G233gat), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n553), .A2(new_n514), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT82), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n553), .A2(new_n550), .A3(new_n554), .ZN(new_n563));
  OAI21_X1  g362(.A(KEYINPUT81), .B1(new_n548), .B2(KEYINPUT17), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AOI22_X1  g364(.A1(new_n565), .A2(new_n549), .B1(new_n553), .B2(new_n514), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n566), .A2(KEYINPUT82), .A3(new_n558), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT18), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n562), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND4_X1  g368(.A1(new_n557), .A2(KEYINPUT18), .A3(new_n558), .A4(new_n559), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT83), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n566), .A2(KEYINPUT83), .A3(KEYINPUT18), .A4(new_n558), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(G113gat), .B(G141gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(G197gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(KEYINPUT11), .B(G169gat), .ZN(new_n577));
  XOR2_X1   g376(.A(new_n576), .B(new_n577), .Z(new_n578));
  XOR2_X1   g377(.A(new_n578), .B(KEYINPUT12), .Z(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n514), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(new_n548), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(new_n559), .ZN(new_n583));
  XOR2_X1   g382(.A(new_n558), .B(KEYINPUT13), .Z(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g384(.A1(new_n569), .A2(new_n574), .A3(new_n580), .A4(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT84), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(KEYINPUT18), .B1(new_n560), .B2(new_n561), .ZN(new_n589));
  AOI22_X1  g388(.A1(new_n589), .A2(new_n567), .B1(new_n583), .B2(new_n584), .ZN(new_n590));
  NAND4_X1  g389(.A1(new_n590), .A2(KEYINPUT84), .A3(new_n580), .A4(new_n574), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n574), .ZN(new_n592));
  AOI22_X1  g391(.A1(new_n588), .A2(new_n591), .B1(new_n579), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n509), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT91), .ZN(new_n595));
  XNOR2_X1  g394(.A(G190gat), .B(G218gat), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT88), .ZN(new_n598));
  NAND2_X1  g397(.A1(G85gat), .A2(G92gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(KEYINPUT7), .ZN(new_n600));
  XNOR2_X1  g399(.A(G99gat), .B(G106gat), .ZN(new_n601));
  NAND2_X1  g400(.A1(G99gat), .A2(G106gat), .ZN(new_n602));
  INV_X1    g401(.A(G85gat), .ZN(new_n603));
  INV_X1    g402(.A(G92gat), .ZN(new_n604));
  AOI22_X1  g403(.A1(KEYINPUT8), .A2(new_n602), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  AND3_X1   g404(.A1(new_n600), .A2(new_n601), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n601), .B1(new_n600), .B2(new_n605), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n598), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n600), .A2(new_n605), .ZN(new_n609));
  INV_X1    g408(.A(new_n601), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n600), .A2(new_n601), .A3(new_n605), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n611), .A2(KEYINPUT88), .A3(new_n612), .ZN(new_n613));
  AND2_X1   g412(.A1(new_n608), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n614), .B1(new_n553), .B2(new_n554), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n615), .B1(new_n564), .B2(new_n563), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT41), .ZN(new_n617));
  NAND2_X1  g416(.A1(G232gat), .A2(G233gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(KEYINPUT86), .ZN(new_n619));
  OAI22_X1  g418(.A1(new_n614), .A2(new_n548), .B1(new_n617), .B2(new_n619), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n597), .B1(new_n616), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n619), .A2(new_n617), .ZN(new_n622));
  XOR2_X1   g421(.A(new_n622), .B(KEYINPUT87), .Z(new_n623));
  XNOR2_X1  g422(.A(G134gat), .B(G162gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n620), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n555), .A2(new_n556), .ZN(new_n627));
  OAI211_X1 g426(.A(new_n626), .B(new_n596), .C1(new_n627), .C2(new_n615), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n621), .A2(new_n625), .A3(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT89), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n621), .A2(new_n628), .ZN(new_n632));
  INV_X1    g431(.A(new_n625), .ZN(new_n633));
  AOI21_X1  g432(.A(KEYINPUT90), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT90), .ZN(new_n635));
  AOI211_X1 g434(.A(new_n635), .B(new_n625), .C1(new_n621), .C2(new_n628), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n595), .B1(new_n631), .B2(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n629), .B(KEYINPUT89), .ZN(new_n639));
  OAI211_X1 g438(.A(new_n639), .B(KEYINPUT91), .C1(new_n634), .C2(new_n636), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g440(.A(G57gat), .B(G64gat), .Z(new_n642));
  NAND2_X1  g441(.A1(new_n466), .A2(new_n270), .ZN(new_n643));
  NAND2_X1  g442(.A1(G71gat), .A2(G78gat), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT9), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n642), .A2(new_n645), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(G57gat), .B(G64gat), .ZN(new_n649));
  OAI211_X1 g448(.A(new_n644), .B(new_n643), .C1(new_n649), .C2(new_n646), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT85), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n648), .A2(new_n650), .A3(KEYINPUT85), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  OR2_X1    g454(.A1(new_n655), .A2(KEYINPUT21), .ZN(new_n656));
  NAND2_X1  g455(.A1(G231gat), .A2(G233gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(G127gat), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n655), .A2(KEYINPUT21), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n581), .A2(new_n660), .ZN(new_n661));
  OR2_X1    g460(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n659), .A2(new_n661), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g463(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(new_n204), .ZN(new_n666));
  XNOR2_X1  g465(.A(G183gat), .B(G211gat), .ZN(new_n667));
  XOR2_X1   g466(.A(new_n666), .B(new_n667), .Z(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n664), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n662), .A2(new_n663), .A3(new_n668), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n641), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n608), .A2(new_n613), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n674), .A2(KEYINPUT10), .A3(new_n655), .ZN(new_n675));
  AND3_X1   g474(.A1(new_n648), .A2(new_n650), .A3(KEYINPUT85), .ZN(new_n676));
  AOI21_X1  g475(.A(KEYINPUT85), .B1(new_n648), .B2(new_n650), .ZN(new_n677));
  OAI22_X1  g476(.A1(new_n676), .A2(new_n677), .B1(new_n606), .B2(new_n607), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n611), .A2(new_n651), .A3(new_n612), .ZN(new_n679));
  AND2_X1   g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  OAI211_X1 g479(.A(KEYINPUT92), .B(new_n675), .C1(new_n680), .C2(KEYINPUT10), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT92), .ZN(new_n682));
  AND3_X1   g481(.A1(new_n674), .A2(KEYINPUT10), .A3(new_n655), .ZN(new_n683));
  AOI21_X1  g482(.A(KEYINPUT10), .B1(new_n678), .B2(new_n679), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n682), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(G230gat), .A2(G233gat), .ZN(new_n686));
  XOR2_X1   g485(.A(new_n686), .B(KEYINPUT93), .Z(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n681), .A2(new_n685), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n680), .A2(new_n687), .ZN(new_n690));
  XNOR2_X1  g489(.A(G120gat), .B(G148gat), .ZN(new_n691));
  XNOR2_X1  g490(.A(G176gat), .B(G204gat), .ZN(new_n692));
  XOR2_X1   g491(.A(new_n691), .B(new_n692), .Z(new_n693));
  AND2_X1   g492(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n689), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n688), .B1(new_n683), .B2(new_n684), .ZN(new_n696));
  AND2_X1   g495(.A1(new_n696), .A2(new_n690), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n695), .B1(new_n697), .B2(new_n693), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n673), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n594), .A2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT94), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n594), .A2(KEYINPUT94), .A3(new_n699), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n417), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(G1gat), .ZN(G1324gat));
  INV_X1    g506(.A(new_n704), .ZN(new_n708));
  OAI211_X1 g507(.A(KEYINPUT97), .B(G8gat), .C1(new_n708), .C2(new_n375), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT97), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n375), .B1(new_n702), .B2(new_n703), .ZN(new_n711));
  INV_X1    g510(.A(G8gat), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n710), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n709), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(KEYINPUT16), .B(G8gat), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT42), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n711), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(KEYINPUT98), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT98), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n711), .A2(new_n720), .A3(new_n717), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n714), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n715), .B(KEYINPUT95), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n704), .A2(new_n422), .A3(new_n724), .ZN(new_n725));
  AND3_X1   g524(.A1(new_n725), .A2(KEYINPUT96), .A3(new_n716), .ZN(new_n726));
  AOI21_X1  g525(.A(KEYINPUT96), .B1(new_n725), .B2(new_n716), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(KEYINPUT99), .B1(new_n723), .B2(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(KEYINPUT42), .B1(new_n711), .B2(new_n724), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(KEYINPUT96), .ZN(new_n731));
  AOI22_X1  g530(.A1(new_n713), .A2(new_n709), .B1(new_n719), .B2(new_n721), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT99), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n731), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n729), .A2(new_n734), .ZN(G1325gat));
  OR3_X1    g534(.A1(new_n708), .A2(G15gat), .A3(new_n495), .ZN(new_n736));
  OAI21_X1  g535(.A(G15gat), .B1(new_n708), .B2(new_n497), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(G1326gat));
  NAND2_X1  g537(.A1(new_n704), .A2(new_n298), .ZN(new_n739));
  XNOR2_X1  g538(.A(KEYINPUT43), .B(G22gat), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n739), .B(new_n740), .ZN(G1327gat));
  INV_X1    g540(.A(new_n641), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n672), .A2(new_n698), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(KEYINPUT100), .ZN(new_n745));
  AND2_X1   g544(.A1(new_n745), .A2(new_n594), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n746), .A2(new_n705), .A3(new_n528), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(KEYINPUT45), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT101), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n505), .A2(new_n508), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n438), .A2(new_n447), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n437), .B1(new_n372), .B2(new_n374), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n298), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n502), .A2(new_n417), .A3(new_n498), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n754), .A2(new_n422), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n497), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n641), .B1(new_n750), .B2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT44), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n749), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  OAI211_X1 g558(.A(KEYINPUT101), .B(KEYINPUT44), .C1(new_n509), .C2(new_n641), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n509), .A2(KEYINPUT102), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n750), .A2(new_n756), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT102), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g564(.A(KEYINPUT103), .B(KEYINPUT44), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n762), .A2(new_n765), .A3(new_n742), .A4(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n761), .A2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(new_n593), .ZN(new_n769));
  AND3_X1   g568(.A1(new_n768), .A2(new_n769), .A3(new_n743), .ZN(new_n770));
  AND2_X1   g569(.A1(new_n770), .A2(new_n705), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n748), .B1(new_n528), .B2(new_n771), .ZN(G1328gat));
  AOI21_X1  g571(.A(new_n518), .B1(new_n770), .B2(new_n422), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n745), .A2(new_n518), .A3(new_n422), .A4(new_n594), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(KEYINPUT46), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT104), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n776), .B(new_n777), .ZN(G1329gat));
  INV_X1    g577(.A(KEYINPUT47), .ZN(new_n779));
  INV_X1    g578(.A(new_n497), .ZN(new_n780));
  AND2_X1   g579(.A1(new_n770), .A2(new_n780), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n781), .A2(new_n525), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n746), .A2(new_n525), .A3(new_n487), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(KEYINPUT105), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n779), .B1(new_n782), .B2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT105), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n783), .B(new_n786), .ZN(new_n787));
  OAI211_X1 g586(.A(new_n787), .B(KEYINPUT47), .C1(new_n525), .C2(new_n781), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n785), .A2(new_n788), .ZN(G1330gat));
  AND3_X1   g588(.A1(new_n746), .A2(new_n523), .A3(new_n298), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n770), .A2(new_n298), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n790), .B1(new_n791), .B2(G50gat), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT48), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n793), .B1(new_n790), .B2(KEYINPUT106), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n792), .B(new_n794), .ZN(G1331gat));
  NAND2_X1  g594(.A1(new_n762), .A2(new_n765), .ZN(new_n796));
  INV_X1    g595(.A(new_n698), .ZN(new_n797));
  NOR4_X1   g596(.A1(new_n796), .A2(new_n769), .A3(new_n673), .A4(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(new_n705), .ZN(new_n799));
  XNOR2_X1  g598(.A(KEYINPUT107), .B(G57gat), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n799), .B(new_n800), .ZN(G1332gat));
  NAND2_X1  g600(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n802));
  AND3_X1   g601(.A1(new_n798), .A2(new_n422), .A3(new_n802), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n803), .B(KEYINPUT108), .ZN(new_n804));
  OR2_X1    g603(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n805));
  XNOR2_X1  g604(.A(new_n804), .B(new_n805), .ZN(G1333gat));
  NAND3_X1  g605(.A1(new_n798), .A2(G71gat), .A3(new_n780), .ZN(new_n807));
  AND2_X1   g606(.A1(new_n798), .A2(new_n487), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n807), .B1(new_n808), .B2(G71gat), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n809), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g609(.A1(new_n798), .A2(new_n298), .ZN(new_n811));
  XNOR2_X1  g610(.A(new_n811), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g611(.A1(new_n769), .A2(new_n672), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n757), .A2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT51), .ZN(new_n815));
  OR3_X1    g614(.A1(new_n814), .A2(KEYINPUT110), .A3(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(KEYINPUT110), .B1(new_n814), .B2(new_n815), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n814), .A2(new_n815), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n816), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n819), .A2(new_n603), .A3(new_n705), .A4(new_n698), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n813), .A2(new_n698), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n768), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n823), .A2(new_n417), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n824), .A2(KEYINPUT109), .ZN(new_n825));
  OAI21_X1  g624(.A(G85gat), .B1(new_n824), .B2(KEYINPUT109), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n820), .B1(new_n825), .B2(new_n826), .ZN(G1336gat));
  NOR3_X1   g626(.A1(new_n375), .A2(G92gat), .A3(new_n797), .ZN(new_n828));
  AOI21_X1  g627(.A(KEYINPUT52), .B1(new_n819), .B2(new_n828), .ZN(new_n829));
  AOI211_X1 g628(.A(new_n375), .B(new_n821), .C1(new_n761), .C2(new_n767), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n829), .B1(new_n604), .B2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT111), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n832), .B1(new_n830), .B2(new_n604), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n768), .A2(new_n422), .A3(new_n822), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n834), .A2(KEYINPUT111), .A3(G92gat), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT112), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n814), .B1(new_n836), .B2(new_n815), .ZN(new_n837));
  AOI211_X1 g636(.A(KEYINPUT112), .B(KEYINPUT51), .C1(new_n757), .C2(new_n813), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n828), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n833), .A2(new_n835), .A3(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT113), .ZN(new_n841));
  AND3_X1   g640(.A1(new_n840), .A2(new_n841), .A3(KEYINPUT52), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n841), .B1(new_n840), .B2(KEYINPUT52), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n831), .B1(new_n842), .B2(new_n843), .ZN(G1337gat));
  INV_X1    g643(.A(KEYINPUT116), .ZN(new_n845));
  OAI21_X1  g644(.A(KEYINPUT114), .B1(new_n823), .B2(new_n497), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT114), .ZN(new_n847));
  NAND4_X1  g646(.A1(new_n768), .A2(new_n847), .A3(new_n780), .A4(new_n822), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  XOR2_X1   g648(.A(KEYINPUT115), .B(G99gat), .Z(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n797), .A2(new_n495), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n851), .B1(new_n819), .B2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n845), .B1(new_n852), .B2(new_n855), .ZN(new_n856));
  AOI211_X1 g655(.A(KEYINPUT116), .B(new_n854), .C1(new_n849), .C2(new_n851), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n856), .A2(new_n857), .ZN(G1338gat));
  XOR2_X1   g657(.A(KEYINPUT119), .B(KEYINPUT53), .Z(new_n859));
  NOR3_X1   g658(.A1(new_n506), .A2(new_n797), .A3(G106gat), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n859), .B1(new_n819), .B2(new_n860), .ZN(new_n861));
  AOI211_X1 g660(.A(new_n506), .B(new_n821), .C1(new_n761), .C2(new_n767), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n861), .B1(new_n294), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(KEYINPUT117), .B1(new_n862), .B2(new_n294), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n768), .A2(new_n298), .A3(new_n822), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT117), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n865), .A2(new_n866), .A3(G106gat), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n860), .B1(new_n837), .B2(new_n838), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n864), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  AND3_X1   g668(.A1(new_n869), .A2(KEYINPUT118), .A3(KEYINPUT53), .ZN(new_n870));
  AOI21_X1  g669(.A(KEYINPUT118), .B1(new_n869), .B2(KEYINPUT53), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n863), .B1(new_n870), .B2(new_n871), .ZN(G1339gat));
  NOR3_X1   g671(.A1(new_n673), .A2(new_n769), .A3(new_n698), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n696), .A2(KEYINPUT54), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n875), .A2(new_n693), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT54), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n683), .A2(new_n684), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n877), .B1(new_n878), .B2(new_n687), .ZN(new_n879));
  AND3_X1   g678(.A1(new_n689), .A2(new_n879), .A3(KEYINPUT120), .ZN(new_n880));
  AOI21_X1  g679(.A(KEYINPUT120), .B1(new_n689), .B2(new_n879), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n876), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT55), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  OAI211_X1 g683(.A(KEYINPUT55), .B(new_n876), .C1(new_n880), .C2(new_n881), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n884), .A2(new_n695), .A3(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(new_n578), .ZN(new_n888));
  OR2_X1    g687(.A1(new_n566), .A2(new_n558), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n583), .A2(new_n584), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n888), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n892), .B1(new_n588), .B2(new_n591), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n887), .A2(new_n893), .A3(new_n640), .A4(new_n638), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n588), .A2(new_n591), .ZN(new_n896));
  INV_X1    g695(.A(new_n892), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n896), .A2(new_n698), .A3(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n898), .B1(new_n593), .B2(new_n886), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n742), .B1(new_n899), .B2(KEYINPUT121), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT121), .ZN(new_n901));
  OAI211_X1 g700(.A(new_n898), .B(new_n901), .C1(new_n593), .C2(new_n886), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n895), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n874), .B1(new_n903), .B2(new_n672), .ZN(new_n904));
  NAND4_X1  g703(.A1(new_n904), .A2(new_n705), .A3(new_n375), .A4(new_n503), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n905), .A2(new_n593), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n906), .B(new_n376), .ZN(G1340gat));
  NOR2_X1   g706(.A1(new_n905), .A2(new_n797), .ZN(new_n908));
  XNOR2_X1  g707(.A(new_n908), .B(new_n377), .ZN(G1341gat));
  INV_X1    g708(.A(new_n672), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n905), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g710(.A(new_n911), .B(new_n382), .ZN(G1342gat));
  NOR2_X1   g711(.A1(new_n905), .A2(new_n641), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(new_n384), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(KEYINPUT56), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT56), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n913), .A2(new_n916), .A3(new_n384), .ZN(new_n917));
  OAI211_X1 g716(.A(new_n915), .B(new_n917), .C1(new_n913), .C2(new_n384), .ZN(G1343gat));
  INV_X1    g717(.A(KEYINPUT57), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n592), .A2(new_n579), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n886), .B1(new_n896), .B2(new_n920), .ZN(new_n921));
  AOI211_X1 g720(.A(new_n797), .B(new_n892), .C1(new_n588), .C2(new_n591), .ZN(new_n922));
  OAI21_X1  g721(.A(KEYINPUT121), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n923), .A2(new_n902), .A3(new_n641), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n672), .B1(new_n924), .B2(new_n894), .ZN(new_n925));
  OAI211_X1 g724(.A(new_n919), .B(new_n298), .C1(new_n925), .C2(new_n873), .ZN(new_n926));
  NOR3_X1   g725(.A1(new_n780), .A2(new_n417), .A3(new_n422), .ZN(new_n927));
  INV_X1    g726(.A(new_n927), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n641), .B1(new_n921), .B2(new_n922), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n672), .B1(new_n929), .B2(new_n894), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n298), .B1(new_n930), .B2(new_n873), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n928), .B1(new_n931), .B2(KEYINPUT57), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n926), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g732(.A(G141gat), .B1(new_n933), .B2(new_n593), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT58), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n924), .A2(new_n894), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(new_n910), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n417), .B1(new_n937), .B2(new_n874), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n497), .A2(new_n298), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n939), .A2(new_n422), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n769), .A2(new_n210), .ZN(new_n942));
  OAI211_X1 g741(.A(new_n934), .B(new_n935), .C1(new_n941), .C2(new_n942), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n941), .A2(new_n942), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n933), .A2(KEYINPUT122), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT122), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n926), .A2(new_n932), .A3(new_n946), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n945), .A2(new_n769), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n944), .B1(new_n948), .B2(G141gat), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n943), .B1(new_n949), .B2(new_n935), .ZN(G1344gat));
  INV_X1    g749(.A(new_n941), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n951), .A2(new_n211), .A3(new_n698), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT59), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(G148gat), .ZN(new_n954));
  AND3_X1   g753(.A1(new_n926), .A2(new_n932), .A3(new_n946), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n946), .B1(new_n926), .B2(new_n932), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n954), .B1(new_n957), .B2(new_n698), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n904), .A2(KEYINPUT57), .A3(new_n298), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n931), .A2(new_n919), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n961), .A2(new_n698), .A3(new_n927), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n953), .B1(new_n962), .B2(G148gat), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n952), .B1(new_n958), .B2(new_n963), .ZN(G1345gat));
  NAND3_X1  g763(.A1(new_n951), .A2(new_n204), .A3(new_n672), .ZN(new_n965));
  NOR3_X1   g764(.A1(new_n955), .A2(new_n956), .A3(new_n910), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n965), .B1(new_n966), .B2(new_n204), .ZN(G1346gat));
  AOI21_X1  g766(.A(G162gat), .B1(new_n951), .B2(new_n742), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n641), .A2(new_n205), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n968), .B1(new_n957), .B2(new_n969), .ZN(G1347gat));
  NAND4_X1  g769(.A1(new_n904), .A2(new_n417), .A3(new_n422), .A4(new_n503), .ZN(new_n971));
  NOR3_X1   g770(.A1(new_n971), .A2(new_n317), .A3(new_n593), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n503), .A2(new_n422), .ZN(new_n973));
  XOR2_X1   g772(.A(new_n973), .B(KEYINPUT123), .Z(new_n974));
  OAI211_X1 g773(.A(new_n417), .B(new_n974), .C1(new_n925), .C2(new_n873), .ZN(new_n975));
  INV_X1    g774(.A(new_n975), .ZN(new_n976));
  AOI21_X1  g775(.A(G169gat), .B1(new_n976), .B2(new_n769), .ZN(new_n977));
  NOR2_X1   g776(.A1(new_n972), .A2(new_n977), .ZN(G1348gat));
  OAI21_X1  g777(.A(G176gat), .B1(new_n971), .B2(new_n797), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n976), .A2(new_n318), .A3(new_n698), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n979), .A2(new_n980), .ZN(G1349gat));
  OAI21_X1  g780(.A(G183gat), .B1(new_n971), .B2(new_n910), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n976), .A2(new_n314), .A3(new_n672), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  XNOR2_X1  g783(.A(new_n984), .B(KEYINPUT60), .ZN(G1350gat));
  AOI21_X1  g784(.A(new_n705), .B1(new_n937), .B2(new_n874), .ZN(new_n986));
  NOR2_X1   g785(.A1(new_n641), .A2(G190gat), .ZN(new_n987));
  NAND4_X1  g786(.A1(new_n986), .A2(KEYINPUT124), .A3(new_n974), .A4(new_n987), .ZN(new_n988));
  INV_X1    g787(.A(KEYINPUT124), .ZN(new_n989));
  INV_X1    g788(.A(new_n987), .ZN(new_n990));
  OAI21_X1  g789(.A(new_n989), .B1(new_n975), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n988), .A2(new_n991), .ZN(new_n992));
  OAI211_X1 g791(.A(KEYINPUT61), .B(G190gat), .C1(new_n971), .C2(new_n641), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND4_X1  g793(.A1(new_n986), .A2(new_n422), .A3(new_n503), .A4(new_n742), .ZN(new_n995));
  AOI21_X1  g794(.A(KEYINPUT61), .B1(new_n995), .B2(G190gat), .ZN(new_n996));
  OAI21_X1  g795(.A(KEYINPUT125), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n995), .A2(G190gat), .ZN(new_n998));
  INV_X1    g797(.A(KEYINPUT61), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g799(.A(KEYINPUT125), .ZN(new_n1001));
  NAND4_X1  g800(.A1(new_n1000), .A2(new_n1001), .A3(new_n993), .A4(new_n992), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n997), .A2(new_n1002), .ZN(G1351gat));
  OAI211_X1 g802(.A(new_n417), .B(new_n422), .C1(new_n925), .C2(new_n873), .ZN(new_n1004));
  NOR2_X1   g803(.A1(new_n1004), .A2(new_n939), .ZN(new_n1005));
  NAND3_X1  g804(.A1(new_n1005), .A2(new_n226), .A3(new_n769), .ZN(new_n1006));
  NOR3_X1   g805(.A1(new_n780), .A2(new_n705), .A3(new_n375), .ZN(new_n1007));
  INV_X1    g806(.A(new_n1007), .ZN(new_n1008));
  AOI211_X1 g807(.A(new_n593), .B(new_n1008), .C1(new_n959), .C2(new_n960), .ZN(new_n1009));
  OAI21_X1  g808(.A(G197gat), .B1(new_n1009), .B2(KEYINPUT126), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n961), .A2(new_n1007), .ZN(new_n1011));
  INV_X1    g810(.A(KEYINPUT126), .ZN(new_n1012));
  NOR3_X1   g811(.A1(new_n1011), .A2(new_n1012), .A3(new_n593), .ZN(new_n1013));
  OAI21_X1  g812(.A(new_n1006), .B1(new_n1010), .B2(new_n1013), .ZN(G1352gat));
  NOR2_X1   g813(.A1(new_n797), .A2(G204gat), .ZN(new_n1015));
  NAND2_X1  g814(.A1(new_n1005), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g815(.A(KEYINPUT62), .ZN(new_n1017));
  XNOR2_X1  g816(.A(new_n1016), .B(new_n1017), .ZN(new_n1018));
  AOI211_X1 g817(.A(new_n797), .B(new_n1008), .C1(new_n959), .C2(new_n960), .ZN(new_n1019));
  INV_X1    g818(.A(KEYINPUT127), .ZN(new_n1020));
  OAI21_X1  g819(.A(G204gat), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  NOR3_X1   g820(.A1(new_n1011), .A2(KEYINPUT127), .A3(new_n797), .ZN(new_n1022));
  OAI21_X1  g821(.A(new_n1018), .B1(new_n1021), .B2(new_n1022), .ZN(G1353gat));
  INV_X1    g822(.A(G211gat), .ZN(new_n1024));
  NAND3_X1  g823(.A1(new_n1005), .A2(new_n1024), .A3(new_n672), .ZN(new_n1025));
  NAND3_X1  g824(.A1(new_n961), .A2(new_n672), .A3(new_n1007), .ZN(new_n1026));
  AND3_X1   g825(.A1(new_n1026), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1027));
  AOI21_X1  g826(.A(KEYINPUT63), .B1(new_n1026), .B2(G211gat), .ZN(new_n1028));
  OAI21_X1  g827(.A(new_n1025), .B1(new_n1027), .B2(new_n1028), .ZN(G1354gat));
  OAI21_X1  g828(.A(G218gat), .B1(new_n1011), .B2(new_n641), .ZN(new_n1030));
  INV_X1    g829(.A(G218gat), .ZN(new_n1031));
  NAND3_X1  g830(.A1(new_n1005), .A2(new_n1031), .A3(new_n742), .ZN(new_n1032));
  NAND2_X1  g831(.A1(new_n1030), .A2(new_n1032), .ZN(G1355gat));
endmodule


