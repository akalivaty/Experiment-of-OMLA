//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 1 0 1 1 0 0 0 0 1 0 0 0 0 1 0 1 0 1 0 0 1 1 0 0 0 0 0 0 0 0 0 1 1 0 1 1 0 1 0 0 1 1 0 0 1 0 0 1 1 1 1 0 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:37 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1287, new_n1288, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1367, new_n1368;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT64), .Z(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT0), .ZN(new_n210));
  OAI21_X1  g0010(.A(G50), .B1(G58), .B2(G68), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT65), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g0016(.A(KEYINPUT66), .B(G68), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G97), .A2(G257), .B1(G116), .B2(G270), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G58), .B2(G232), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G77), .A2(G244), .ZN(new_n224));
  NAND4_X1  g0024(.A1(new_n221), .A2(new_n222), .A3(new_n223), .A4(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n207), .B1(new_n220), .B2(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n210), .B(new_n216), .C1(new_n226), .C2(KEYINPUT1), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT2), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G226), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n231), .B(G232), .Z(new_n232));
  XOR2_X1   g0032(.A(G250), .B(G257), .Z(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n232), .B(new_n235), .Z(G358));
  XNOR2_X1  g0036(.A(G87), .B(G97), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT67), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XOR2_X1   g0041(.A(G50), .B(G58), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G351));
  XNOR2_X1  g0044(.A(KEYINPUT3), .B(G33), .ZN(new_n245));
  NAND3_X1  g0045(.A1(new_n245), .A2(G223), .A3(G1698), .ZN(new_n246));
  INV_X1    g0046(.A(G1698), .ZN(new_n247));
  NAND3_X1  g0047(.A1(new_n245), .A2(G222), .A3(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(KEYINPUT3), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT3), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G77), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n246), .A2(new_n248), .A3(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT69), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  AND2_X1   g0057(.A1(G33), .A2(G41), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(new_n213), .ZN(new_n259));
  NAND4_X1  g0059(.A1(new_n246), .A2(new_n248), .A3(KEYINPUT69), .A4(new_n254), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n257), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT68), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n262), .B1(new_n258), .B2(new_n213), .ZN(new_n263));
  AND2_X1   g0063(.A1(G1), .A2(G13), .ZN(new_n264));
  NAND2_X1  g0064(.A1(G33), .A2(G41), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n264), .A2(KEYINPUT68), .A3(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G41), .ZN(new_n267));
  INV_X1    g0067(.A(G45), .ZN(new_n268));
  AOI21_X1  g0068(.A(G1), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND4_X1  g0069(.A1(new_n263), .A2(new_n266), .A3(G274), .A4(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G1), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n272), .B1(G41), .B2(G45), .ZN(new_n273));
  AND3_X1   g0073(.A1(new_n263), .A2(new_n273), .A3(new_n266), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n271), .B1(G226), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n261), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G169), .ZN(new_n277));
  INV_X1    g0077(.A(G179), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n277), .B1(new_n278), .B2(new_n276), .ZN(new_n279));
  NOR2_X1   g0079(.A1(G20), .A2(G33), .ZN(new_n280));
  AOI22_X1  g0080(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n280), .ZN(new_n281));
  XNOR2_X1  g0081(.A(KEYINPUT8), .B(G58), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n214), .A2(G33), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n281), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  OAI21_X1  g0084(.A(KEYINPUT70), .B1(new_n207), .B2(new_n249), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT70), .ZN(new_n286));
  NAND4_X1  g0086(.A1(new_n286), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n285), .A2(new_n213), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n284), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n288), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n272), .A2(G20), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n290), .A2(G50), .A3(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n272), .A2(G13), .A3(G20), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n202), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n289), .A2(new_n292), .A3(new_n295), .ZN(new_n296));
  AND2_X1   g0096(.A1(new_n279), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n290), .A2(new_n291), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(G77), .ZN(new_n300));
  NAND2_X1  g0100(.A1(G20), .A2(G77), .ZN(new_n301));
  INV_X1    g0101(.A(new_n280), .ZN(new_n302));
  XNOR2_X1  g0102(.A(KEYINPUT15), .B(G87), .ZN(new_n303));
  OAI221_X1 g0103(.A(new_n301), .B1(new_n282), .B2(new_n302), .C1(new_n283), .C2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(new_n288), .ZN(new_n305));
  INV_X1    g0105(.A(G77), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n294), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n300), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n271), .B1(G244), .B2(new_n274), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n245), .A2(G232), .A3(new_n247), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n245), .A2(G238), .A3(G1698), .ZN(new_n312));
  OR2_X1    g0112(.A1(KEYINPUT71), .A2(G107), .ZN(new_n313));
  NAND2_X1  g0113(.A1(KEYINPUT71), .A2(G107), .ZN(new_n314));
  AND2_X1   g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n311), .B(new_n312), .C1(new_n245), .C2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(new_n259), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n310), .A2(G179), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n310), .A2(new_n317), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(G169), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n309), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  XOR2_X1   g0122(.A(KEYINPUT72), .B(G200), .Z(new_n323));
  NAND2_X1  g0123(.A1(new_n319), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n324), .B1(G190), .B2(new_n319), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(new_n309), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n322), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT9), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n296), .A2(new_n328), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n289), .A2(KEYINPUT9), .A3(new_n292), .A4(new_n295), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n323), .B1(new_n261), .B2(new_n275), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT10), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n261), .A2(G190), .A3(new_n275), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n332), .A2(new_n334), .A3(new_n335), .A4(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT73), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n331), .A2(new_n333), .ZN(new_n340));
  NAND4_X1  g0140(.A1(new_n340), .A2(KEYINPUT73), .A3(new_n335), .A4(new_n336), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n340), .A2(new_n336), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(KEYINPUT10), .ZN(new_n344));
  AOI211_X1 g0144(.A(new_n297), .B(new_n327), .C1(new_n342), .C2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n274), .A2(G232), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(new_n270), .ZN(new_n347));
  INV_X1    g0147(.A(new_n259), .ZN(new_n348));
  OAI21_X1  g0148(.A(KEYINPUT80), .B1(new_n249), .B2(KEYINPUT3), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT80), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n350), .A2(new_n251), .A3(G33), .ZN(new_n351));
  AND3_X1   g0151(.A1(new_n349), .A2(new_n351), .A3(new_n250), .ZN(new_n352));
  MUX2_X1   g0152(.A(G223), .B(G226), .S(G1698), .Z(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(G33), .A2(G87), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n348), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n347), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(new_n278), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n358), .B1(G169), .B2(new_n357), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT16), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT7), .ZN(new_n361));
  NOR3_X1   g0161(.A1(new_n245), .A2(new_n361), .A3(G20), .ZN(new_n362));
  AOI21_X1  g0162(.A(KEYINPUT7), .B1(new_n253), .B2(new_n214), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n364), .A2(new_n218), .ZN(new_n365));
  INV_X1    g0165(.A(G159), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n302), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n201), .B1(new_n217), .B2(G58), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n368), .B1(new_n369), .B2(new_n214), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n360), .B1(new_n365), .B2(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n349), .A2(new_n351), .A3(new_n250), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(new_n214), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(KEYINPUT7), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n372), .A2(new_n361), .A3(new_n214), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n374), .A2(G68), .A3(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n370), .ZN(new_n377));
  AND4_X1   g0177(.A1(KEYINPUT81), .A2(new_n376), .A3(KEYINPUT16), .A4(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(G68), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n379), .B1(new_n373), .B2(KEYINPUT7), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n370), .B1(new_n380), .B2(new_n375), .ZN(new_n381));
  AOI21_X1  g0181(.A(KEYINPUT81), .B1(new_n381), .B2(KEYINPUT16), .ZN(new_n382));
  OAI211_X1 g0182(.A(new_n371), .B(new_n288), .C1(new_n378), .C2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(new_n282), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n384), .A2(new_n294), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n385), .B1(new_n298), .B2(new_n384), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n359), .B1(new_n383), .B2(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(KEYINPUT82), .B1(new_n388), .B2(KEYINPUT18), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(KEYINPUT18), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n376), .A2(new_n377), .A3(KEYINPUT16), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT81), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n381), .A2(KEYINPUT81), .A3(KEYINPUT16), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n290), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n386), .B1(new_n396), .B2(new_n371), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT82), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT18), .ZN(new_n399));
  NOR4_X1   g0199(.A1(new_n397), .A2(new_n398), .A3(new_n399), .A4(new_n359), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n391), .A2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(G190), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n357), .A2(new_n403), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n404), .B1(G200), .B2(new_n357), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n397), .A2(KEYINPUT17), .A3(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n383), .A2(new_n387), .A3(new_n405), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT17), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n406), .A2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n345), .A2(new_n402), .A3(new_n411), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n217), .A2(new_n214), .ZN(new_n413));
  OAI22_X1  g0213(.A1(new_n302), .A2(new_n202), .B1(new_n283), .B2(new_n306), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n288), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  XNOR2_X1  g0215(.A(new_n415), .B(KEYINPUT11), .ZN(new_n416));
  OAI21_X1  g0216(.A(KEYINPUT12), .B1(new_n217), .B2(new_n293), .ZN(new_n417));
  OAI21_X1  g0217(.A(G68), .B1(new_n299), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n417), .B1(KEYINPUT12), .B2(new_n293), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n416), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(G33), .A2(G97), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n250), .A2(new_n252), .A3(G226), .A4(new_n247), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n250), .A2(new_n252), .A3(G232), .A4(G1698), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n422), .B(new_n423), .C1(new_n424), .C2(KEYINPUT74), .ZN(new_n425));
  AND2_X1   g0225(.A1(new_n424), .A2(KEYINPUT74), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n259), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  NOR3_X1   g0228(.A1(new_n258), .A2(new_n262), .A3(new_n213), .ZN(new_n429));
  AOI21_X1  g0229(.A(KEYINPUT68), .B1(new_n264), .B2(new_n265), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT75), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n431), .A2(new_n432), .A3(G274), .A4(new_n269), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n431), .A2(G238), .A3(new_n273), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n270), .A2(KEYINPUT75), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  OAI21_X1  g0236(.A(KEYINPUT13), .B1(new_n428), .B2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  AOI22_X1  g0238(.A1(new_n274), .A2(G238), .B1(new_n270), .B2(KEYINPUT75), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT13), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n427), .A2(new_n439), .A3(new_n440), .A4(new_n433), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(G190), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n421), .B1(new_n438), .B2(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n427), .A2(new_n439), .A3(new_n433), .ZN(new_n444));
  AND3_X1   g0244(.A1(new_n444), .A2(KEYINPUT76), .A3(KEYINPUT13), .ZN(new_n445));
  AOI21_X1  g0245(.A(KEYINPUT76), .B1(new_n444), .B2(KEYINPUT13), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n441), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n443), .B1(new_n447), .B2(G200), .ZN(new_n448));
  INV_X1    g0248(.A(new_n441), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT76), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n437), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n444), .A2(KEYINPUT76), .A3(KEYINPUT13), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n449), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(KEYINPUT77), .A2(G169), .ZN(new_n454));
  OAI21_X1  g0254(.A(KEYINPUT14), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT14), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n447), .A2(KEYINPUT77), .A3(new_n456), .A4(G169), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT78), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n441), .A2(G179), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n458), .B1(new_n438), .B2(new_n459), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n437), .A2(KEYINPUT78), .A3(G179), .A4(new_n441), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n455), .A2(new_n457), .A3(new_n462), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n448), .B1(new_n463), .B2(new_n420), .ZN(new_n464));
  AND2_X1   g0264(.A1(new_n464), .A2(KEYINPUT79), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n464), .A2(KEYINPUT79), .ZN(new_n466));
  NOR3_X1   g0266(.A1(new_n412), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n249), .A2(G97), .ZN(new_n469));
  NAND2_X1  g0269(.A1(G33), .A2(G283), .ZN(new_n470));
  AOI21_X1  g0270(.A(G20), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(G116), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(KEYINPUT87), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT87), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(G116), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n214), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n288), .B1(new_n471), .B2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT20), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n288), .B(KEYINPUT20), .C1(new_n471), .C2(new_n476), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n272), .A2(G33), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n293), .A2(new_n482), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n288), .A2(new_n483), .ZN(new_n484));
  XNOR2_X1  g0284(.A(KEYINPUT87), .B(G116), .ZN(new_n485));
  AOI22_X1  g0285(.A1(new_n484), .A2(G116), .B1(new_n294), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n481), .A2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n272), .A2(G45), .ZN(new_n489));
  NOR2_X1   g0289(.A1(KEYINPUT5), .A2(G41), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(KEYINPUT5), .A2(G41), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n489), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n431), .A2(KEYINPUT85), .A3(G274), .A4(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT85), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n263), .A2(G274), .A3(new_n266), .ZN(new_n496));
  INV_X1    g0296(.A(new_n489), .ZN(new_n497));
  INV_X1    g0297(.A(new_n492), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n497), .B1(new_n498), .B2(new_n490), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n495), .B1(new_n496), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n263), .A2(new_n266), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n501), .A2(new_n493), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n494), .A2(new_n500), .B1(G270), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(G264), .A2(G1698), .ZN(new_n504));
  INV_X1    g0304(.A(G257), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n504), .B1(new_n505), .B2(G1698), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n506), .A2(new_n349), .A3(new_n351), .A4(new_n250), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n253), .A2(G303), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT89), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n507), .A2(new_n508), .A3(KEYINPUT89), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n511), .A2(new_n259), .A3(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n503), .A2(G179), .A3(new_n513), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n488), .A2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(G169), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n516), .B1(new_n481), .B2(new_n486), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n494), .A2(new_n500), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n502), .A2(G270), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n513), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n517), .A2(new_n520), .A3(KEYINPUT21), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(KEYINPUT90), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT90), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n517), .A2(new_n520), .A3(new_n523), .A4(KEYINPUT21), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n515), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n520), .A2(G200), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n526), .A2(KEYINPUT92), .A3(new_n488), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT92), .ZN(new_n528));
  INV_X1    g0328(.A(G200), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n529), .B1(new_n503), .B2(new_n513), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n528), .B1(new_n530), .B2(new_n487), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n503), .A2(G190), .A3(new_n513), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n527), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT21), .ZN(new_n534));
  AND3_X1   g0334(.A1(new_n517), .A2(KEYINPUT91), .A3(new_n520), .ZN(new_n535));
  AOI21_X1  g0335(.A(KEYINPUT91), .B1(new_n517), .B2(new_n520), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n525), .A2(new_n533), .A3(new_n537), .ZN(new_n538));
  AND2_X1   g0338(.A1(new_n287), .A2(new_n213), .ZN(new_n539));
  INV_X1    g0339(.A(new_n483), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n539), .A2(new_n540), .A3(KEYINPUT83), .A4(new_n285), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT83), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n542), .B1(new_n288), .B2(new_n483), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n541), .A2(new_n543), .A3(G97), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n293), .A2(G97), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT6), .ZN(new_n547));
  INV_X1    g0347(.A(G97), .ZN(new_n548));
  INV_X1    g0348(.A(G107), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NOR2_X1   g0350(.A1(G97), .A2(G107), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n547), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n549), .A2(KEYINPUT6), .A3(G97), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n554), .A2(G20), .B1(G77), .B2(new_n280), .ZN(new_n555));
  INV_X1    g0355(.A(new_n315), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n556), .B1(new_n362), .B2(new_n363), .ZN(new_n557));
  AND2_X1   g0357(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n544), .B(new_n546), .C1(new_n558), .C2(new_n290), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n349), .A2(new_n351), .A3(G244), .A4(new_n250), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(KEYINPUT4), .B1(new_n561), .B2(new_n247), .ZN(new_n562));
  AND2_X1   g0362(.A1(KEYINPUT4), .A2(G244), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n250), .A2(new_n252), .A3(new_n563), .A4(new_n247), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT84), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n245), .A2(KEYINPUT84), .A3(new_n247), .A4(new_n563), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n245), .A2(G250), .A3(G1698), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n566), .A2(new_n567), .A3(new_n470), .A4(new_n568), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n259), .B1(new_n562), .B2(new_n569), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n494), .A2(new_n500), .B1(G257), .B2(new_n502), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n529), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n570), .A2(new_n571), .A3(new_n403), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n559), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n290), .B1(new_n555), .B2(new_n557), .ZN(new_n576));
  INV_X1    g0376(.A(new_n544), .ZN(new_n577));
  NOR3_X1   g0377(.A1(new_n576), .A2(new_n577), .A3(new_n545), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n572), .A2(G169), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n570), .A2(new_n571), .A3(G179), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n578), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n575), .A2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(G264), .ZN(new_n583));
  NOR3_X1   g0383(.A1(new_n501), .A2(new_n493), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(G257), .A2(G1698), .ZN(new_n585));
  INV_X1    g0385(.A(G250), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n585), .B1(new_n586), .B2(G1698), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n587), .A2(new_n349), .A3(new_n351), .A4(new_n250), .ZN(new_n588));
  NAND2_X1  g0388(.A1(G33), .A2(G294), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n348), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n584), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n518), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(G169), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT93), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n594), .B1(new_n584), .B2(new_n590), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n588), .A2(new_n589), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n259), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n431), .A2(G264), .A3(new_n499), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n597), .A2(new_n598), .A3(KEYINPUT93), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n595), .A2(new_n599), .A3(G179), .A4(new_n518), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT22), .ZN(new_n601));
  INV_X1    g0401(.A(G87), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n349), .A2(new_n603), .A3(new_n351), .A4(new_n250), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n473), .A2(new_n475), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(G33), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n214), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n313), .A2(G20), .A3(new_n314), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(KEYINPUT23), .ZN(new_n610));
  OR3_X1    g0410(.A1(new_n214), .A2(KEYINPUT23), .A3(G107), .ZN(new_n611));
  AND2_X1   g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n214), .A2(G87), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n601), .B1(new_n253), .B2(new_n613), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n608), .A2(new_n612), .A3(KEYINPUT24), .A4(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT24), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n614), .A2(new_n610), .A3(new_n611), .ZN(new_n617));
  AOI21_X1  g0417(.A(G20), .B1(new_n604), .B2(new_n606), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n615), .A2(new_n619), .A3(new_n288), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n541), .A2(new_n543), .A3(G107), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n293), .A2(G107), .ZN(new_n622));
  XNOR2_X1  g0422(.A(new_n622), .B(KEYINPUT25), .ZN(new_n623));
  AND2_X1   g0423(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n593), .A2(new_n600), .B1(new_n620), .B2(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n595), .A2(new_n599), .A3(new_n518), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  OAI22_X1  g0427(.A1(new_n627), .A2(G200), .B1(G190), .B2(new_n592), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n620), .A2(new_n624), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n625), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT19), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n313), .A2(new_n602), .A3(new_n548), .A4(new_n314), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n422), .A2(new_n214), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n632), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NOR3_X1   g0435(.A1(new_n422), .A2(KEYINPUT19), .A3(G20), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n214), .A2(G68), .ZN(new_n637));
  OAI22_X1  g0437(.A1(new_n635), .A2(new_n636), .B1(new_n372), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n288), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n303), .A2(new_n294), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n541), .A2(new_n543), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n639), .B(new_n640), .C1(new_n303), .C2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n497), .A2(G274), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n489), .A2(G250), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n501), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n606), .B1(new_n560), .B2(new_n247), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT86), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n219), .A2(G1698), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n352), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n349), .A2(new_n351), .A3(new_n250), .A4(new_n649), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(KEYINPUT86), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n647), .B1(new_n650), .B2(new_n652), .ZN(new_n653));
  OAI211_X1 g0453(.A(new_n278), .B(new_n646), .C1(new_n653), .C2(new_n348), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n650), .A2(new_n652), .ZN(new_n655));
  INV_X1    g0455(.A(new_n647), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n645), .B1(new_n657), .B2(new_n259), .ZN(new_n658));
  OAI211_X1 g0458(.A(new_n642), .B(new_n654), .C1(new_n658), .C2(G169), .ZN(new_n659));
  INV_X1    g0459(.A(new_n323), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n348), .B1(new_n655), .B2(new_n656), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n660), .B1(new_n661), .B2(new_n645), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n541), .A2(new_n543), .A3(G87), .ZN(new_n663));
  AND3_X1   g0463(.A1(new_n639), .A2(new_n640), .A3(new_n663), .ZN(new_n664));
  OAI211_X1 g0464(.A(G190), .B(new_n646), .C1(new_n653), .C2(new_n348), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n662), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT88), .ZN(new_n667));
  AND3_X1   g0467(.A1(new_n659), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n667), .B1(new_n659), .B2(new_n666), .ZN(new_n669));
  OAI211_X1 g0469(.A(new_n582), .B(new_n631), .C1(new_n668), .C2(new_n669), .ZN(new_n670));
  NOR3_X1   g0470(.A1(new_n468), .A2(new_n538), .A3(new_n670), .ZN(G372));
  INV_X1    g0471(.A(new_n442), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n420), .B1(new_n672), .B2(new_n437), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n673), .B1(new_n453), .B2(new_n529), .ZN(new_n674));
  AOI22_X1  g0474(.A1(new_n463), .A2(new_n420), .B1(new_n321), .B2(new_n674), .ZN(new_n675));
  AOI211_X1 g0475(.A(new_n399), .B(new_n359), .C1(new_n383), .C2(new_n387), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n383), .A2(new_n387), .ZN(new_n677));
  INV_X1    g0477(.A(new_n359), .ZN(new_n678));
  AOI21_X1  g0478(.A(KEYINPUT18), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  OAI22_X1  g0479(.A1(new_n675), .A2(new_n410), .B1(new_n676), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n342), .A2(new_n344), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n297), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n659), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n659), .A2(new_n666), .ZN(new_n684));
  INV_X1    g0484(.A(new_n580), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n516), .B1(new_n570), .B2(new_n571), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n559), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT26), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n683), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n684), .A2(KEYINPUT88), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n659), .A2(new_n666), .A3(new_n667), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n687), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n690), .B1(new_n693), .B2(new_n689), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n593), .A2(new_n600), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(new_n629), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT94), .ZN(new_n697));
  AND3_X1   g0497(.A1(new_n525), .A2(new_n697), .A3(new_n537), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n697), .B1(new_n525), .B2(new_n537), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n696), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  AND2_X1   g0500(.A1(new_n659), .A2(new_n666), .ZN(new_n701));
  INV_X1    g0501(.A(new_n592), .ZN(new_n702));
  AOI22_X1  g0502(.A1(new_n702), .A2(new_n403), .B1(new_n626), .B2(new_n529), .ZN(new_n703));
  OAI211_X1 g0503(.A(new_n582), .B(new_n701), .C1(new_n629), .C2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n694), .B1(new_n700), .B2(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n682), .B1(new_n468), .B2(new_n706), .ZN(G369));
  NAND3_X1  g0507(.A1(new_n272), .A2(new_n214), .A3(G13), .ZN(new_n708));
  OR2_X1    g0508(.A1(new_n708), .A2(KEYINPUT27), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(KEYINPUT27), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n709), .A2(G213), .A3(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT95), .ZN(new_n713));
  OR2_X1    g0513(.A1(new_n713), .A2(G343), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(G343), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n712), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n631), .B1(new_n630), .B2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n717), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n695), .A2(new_n629), .A3(new_n719), .ZN(new_n720));
  OR2_X1    g0520(.A1(new_n720), .A2(KEYINPUT96), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(KEYINPUT96), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n718), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n719), .B1(new_n525), .B2(new_n537), .ZN(new_n724));
  AOI22_X1  g0524(.A1(new_n723), .A2(new_n724), .B1(new_n625), .B2(new_n717), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n525), .A2(new_n537), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(KEYINPUT94), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n525), .A2(new_n697), .A3(new_n537), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n729), .A2(new_n487), .A3(new_n719), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n538), .B1(new_n488), .B2(new_n717), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n730), .A2(G330), .A3(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n723), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n725), .B1(new_n732), .B2(new_n733), .ZN(G399));
  INV_X1    g0534(.A(new_n208), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(G41), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n633), .A2(G116), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n737), .A2(G1), .A3(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n739), .B1(new_n211), .B2(new_n737), .ZN(new_n740));
  XNOR2_X1  g0540(.A(new_n740), .B(KEYINPUT28), .ZN(new_n741));
  INV_X1    g0541(.A(G330), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT31), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n646), .B1(new_n653), .B2(new_n348), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n572), .A2(new_n744), .A3(new_n520), .A4(new_n278), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(new_n627), .ZN(new_n746));
  NOR2_X1   g0546(.A1(KEYINPUT98), .A2(KEYINPUT30), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  AND2_X1   g0548(.A1(new_n595), .A2(new_n599), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n749), .A2(new_n658), .A3(new_n570), .A4(new_n571), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n748), .B1(new_n750), .B2(new_n514), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n570), .A2(new_n571), .A3(new_n595), .A4(new_n599), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(new_n744), .ZN(new_n753));
  INV_X1    g0553(.A(new_n514), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n753), .A2(new_n754), .A3(new_n747), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n746), .B1(new_n751), .B2(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n743), .B1(new_n756), .B2(new_n717), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n747), .B1(new_n753), .B2(new_n754), .ZN(new_n758));
  NOR4_X1   g0558(.A1(new_n752), .A2(new_n514), .A3(new_n744), .A4(new_n748), .ZN(new_n759));
  OAI22_X1  g0559(.A1(new_n758), .A2(new_n759), .B1(new_n627), .B2(new_n745), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(new_n719), .ZN(new_n761));
  XNOR2_X1  g0561(.A(KEYINPUT97), .B(KEYINPUT31), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n757), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  AND3_X1   g0564(.A1(new_n525), .A2(new_n533), .A3(new_n537), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n691), .A2(new_n692), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n696), .B1(new_n629), .B2(new_n703), .ZN(new_n767));
  INV_X1    g0567(.A(new_n574), .ZN(new_n768));
  AOI21_X1  g0568(.A(G200), .B1(new_n570), .B2(new_n571), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n578), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(new_n687), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n767), .A2(new_n771), .ZN(new_n772));
  NAND4_X1  g0572(.A1(new_n765), .A2(new_n766), .A3(new_n772), .A4(new_n717), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n742), .B1(new_n764), .B2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(KEYINPUT29), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n775), .B1(new_n706), .B2(new_n719), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n766), .A2(new_n689), .A3(new_n581), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n701), .A2(new_n581), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n683), .B1(new_n778), .B2(KEYINPUT26), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n726), .A2(new_n625), .ZN(new_n780));
  OAI211_X1 g0580(.A(new_n777), .B(new_n779), .C1(new_n704), .C2(new_n780), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n781), .A2(KEYINPUT29), .A3(new_n717), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n774), .B1(new_n776), .B2(new_n782), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n741), .B1(new_n783), .B2(G1), .ZN(G364));
  AND2_X1   g0584(.A1(new_n214), .A2(G13), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(G45), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n737), .A2(G1), .A3(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n214), .A2(G190), .ZN(new_n788));
  NOR2_X1   g0588(.A1(G179), .A2(G200), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  OR2_X1    g0591(.A1(new_n791), .A2(KEYINPUT102), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n791), .A2(KEYINPUT102), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n660), .A2(new_n278), .A3(new_n788), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n795), .A2(G329), .B1(G283), .B2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(G303), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n214), .A2(new_n403), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n660), .A2(new_n278), .A3(new_n800), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n798), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n278), .A2(new_n529), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(new_n788), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(KEYINPUT33), .A2(G317), .ZN(new_n806));
  AND2_X1   g0606(.A1(KEYINPUT33), .A2(G317), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n805), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(G311), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n278), .A2(G200), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n788), .A2(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n808), .B1(new_n809), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n803), .A2(new_n800), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n812), .B1(G326), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n800), .A2(new_n810), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n245), .B1(new_n817), .B2(G322), .ZN(new_n818));
  INV_X1    g0618(.A(G294), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n789), .A2(G190), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(G20), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  OAI211_X1 g0622(.A(new_n815), .B(new_n818), .C1(new_n819), .C2(new_n822), .ZN(new_n823));
  AOI22_X1  g0623(.A1(G50), .A2(new_n814), .B1(new_n817), .B2(G58), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n805), .A2(G68), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n821), .A2(G97), .ZN(new_n826));
  INV_X1    g0626(.A(new_n811), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n253), .B1(new_n827), .B2(G77), .ZN(new_n828));
  NAND4_X1  g0628(.A1(new_n824), .A2(new_n825), .A3(new_n826), .A4(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n797), .A2(G107), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n790), .A2(new_n366), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(KEYINPUT32), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n830), .B(new_n832), .C1(new_n602), .C2(new_n801), .ZN(new_n833));
  OAI22_X1  g0633(.A1(new_n802), .A2(new_n823), .B1(new_n829), .B2(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n213), .B1(G20), .B2(new_n516), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n787), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n735), .A2(new_n253), .ZN(new_n837));
  AOI22_X1  g0637(.A1(G355), .A2(new_n837), .B1(new_n472), .B2(new_n735), .ZN(new_n838));
  XNOR2_X1  g0638(.A(new_n838), .B(KEYINPUT100), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n352), .A2(new_n735), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n243), .A2(new_n268), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n212), .A2(G45), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n840), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(KEYINPUT101), .B1(new_n839), .B2(new_n843), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n839), .A2(KEYINPUT101), .A3(new_n843), .ZN(new_n845));
  NOR2_X1   g0645(.A1(G13), .A2(G33), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n847), .A2(G20), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n848), .A2(new_n835), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n845), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n730), .A2(new_n731), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n848), .ZN(new_n853));
  OAI221_X1 g0653(.A(new_n836), .B1(new_n844), .B2(new_n850), .C1(new_n852), .C2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n787), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n852), .A2(G330), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT99), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n855), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n856), .B1(new_n857), .B2(new_n732), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n854), .B1(new_n859), .B2(new_n860), .ZN(G396));
  NOR2_X1   g0661(.A1(new_n835), .A2(new_n846), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n787), .B1(new_n306), .B2(new_n862), .ZN(new_n863));
  XNOR2_X1  g0663(.A(new_n863), .B(KEYINPUT103), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n797), .A2(G87), .ZN(new_n865));
  OAI221_X1 g0665(.A(new_n865), .B1(new_n549), .B2(new_n801), .C1(new_n809), .C2(new_n794), .ZN(new_n866));
  AOI22_X1  g0666(.A1(G283), .A2(new_n805), .B1(new_n827), .B2(new_n605), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n867), .B1(new_n819), .B2(new_n816), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n826), .B(new_n253), .C1(new_n799), .C2(new_n813), .ZN(new_n869));
  NOR3_X1   g0669(.A1(new_n866), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n796), .A2(new_n379), .ZN(new_n871));
  INV_X1    g0671(.A(new_n801), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n871), .B1(G50), .B2(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n372), .B1(G58), .B2(new_n821), .ZN(new_n874));
  INV_X1    g0674(.A(G132), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n873), .B(new_n874), .C1(new_n875), .C2(new_n794), .ZN(new_n876));
  XOR2_X1   g0676(.A(new_n876), .B(KEYINPUT104), .Z(new_n877));
  AOI22_X1  g0677(.A1(new_n814), .A2(G137), .B1(new_n827), .B2(G159), .ZN(new_n878));
  INV_X1    g0678(.A(G143), .ZN(new_n879));
  INV_X1    g0679(.A(G150), .ZN(new_n880));
  OAI221_X1 g0680(.A(new_n878), .B1(new_n879), .B2(new_n816), .C1(new_n880), .C2(new_n804), .ZN(new_n881));
  XNOR2_X1  g0681(.A(new_n881), .B(KEYINPUT34), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n870), .B1(new_n877), .B2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n835), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n322), .A2(new_n719), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n326), .B1(new_n309), .B2(new_n717), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(new_n322), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  OAI221_X1 g0690(.A(new_n864), .B1(new_n883), .B2(new_n884), .C1(new_n890), .C2(new_n847), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n700), .A2(new_n705), .ZN(new_n892));
  INV_X1    g0692(.A(new_n694), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n719), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n894), .B(new_n889), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(new_n774), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n787), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n895), .A2(new_n774), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n891), .B1(new_n897), .B2(new_n898), .ZN(G384));
  OAI211_X1 g0699(.A(G116), .B(new_n215), .C1(new_n554), .C2(KEYINPUT35), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n900), .B1(KEYINPUT35), .B2(new_n554), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n901), .B(KEYINPUT36), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n217), .A2(G58), .ZN(new_n903));
  INV_X1    g0703(.A(new_n211), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n903), .A2(G77), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n202), .A2(G68), .ZN(new_n906));
  AOI211_X1 g0706(.A(new_n272), .B(G13), .C1(new_n905), .C2(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n902), .A2(new_n907), .ZN(new_n908));
  NOR3_X1   g0708(.A1(new_n756), .A2(KEYINPUT31), .A3(new_n717), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  NOR3_X1   g0710(.A1(new_n670), .A2(new_n538), .A3(new_n719), .ZN(new_n911));
  INV_X1    g0711(.A(new_n762), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n761), .A2(new_n912), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n890), .B(new_n910), .C1(new_n911), .C2(new_n913), .ZN(new_n914));
  NAND4_X1  g0714(.A1(new_n455), .A2(new_n674), .A3(new_n457), .A4(new_n462), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n421), .A2(new_n717), .ZN(new_n916));
  AND2_X1   g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AOI211_X1 g0717(.A(new_n448), .B(new_n916), .C1(new_n463), .C2(new_n420), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT105), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n917), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n916), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n464), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(KEYINPUT105), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n914), .B1(new_n920), .B2(new_n923), .ZN(new_n924));
  OR2_X1    g0724(.A1(new_n381), .A2(KEYINPUT16), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n386), .B1(new_n396), .B2(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n926), .A2(new_n711), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n928), .B1(new_n402), .B2(new_n411), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n677), .B1(new_n678), .B2(new_n712), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n407), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n931), .A2(KEYINPUT37), .ZN(new_n932));
  AND3_X1   g0732(.A1(new_n383), .A2(new_n387), .A3(new_n405), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n288), .B(new_n925), .C1(new_n378), .C2(new_n382), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n359), .B1(new_n934), .B2(new_n387), .ZN(new_n935));
  OAI21_X1  g0735(.A(KEYINPUT106), .B1(new_n933), .B2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT106), .ZN(new_n937));
  OAI211_X1 g0737(.A(new_n407), .B(new_n937), .C1(new_n926), .C2(new_n359), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n936), .A2(new_n938), .A3(new_n928), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n932), .B1(KEYINPUT37), .B2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT38), .ZN(new_n941));
  NOR3_X1   g0741(.A1(new_n929), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n939), .A2(KEYINPUT37), .ZN(new_n943));
  INV_X1    g0743(.A(new_n932), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n400), .B1(new_n390), .B2(new_n389), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n927), .B1(new_n946), .B2(new_n410), .ZN(new_n947));
  AOI21_X1  g0747(.A(KEYINPUT38), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n924), .B1(new_n942), .B2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT40), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n945), .A2(new_n947), .A3(KEYINPUT38), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n397), .A2(new_n711), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n679), .A2(new_n676), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n952), .B1(new_n953), .B2(new_n410), .ZN(new_n954));
  AOI22_X1  g0754(.A1(new_n383), .A2(new_n387), .B1(new_n359), .B2(new_n711), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT107), .ZN(new_n956));
  OAI21_X1  g0756(.A(KEYINPUT37), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n931), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n931), .A2(new_n957), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n954), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(new_n941), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n950), .B1(new_n951), .B2(new_n961), .ZN(new_n962));
  AOI22_X1  g0762(.A1(new_n949), .A2(new_n950), .B1(new_n924), .B2(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n762), .B1(new_n760), .B2(new_n719), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n909), .B1(new_n773), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n467), .A2(new_n965), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n963), .B(new_n966), .Z(new_n967));
  NOR2_X1   g0767(.A1(new_n967), .A2(new_n742), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n463), .A2(new_n420), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n969), .A2(new_n719), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(KEYINPUT39), .B1(new_n942), .B2(new_n948), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT39), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n951), .A2(new_n973), .A3(new_n961), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n971), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n941), .B1(new_n929), .B2(new_n940), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n951), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n704), .B1(new_n729), .B2(new_n696), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n717), .B1(new_n978), .B2(new_n694), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n886), .B1(new_n979), .B2(new_n889), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n920), .A2(new_n923), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n977), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n953), .A2(new_n711), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n975), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n467), .A2(new_n776), .A3(new_n782), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(new_n682), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n985), .B(new_n987), .ZN(new_n988));
  OAI22_X1  g0788(.A1(new_n968), .A2(new_n988), .B1(new_n272), .B2(new_n785), .ZN(new_n989));
  AND2_X1   g0789(.A1(new_n968), .A2(new_n988), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n908), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n991), .B(KEYINPUT108), .Z(G367));
  NAND2_X1  g0792(.A1(new_n723), .A2(new_n724), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n582), .B1(new_n578), .B2(new_n717), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n687), .B2(new_n717), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  AND2_X1   g0797(.A1(new_n997), .A2(KEYINPUT42), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n687), .B1(new_n995), .B2(new_n696), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n999), .A2(new_n717), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(new_n997), .B2(KEYINPUT42), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT43), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n664), .A2(new_n717), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n659), .A2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(new_n701), .B2(new_n1003), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n998), .A2(new_n1001), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(new_n1002), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1006), .B(new_n1007), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n732), .A2(new_n733), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(new_n996), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1008), .B(new_n1010), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n736), .B(KEYINPUT41), .Z(new_n1012));
  XNOR2_X1  g0812(.A(new_n732), .B(new_n733), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n724), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n994), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  OR3_X1    g0815(.A1(new_n725), .A2(KEYINPUT44), .A3(new_n996), .ZN(new_n1016));
  OAI21_X1  g0816(.A(KEYINPUT44), .B1(new_n725), .B2(new_n996), .ZN(new_n1017));
  AND3_X1   g0817(.A1(new_n725), .A2(KEYINPUT45), .A3(new_n996), .ZN(new_n1018));
  AOI21_X1  g0818(.A(KEYINPUT45), .B1(new_n725), .B2(new_n996), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n1016), .B(new_n1017), .C1(new_n1018), .C2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1015), .A2(new_n783), .A3(new_n1020), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT109), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1012), .B1(new_n1022), .B2(new_n783), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n786), .A2(G1), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1011), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n814), .A2(G311), .B1(new_n805), .B2(G294), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n1026), .B(new_n372), .C1(new_n315), .C2(new_n822), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n797), .A2(G97), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(G303), .A2(new_n817), .B1(new_n791), .B2(G317), .ZN(new_n1029));
  INV_X1    g0829(.A(G283), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n1028), .B(new_n1029), .C1(new_n1030), .C2(new_n811), .ZN(new_n1031));
  OAI21_X1  g0831(.A(KEYINPUT46), .B1(new_n801), .B2(new_n472), .ZN(new_n1032));
  OR3_X1    g0832(.A1(new_n801), .A2(KEYINPUT46), .A3(new_n485), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n1027), .B(new_n1031), .C1(new_n1032), .C2(new_n1033), .ZN(new_n1034));
  AND2_X1   g0834(.A1(new_n1034), .A2(KEYINPUT110), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n1034), .A2(KEYINPUT110), .ZN(new_n1036));
  INV_X1    g0836(.A(G137), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n245), .B1(new_n790), .B2(new_n1037), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n804), .A2(new_n366), .B1(new_n811), .B2(new_n202), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n1038), .B(new_n1039), .C1(G143), .C2(new_n814), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n821), .A2(G68), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1041), .B1(new_n880), .B2(new_n816), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT111), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n872), .A2(G58), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n797), .A2(G77), .ZN(new_n1045));
  AND4_X1   g0845(.A1(new_n1040), .A2(new_n1043), .A3(new_n1044), .A4(new_n1045), .ZN(new_n1046));
  NOR3_X1   g0846(.A1(new_n1035), .A2(new_n1036), .A3(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n884), .B1(new_n1047), .B2(KEYINPUT47), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1048), .B1(KEYINPUT47), .B2(new_n1047), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1005), .A2(new_n848), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n840), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n849), .B1(new_n208), .B2(new_n303), .C1(new_n1051), .C2(new_n235), .ZN(new_n1052));
  NAND4_X1  g0852(.A1(new_n1049), .A2(new_n1050), .A3(new_n855), .A4(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1025), .A2(new_n1053), .ZN(G387));
  AOI21_X1  g0854(.A(new_n737), .B1(new_n1015), .B2(new_n783), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1055), .B1(new_n783), .B2(new_n1015), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n733), .A2(new_n848), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n837), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n1058), .A2(new_n738), .B1(G107), .B2(new_n208), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n232), .A2(G45), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n738), .ZN(new_n1061));
  AOI211_X1 g0861(.A(G45), .B(new_n1061), .C1(G68), .C2(G77), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n282), .A2(G50), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT50), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1051), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1059), .B1(new_n1060), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT112), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n849), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(new_n1067), .B2(new_n1066), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n872), .A2(G77), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n827), .A2(G68), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(G50), .A2(new_n817), .B1(new_n805), .B2(new_n384), .ZN(new_n1072));
  NAND4_X1  g0872(.A1(new_n1028), .A2(new_n1070), .A3(new_n1071), .A4(new_n1072), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n822), .A2(new_n303), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n813), .A2(new_n366), .B1(new_n790), .B2(new_n880), .ZN(new_n1075));
  OR4_X1    g0875(.A1(new_n372), .A2(new_n1073), .A3(new_n1074), .A4(new_n1075), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n872), .A2(G294), .B1(G283), .B2(new_n821), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n814), .A2(G322), .B1(new_n827), .B2(G303), .ZN(new_n1078));
  INV_X1    g0878(.A(G317), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n1078), .B1(new_n809), .B2(new_n804), .C1(new_n1079), .C2(new_n816), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT48), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1077), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(new_n1081), .B2(new_n1080), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(KEYINPUT113), .B(KEYINPUT49), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(new_n1083), .B(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n352), .B1(G326), .B2(new_n791), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1086), .B1(new_n485), .B2(new_n796), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1076), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n787), .B(new_n1069), .C1(new_n1088), .C2(new_n835), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n1015), .A2(new_n1024), .B1(new_n1057), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1056), .A2(new_n1090), .ZN(G393));
  INV_X1    g0891(.A(KEYINPUT114), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1092), .B1(new_n1020), .B2(new_n1009), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1020), .A2(new_n1009), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n1095), .B(new_n1024), .C1(KEYINPUT114), .C2(new_n1094), .ZN(new_n1096));
  OR2_X1    g0896(.A1(new_n240), .A2(new_n1051), .ZN(new_n1097));
  AOI211_X1 g0897(.A(new_n835), .B(new_n848), .C1(G97), .C2(new_n735), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n787), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(G303), .A2(new_n805), .B1(new_n791), .B2(G322), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1100), .B(new_n253), .C1(new_n819), .C2(new_n811), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n813), .A2(new_n1079), .B1(new_n816), .B2(new_n809), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT52), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1103), .B(new_n830), .C1(new_n1030), .C2(new_n801), .ZN(new_n1104));
  AOI211_X1 g0904(.A(new_n1101), .B(new_n1104), .C1(new_n605), .C2(new_n821), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(new_n1105), .B(KEYINPUT116), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n372), .B1(new_n791), .B2(G143), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n865), .B(new_n1107), .C1(new_n218), .C2(new_n801), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1108), .B(KEYINPUT115), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n813), .A2(new_n880), .B1(new_n816), .B2(new_n366), .ZN(new_n1110));
  XOR2_X1   g0910(.A(new_n1110), .B(KEYINPUT51), .Z(new_n1111));
  NOR2_X1   g0911(.A1(new_n822), .A2(new_n306), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n804), .A2(new_n202), .B1(new_n811), .B2(new_n282), .ZN(new_n1113));
  NOR3_X1   g0913(.A1(new_n1111), .A2(new_n1112), .A3(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1106), .B1(new_n1109), .B2(new_n1114), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n1099), .B1(new_n996), .B2(new_n853), .C1(new_n1115), .C2(new_n884), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1096), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT117), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(new_n1117), .B(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1015), .A2(new_n783), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1095), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1094), .A2(KEYINPUT114), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1120), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(KEYINPUT118), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  OAI211_X1 g0925(.A(KEYINPUT118), .B(new_n1120), .C1(new_n1121), .C2(new_n1122), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1125), .A2(new_n1126), .A3(new_n736), .A4(new_n1022), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1119), .A2(new_n1127), .ZN(G390));
  INV_X1    g0928(.A(G128), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n813), .A2(new_n1129), .B1(new_n804), .B2(new_n1037), .ZN(new_n1130));
  OAI221_X1 g0930(.A(new_n245), .B1(new_n816), .B2(new_n875), .C1(new_n822), .C2(new_n366), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(KEYINPUT54), .B(G143), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  AOI211_X1 g0933(.A(new_n1130), .B(new_n1131), .C1(new_n827), .C2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n801), .A2(new_n880), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1135), .B(KEYINPUT53), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n795), .A2(G125), .B1(G50), .B2(new_n797), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1134), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n814), .A2(G283), .B1(new_n827), .B2(G97), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1139), .B1(new_n315), .B2(new_n804), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(new_n1140), .B(KEYINPUT120), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n245), .B1(new_n872), .B2(G87), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1141), .B1(KEYINPUT121), .B2(new_n1143), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n1112), .B(new_n871), .C1(G116), .C2(new_n817), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1143), .A2(KEYINPUT121), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n1145), .B(new_n1146), .C1(new_n819), .C2(new_n794), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1138), .B1(new_n1144), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT122), .ZN(new_n1149));
  OR2_X1    g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1150), .A2(new_n835), .A3(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n862), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1152), .B(new_n855), .C1(new_n384), .C2(new_n1153), .ZN(new_n1154));
  XOR2_X1   g0954(.A(new_n1154), .B(KEYINPUT123), .Z(new_n1155));
  INV_X1    g0955(.A(new_n974), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n973), .B1(new_n976), .B2(new_n951), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1155), .B1(new_n1159), .B2(new_n847), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n885), .B1(new_n894), .B2(new_n890), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n969), .A2(new_n919), .A3(new_n674), .A4(new_n921), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n915), .A2(new_n916), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n919), .B1(new_n464), .B2(new_n921), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n971), .B1(new_n1161), .B2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1167), .A2(new_n972), .A3(new_n974), .ZN(new_n1168));
  OAI21_X1  g0968(.A(KEYINPUT119), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT119), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n923), .A2(new_n1170), .A3(new_n1162), .A4(new_n1163), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1169), .A2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n781), .A2(new_n717), .A3(new_n888), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(new_n886), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n970), .B1(new_n951), .B2(new_n961), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  OAI211_X1 g0977(.A(G330), .B(new_n890), .C1(new_n763), .C2(new_n911), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n981), .A2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1168), .A2(new_n1177), .A3(new_n1180), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n1158), .A2(new_n1167), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n889), .B(new_n909), .C1(new_n773), .C2(new_n964), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n981), .A2(G330), .A3(new_n1183), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1181), .B1(new_n1182), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1024), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1160), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n467), .A2(G330), .A3(new_n965), .ZN(new_n1188));
  AND3_X1   g0988(.A1(new_n986), .A2(new_n1188), .A3(new_n682), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1174), .B1(new_n981), .B2(new_n1179), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1183), .A2(G330), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1169), .A2(new_n1171), .A3(new_n1191), .ZN(new_n1192));
  AND2_X1   g0992(.A1(new_n1190), .A2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1166), .A2(new_n1178), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1161), .B1(new_n1184), .B2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1189), .B1(new_n1193), .B2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n737), .B1(new_n1185), .B2(new_n1196), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n986), .A2(new_n1188), .A3(new_n682), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1184), .A2(new_n1194), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1199), .A2(new_n980), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1190), .A2(new_n1192), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1198), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n1202), .B(new_n1181), .C1(new_n1182), .C2(new_n1184), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1187), .B1(new_n1197), .B2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(G378));
  OR2_X1    g1005(.A1(new_n975), .A2(new_n984), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n949), .A2(new_n950), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n951), .A2(new_n961), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1208), .A2(KEYINPUT40), .A3(new_n924), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n297), .B1(new_n342), .B2(new_n344), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n296), .A2(new_n712), .ZN(new_n1211));
  XOR2_X1   g1011(.A(new_n1210), .B(new_n1211), .Z(new_n1212));
  XNOR2_X1  g1012(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(new_n1212), .B(new_n1213), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1207), .A2(G330), .A3(new_n1209), .A4(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1214), .B1(new_n963), .B2(G330), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1206), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1183), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(new_n951), .B2(new_n976), .ZN(new_n1220));
  OAI211_X1 g1020(.A(G330), .B(new_n1209), .C1(new_n1220), .C2(KEYINPUT40), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1214), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1223), .A2(new_n985), .A3(new_n1215), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1218), .A2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT57), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1203), .A2(new_n1189), .ZN(new_n1227));
  AND3_X1   g1027(.A1(new_n1225), .A2(new_n1226), .A3(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1226), .B1(new_n1225), .B2(new_n1227), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n736), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n372), .A2(new_n267), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n797), .A2(G58), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  AOI211_X1 g1033(.A(new_n1231), .B(new_n1233), .C1(G283), .C2(new_n795), .ZN(new_n1234));
  OAI22_X1  g1034(.A1(new_n804), .A2(new_n548), .B1(new_n811), .B2(new_n303), .ZN(new_n1235));
  XOR2_X1   g1035(.A(new_n1235), .B(KEYINPUT124), .Z(new_n1236));
  OAI221_X1 g1036(.A(new_n1041), .B1(new_n549), .B2(new_n816), .C1(new_n472), .C2(new_n813), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(G77), .B2(new_n872), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1234), .A2(new_n1236), .A3(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT58), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1231), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1242));
  AND2_X1   g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n816), .A2(new_n1129), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n804), .A2(new_n875), .B1(new_n811), .B2(new_n1037), .ZN(new_n1245));
  AOI211_X1 g1045(.A(new_n1244), .B(new_n1245), .C1(G125), .C2(new_n814), .ZN(new_n1246));
  OAI221_X1 g1046(.A(new_n1246), .B1(new_n880), .B2(new_n822), .C1(new_n801), .C2(new_n1132), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1247), .A2(KEYINPUT59), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1247), .A2(KEYINPUT59), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n797), .A2(G159), .ZN(new_n1250));
  AOI211_X1 g1050(.A(G33), .B(G41), .C1(new_n791), .C2(G124), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1249), .A2(new_n1250), .A3(new_n1251), .ZN(new_n1252));
  OAI221_X1 g1052(.A(new_n1243), .B1(new_n1240), .B2(new_n1239), .C1(new_n1248), .C2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(new_n835), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n787), .B1(new_n202), .B2(new_n862), .ZN(new_n1255));
  OAI211_X1 g1055(.A(new_n1254), .B(new_n1255), .C1(new_n1214), .C2(new_n847), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1257), .B1(new_n1225), .B2(new_n1024), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1230), .A2(new_n1258), .ZN(G375));
  NOR2_X1   g1059(.A1(new_n1193), .A2(new_n1195), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1169), .A2(new_n1171), .A3(new_n846), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n855), .B1(G68), .B2(new_n1153), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n253), .B1(new_n813), .B2(new_n819), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1074), .A2(new_n1264), .ZN(new_n1265));
  AOI22_X1  g1065(.A1(new_n556), .A2(new_n827), .B1(new_n805), .B2(new_n605), .ZN(new_n1266));
  OAI211_X1 g1066(.A(new_n1265), .B(new_n1266), .C1(new_n1030), .C2(new_n816), .ZN(new_n1267));
  OAI221_X1 g1067(.A(new_n1045), .B1(new_n548), .B2(new_n801), .C1(new_n799), .C2(new_n794), .ZN(new_n1268));
  OAI221_X1 g1068(.A(new_n1232), .B1(new_n366), .B2(new_n801), .C1(new_n1129), .C2(new_n794), .ZN(new_n1269));
  AOI22_X1  g1069(.A1(G132), .A2(new_n814), .B1(new_n817), .B2(G137), .ZN(new_n1270));
  AOI22_X1  g1070(.A1(new_n805), .A2(new_n1133), .B1(new_n827), .B2(G150), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n372), .B1(G50), .B2(new_n821), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1270), .A2(new_n1271), .A3(new_n1272), .ZN(new_n1273));
  OAI22_X1  g1073(.A1(new_n1267), .A2(new_n1268), .B1(new_n1269), .B2(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1263), .B1(new_n1274), .B2(new_n835), .ZN(new_n1275));
  AOI22_X1  g1075(.A1(new_n1261), .A2(new_n1024), .B1(new_n1262), .B2(new_n1275), .ZN(new_n1276));
  OR2_X1    g1076(.A1(new_n1202), .A2(new_n1012), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1260), .A2(new_n1198), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1276), .B1(new_n1277), .B2(new_n1279), .ZN(G381));
  NOR2_X1   g1080(.A1(G375), .A2(G378), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1025), .A2(new_n1119), .A3(new_n1127), .A4(new_n1053), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  OR2_X1    g1083(.A1(G393), .A2(G396), .ZN(new_n1284));
  NOR3_X1   g1084(.A1(new_n1284), .A2(G381), .A3(G384), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1281), .A2(new_n1283), .A3(new_n1285), .ZN(G407));
  INV_X1    g1086(.A(new_n1281), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n714), .A2(new_n715), .A3(G213), .ZN(new_n1288));
  OAI211_X1 g1088(.A(G407), .B(G213), .C1(new_n1287), .C2(new_n1288), .ZN(G409));
  INV_X1    g1089(.A(KEYINPUT127), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(G387), .A2(G390), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(new_n1282), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(G393), .A2(G396), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1284), .A2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1292), .A2(new_n1295), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1291), .A2(new_n1282), .A3(new_n1294), .ZN(new_n1297));
  AND2_X1   g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT126), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT62), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1230), .A2(G378), .A3(new_n1258), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1258), .ZN(new_n1303));
  AND3_X1   g1103(.A1(new_n1168), .A2(new_n1177), .A3(new_n1180), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1184), .B1(new_n1168), .B2(new_n1177), .ZN(new_n1305));
  NOR3_X1   g1105(.A1(new_n1304), .A2(new_n1305), .A3(new_n1196), .ZN(new_n1306));
  AND3_X1   g1106(.A1(new_n1223), .A2(new_n985), .A3(new_n1215), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n985), .B1(new_n1223), .B2(new_n1215), .ZN(new_n1308));
  OAI22_X1  g1108(.A1(new_n1306), .A2(new_n1198), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n1309), .A2(new_n1012), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1204), .B1(new_n1303), .B2(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1302), .A2(new_n1311), .ZN(new_n1312));
  XNOR2_X1  g1112(.A(new_n1278), .B(KEYINPUT60), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1313), .A2(new_n736), .A3(new_n1196), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1314), .A2(G384), .A3(new_n1276), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1315), .ZN(new_n1316));
  AOI21_X1  g1116(.A(G384), .B1(new_n1314), .B2(new_n1276), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  NOR2_X1   g1118(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1319), .ZN(new_n1320));
  AND4_X1   g1120(.A1(new_n1288), .A2(new_n1312), .A3(new_n1318), .A4(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1288), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1322), .B1(new_n1302), .B2(new_n1311), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1320), .B1(new_n1323), .B2(new_n1318), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1301), .B1(new_n1321), .B2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1312), .A2(new_n1288), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1317), .ZN(new_n1327));
  NAND4_X1  g1127(.A1(new_n1327), .A2(G2897), .A3(new_n1322), .A4(new_n1315), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1322), .A2(G2897), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1329), .B1(new_n1316), .B2(new_n1317), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1328), .A2(new_n1330), .ZN(new_n1331));
  AOI21_X1  g1131(.A(KEYINPUT61), .B1(new_n1326), .B2(new_n1331), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1298), .B1(new_n1325), .B2(new_n1332), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT61), .ZN(new_n1334));
  AND3_X1   g1134(.A1(new_n1296), .A2(new_n1334), .A3(new_n1297), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1309), .A2(KEYINPUT57), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1225), .A2(new_n1226), .A3(new_n1227), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n737), .B1(new_n1336), .B2(new_n1337), .ZN(new_n1338));
  NOR3_X1   g1138(.A1(new_n1338), .A2(new_n1204), .A3(new_n1303), .ZN(new_n1339));
  INV_X1    g1139(.A(new_n1311), .ZN(new_n1340));
  OAI211_X1 g1140(.A(KEYINPUT125), .B(new_n1288), .C1(new_n1339), .C2(new_n1340), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1341), .A2(new_n1331), .ZN(new_n1342));
  NOR2_X1   g1142(.A1(new_n1323), .A2(KEYINPUT125), .ZN(new_n1343));
  OAI21_X1  g1143(.A(new_n1335), .B1(new_n1342), .B2(new_n1343), .ZN(new_n1344));
  INV_X1    g1144(.A(KEYINPUT63), .ZN(new_n1345));
  AND3_X1   g1145(.A1(new_n1323), .A2(new_n1345), .A3(new_n1318), .ZN(new_n1346));
  AOI21_X1  g1146(.A(new_n1345), .B1(new_n1323), .B2(new_n1318), .ZN(new_n1347));
  NOR2_X1   g1147(.A1(new_n1346), .A2(new_n1347), .ZN(new_n1348));
  NOR2_X1   g1148(.A1(new_n1344), .A2(new_n1348), .ZN(new_n1349));
  OAI21_X1  g1149(.A(new_n1290), .B1(new_n1333), .B2(new_n1349), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1312), .A2(new_n1288), .A3(new_n1318), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1351), .A2(KEYINPUT63), .ZN(new_n1352));
  NAND3_X1  g1152(.A1(new_n1323), .A2(new_n1345), .A3(new_n1318), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1352), .A2(new_n1353), .ZN(new_n1354));
  INV_X1    g1154(.A(KEYINPUT125), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1326), .A2(new_n1355), .ZN(new_n1356));
  NAND3_X1  g1156(.A1(new_n1356), .A2(new_n1331), .A3(new_n1341), .ZN(new_n1357));
  NAND3_X1  g1157(.A1(new_n1354), .A2(new_n1357), .A3(new_n1335), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1326), .A2(new_n1331), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1359), .A2(new_n1334), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1351), .A2(new_n1319), .ZN(new_n1361));
  NAND3_X1  g1161(.A1(new_n1323), .A2(new_n1318), .A3(new_n1320), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1361), .A2(new_n1362), .ZN(new_n1363));
  AOI21_X1  g1163(.A(new_n1360), .B1(new_n1363), .B2(new_n1301), .ZN(new_n1364));
  OAI211_X1 g1164(.A(KEYINPUT127), .B(new_n1358), .C1(new_n1364), .C2(new_n1298), .ZN(new_n1365));
  NAND2_X1  g1165(.A1(new_n1350), .A2(new_n1365), .ZN(G405));
  XNOR2_X1  g1166(.A(new_n1298), .B(new_n1318), .ZN(new_n1367));
  XNOR2_X1  g1167(.A(G375), .B(G378), .ZN(new_n1368));
  XNOR2_X1  g1168(.A(new_n1367), .B(new_n1368), .ZN(G402));
endmodule


