//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 0 1 1 1 1 0 1 0 1 1 1 0 0 0 0 0 0 1 1 1 0 1 1 0 0 1 1 0 0 1 0 1 0 0 0 1 1 0 1 1 0 0 1 1 1 0 0 0 1 1 1 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:58 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1264, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1325, new_n1326;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XOR2_X1   g0014(.A(new_n214), .B(KEYINPUT64), .Z(new_n215));
  XOR2_X1   g0015(.A(new_n215), .B(KEYINPUT0), .Z(new_n216));
  AND2_X1   g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(G20), .ZN(new_n218));
  OR2_X1    g0018(.A1(new_n201), .A2(KEYINPUT65), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n201), .A2(KEYINPUT65), .ZN(new_n220));
  NAND3_X1  g0020(.A1(new_n219), .A2(G50), .A3(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n222));
  INV_X1    g0022(.A(G68), .ZN(new_n223));
  INV_X1    g0023(.A(G238), .ZN(new_n224));
  INV_X1    g0024(.A(G77), .ZN(new_n225));
  INV_X1    g0025(.A(G244), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n222), .B1(new_n223), .B2(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(KEYINPUT66), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n230));
  NAND3_X1  g0030(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n227), .A2(KEYINPUT66), .ZN(new_n232));
  OAI21_X1  g0032(.A(new_n212), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  OAI221_X1 g0033(.A(new_n216), .B1(new_n218), .B2(new_n221), .C1(KEYINPUT1), .C2(new_n233), .ZN(new_n234));
  AOI21_X1  g0034(.A(new_n234), .B1(KEYINPUT1), .B2(new_n233), .ZN(G361));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT67), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  INV_X1    g0040(.A(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(KEYINPUT2), .B(G226), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n239), .B(new_n244), .ZN(G358));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XOR2_X1   g0046(.A(G107), .B(G116), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n202), .A2(G68), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n223), .A2(G50), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G58), .B(G77), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XOR2_X1   g0053(.A(new_n248), .B(new_n253), .Z(G351));
  INV_X1    g0054(.A(G41), .ZN(new_n255));
  INV_X1    g0055(.A(G45), .ZN(new_n256));
  AOI21_X1  g0056(.A(G1), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(G33), .A2(G41), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n258), .A2(G1), .A3(G13), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n257), .A2(new_n259), .A3(G274), .ZN(new_n260));
  INV_X1    g0060(.A(G226), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n260), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  OR2_X1    g0064(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n265));
  INV_X1    g0065(.A(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(KEYINPUT3), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT3), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n270));
  NAND4_X1  g0070(.A1(new_n265), .A2(new_n267), .A3(new_n269), .A4(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G222), .ZN(new_n273));
  XNOR2_X1  g0073(.A(KEYINPUT3), .B(G33), .ZN(new_n274));
  INV_X1    g0074(.A(G223), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(G1698), .ZN(new_n276));
  OAI221_X1 g0076(.A(new_n273), .B1(new_n225), .B2(new_n274), .C1(new_n275), .C2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n259), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n264), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(KEYINPUT10), .B1(new_n279), .B2(G190), .ZN(new_n280));
  XNOR2_X1  g0080(.A(KEYINPUT8), .B(G58), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n210), .A2(G33), .ZN(new_n282));
  INV_X1    g0082(.A(G150), .ZN(new_n283));
  NOR2_X1   g0083(.A1(G20), .A2(G33), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  OAI22_X1  g0085(.A1(new_n281), .A2(new_n282), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n286), .B1(G20), .B2(new_n203), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n217), .B1(new_n211), .B2(G33), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G13), .ZN(new_n290));
  NOR3_X1   g0090(.A1(new_n290), .A2(new_n210), .A3(G1), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n288), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n209), .A2(G20), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(G50), .ZN(new_n295));
  OAI22_X1  g0095(.A1(new_n293), .A2(new_n295), .B1(G50), .B2(new_n292), .ZN(new_n296));
  OR2_X1    g0096(.A1(new_n289), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(KEYINPUT9), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n289), .A2(new_n296), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT9), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n298), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(KEYINPUT69), .ZN(new_n303));
  INV_X1    g0103(.A(G200), .ZN(new_n304));
  OR2_X1    g0104(.A1(new_n279), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT69), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n298), .A2(new_n306), .A3(new_n301), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n280), .A2(new_n303), .A3(new_n305), .A4(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n279), .A2(G190), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n302), .A2(new_n309), .A3(new_n305), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(KEYINPUT10), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G179), .ZN(new_n313));
  AND2_X1   g0113(.A1(new_n279), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n297), .B1(new_n279), .B2(G169), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(G20), .A2(G77), .ZN(new_n318));
  INV_X1    g0118(.A(G87), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(KEYINPUT15), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT15), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(G87), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  OAI221_X1 g0124(.A(new_n318), .B1(new_n281), .B2(new_n285), .C1(new_n324), .C2(new_n282), .ZN(new_n325));
  INV_X1    g0125(.A(new_n288), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n294), .A2(G77), .ZN(new_n328));
  OAI221_X1 g0128(.A(new_n327), .B1(G77), .B2(new_n292), .C1(new_n293), .C2(new_n328), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n260), .B1(new_n226), .B2(new_n263), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n267), .A2(new_n269), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(G107), .ZN(new_n332));
  OAI221_X1 g0132(.A(new_n332), .B1(new_n271), .B2(new_n241), .C1(new_n224), .C2(new_n276), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n330), .B1(new_n333), .B2(new_n278), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n329), .B1(G169), .B2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n334), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n336), .A2(G179), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n329), .B1(G200), .B2(new_n336), .ZN(new_n340));
  INV_X1    g0140(.A(G190), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n340), .B1(new_n341), .B2(new_n336), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n312), .A2(new_n317), .A3(new_n339), .A4(new_n342), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n267), .A2(new_n269), .A3(G232), .A4(G1698), .ZN(new_n344));
  NAND2_X1  g0144(.A1(G33), .A2(G97), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n344), .B(new_n345), .C1(new_n271), .C2(new_n261), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(new_n278), .ZN(new_n347));
  AND3_X1   g0147(.A1(new_n259), .A2(G238), .A3(new_n262), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT70), .ZN(new_n349));
  AND2_X1   g0149(.A1(G33), .A2(G41), .ZN(new_n350));
  NAND2_X1  g0150(.A1(G1), .A2(G13), .ZN(new_n351));
  OAI21_X1  g0151(.A(G274), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n349), .B1(new_n352), .B2(new_n262), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n257), .A2(new_n259), .A3(KEYINPUT70), .A4(G274), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n348), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT13), .ZN(new_n356));
  AND3_X1   g0156(.A1(new_n347), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n356), .B1(new_n347), .B2(new_n355), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(G169), .ZN(new_n360));
  OAI21_X1  g0160(.A(KEYINPUT14), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT14), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n362), .B(G169), .C1(new_n357), .C2(new_n358), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT73), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n364), .B1(new_n359), .B2(G179), .ZN(new_n365));
  NOR4_X1   g0165(.A1(new_n357), .A2(new_n358), .A3(KEYINPUT73), .A4(new_n313), .ZN(new_n366));
  OAI211_X1 g0166(.A(new_n361), .B(new_n363), .C1(new_n365), .C2(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n210), .A2(G33), .A3(G77), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT71), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n223), .A2(G20), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n284), .A2(G50), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n369), .B1(new_n368), .B2(new_n370), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n326), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT11), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  OAI211_X1 g0177(.A(new_n326), .B(KEYINPUT11), .C1(new_n373), .C2(new_n374), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  OR2_X1    g0179(.A1(new_n379), .A2(KEYINPUT72), .ZN(new_n380));
  NOR3_X1   g0180(.A1(new_n292), .A2(KEYINPUT12), .A3(G68), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT12), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n382), .B1(new_n291), .B2(new_n223), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n294), .A2(G68), .ZN(new_n384));
  OAI22_X1  g0184(.A1(new_n381), .A2(new_n383), .B1(new_n293), .B2(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n385), .B1(new_n379), .B2(KEYINPUT72), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n380), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n367), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(G200), .B1(new_n357), .B2(new_n358), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n347), .A2(new_n355), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(KEYINPUT13), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n347), .A2(new_n355), .A3(new_n356), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n391), .A2(G190), .A3(new_n392), .ZN(new_n393));
  AND4_X1   g0193(.A1(new_n380), .A2(new_n389), .A3(new_n393), .A4(new_n386), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n388), .A2(new_n395), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n343), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT17), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT78), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n267), .A2(new_n269), .A3(G226), .A4(G1698), .ZN(new_n400));
  NAND2_X1  g0200(.A1(G33), .A2(G87), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n400), .B(new_n401), .C1(new_n271), .C2(new_n275), .ZN(new_n402));
  AND2_X1   g0202(.A1(new_n402), .A2(new_n278), .ZN(new_n403));
  OAI21_X1  g0203(.A(KEYINPUT77), .B1(new_n263), .B2(new_n241), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT77), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n259), .A2(new_n262), .A3(new_n405), .A4(G232), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n404), .A2(new_n260), .A3(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n399), .B1(new_n403), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n255), .A2(new_n256), .ZN(new_n409));
  AOI22_X1  g0209(.A1(new_n209), .A2(new_n409), .B1(new_n217), .B2(new_n258), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n405), .B1(new_n410), .B2(G232), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n406), .A2(new_n260), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n402), .A2(new_n278), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n413), .A2(new_n414), .A3(KEYINPUT78), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n408), .A2(new_n304), .A3(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT80), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n403), .A2(KEYINPUT76), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT76), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n414), .A2(new_n419), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n407), .A2(G190), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n418), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  AND3_X1   g0222(.A1(new_n416), .A2(new_n417), .A3(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n417), .B1(new_n416), .B2(new_n422), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(G58), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n426), .A2(new_n223), .ZN(new_n427));
  OAI21_X1  g0227(.A(G20), .B1(new_n427), .B2(new_n201), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n284), .A2(G159), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT16), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n331), .A2(KEYINPUT74), .A3(KEYINPUT7), .A4(new_n210), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT7), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n434), .B1(new_n274), .B2(G20), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(G20), .B1(new_n267), .B2(new_n269), .ZN(new_n437));
  AOI21_X1  g0237(.A(KEYINPUT74), .B1(new_n437), .B2(KEYINPUT7), .ZN(new_n438));
  OAI211_X1 g0238(.A(KEYINPUT75), .B(G68), .C1(new_n436), .C2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n331), .A2(KEYINPUT7), .A3(new_n210), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT74), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n443), .A2(new_n435), .A3(new_n433), .ZN(new_n444));
  AOI21_X1  g0244(.A(KEYINPUT75), .B1(new_n444), .B2(G68), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n432), .B1(new_n440), .B2(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n223), .B1(new_n435), .B2(new_n441), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n431), .B1(new_n447), .B2(new_n430), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n446), .A2(new_n448), .A3(new_n326), .ZN(new_n449));
  INV_X1    g0249(.A(new_n281), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(new_n294), .ZN(new_n451));
  OAI22_X1  g0251(.A1(new_n293), .A2(new_n451), .B1(new_n292), .B2(new_n450), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n449), .A2(new_n453), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n398), .B1(new_n425), .B2(new_n454), .ZN(new_n455));
  AND3_X1   g0255(.A1(new_n413), .A2(new_n414), .A3(KEYINPUT78), .ZN(new_n456));
  AOI21_X1  g0256(.A(KEYINPUT78), .B1(new_n413), .B2(new_n414), .ZN(new_n457));
  NOR3_X1   g0257(.A1(new_n456), .A2(new_n457), .A3(G169), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n407), .A2(G179), .ZN(new_n459));
  AND3_X1   g0259(.A1(new_n418), .A2(new_n420), .A3(new_n459), .ZN(new_n460));
  OAI21_X1  g0260(.A(KEYINPUT79), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n408), .A2(new_n360), .A3(new_n415), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n418), .A2(new_n420), .A3(new_n459), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT79), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n461), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g0266(.A(G68), .B1(new_n436), .B2(new_n438), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT75), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(new_n439), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n288), .B1(new_n470), .B2(new_n432), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n452), .B1(new_n471), .B2(new_n448), .ZN(new_n472));
  OAI21_X1  g0272(.A(KEYINPUT18), .B1(new_n466), .B2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT18), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n454), .A2(new_n461), .A3(new_n474), .A4(new_n465), .ZN(new_n475));
  NOR3_X1   g0275(.A1(new_n456), .A2(new_n457), .A3(G200), .ZN(new_n476));
  AND3_X1   g0276(.A1(new_n418), .A2(new_n420), .A3(new_n421), .ZN(new_n477));
  OAI21_X1  g0277(.A(KEYINPUT80), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n416), .A2(new_n417), .A3(new_n422), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n480), .A2(KEYINPUT17), .A3(new_n472), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n455), .A2(new_n473), .A3(new_n475), .A4(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n397), .A2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n209), .A2(G33), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n288), .A2(new_n292), .A3(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(G116), .ZN(new_n489));
  INV_X1    g0289(.A(G116), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n291), .A2(new_n490), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n210), .A2(G116), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n288), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(G33), .A2(G283), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n494), .B(new_n210), .C1(G33), .C2(new_n205), .ZN(new_n495));
  AND3_X1   g0295(.A1(new_n493), .A2(KEYINPUT20), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(KEYINPUT20), .B1(new_n493), .B2(new_n495), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n489), .B(new_n491), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n274), .A2(G264), .A3(G1698), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n331), .A2(G303), .ZN(new_n500));
  INV_X1    g0300(.A(G257), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n499), .B(new_n500), .C1(new_n501), .C2(new_n271), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n278), .ZN(new_n503));
  XNOR2_X1  g0303(.A(KEYINPUT5), .B(G41), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n209), .A2(G45), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n507), .A2(G270), .A3(new_n259), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n504), .A2(new_n506), .A3(G274), .A4(new_n259), .ZN(new_n509));
  AND2_X1   g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n360), .B1(new_n503), .B2(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(KEYINPUT86), .B1(new_n498), .B2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT21), .ZN(new_n513));
  AND2_X1   g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n508), .A2(new_n509), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n515), .B1(new_n278), .B2(new_n502), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n498), .A2(G179), .A3(new_n516), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n517), .B1(new_n512), .B2(new_n513), .ZN(new_n518));
  AND2_X1   g0318(.A1(new_n516), .A2(G190), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n516), .A2(new_n304), .ZN(new_n520));
  NOR3_X1   g0320(.A1(new_n519), .A2(new_n520), .A3(new_n498), .ZN(new_n521));
  NOR3_X1   g0321(.A1(new_n514), .A2(new_n518), .A3(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n274), .A2(G257), .A3(G1698), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(KEYINPUT89), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT89), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n274), .A2(new_n525), .A3(G257), .A4(G1698), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(G250), .ZN(new_n528));
  INV_X1    g0328(.A(G294), .ZN(new_n529));
  OAI22_X1  g0329(.A1(new_n271), .A2(new_n528), .B1(new_n266), .B2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n527), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n278), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n278), .B1(new_n506), .B2(new_n504), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(G264), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n533), .A2(G179), .A3(new_n509), .A4(new_n535), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n259), .B1(new_n527), .B2(new_n531), .ZN(new_n537));
  INV_X1    g0337(.A(new_n509), .ZN(new_n538));
  INV_X1    g0338(.A(new_n535), .ZN(new_n539));
  NOR3_X1   g0339(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n536), .B1(new_n540), .B2(new_n360), .ZN(new_n541));
  AOI21_X1  g0341(.A(KEYINPUT25), .B1(new_n291), .B2(new_n206), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n291), .A2(KEYINPUT25), .A3(new_n206), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n488), .A2(G107), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n274), .A2(new_n210), .A3(G87), .ZN(new_n546));
  AND2_X1   g0346(.A1(KEYINPUT87), .A2(KEYINPUT22), .ZN(new_n547));
  NOR2_X1   g0347(.A1(KEYINPUT87), .A2(KEYINPUT22), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n274), .A2(new_n210), .A3(G87), .A4(new_n547), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT23), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n552), .B1(G20), .B2(new_n206), .ZN(new_n553));
  OR2_X1    g0353(.A1(new_n553), .A2(KEYINPUT88), .ZN(new_n554));
  OAI211_X1 g0354(.A(KEYINPUT88), .B(KEYINPUT23), .C1(new_n210), .C2(G107), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n210), .A2(G33), .A3(G116), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n552), .A2(new_n206), .A3(G20), .ZN(new_n557));
  AND3_X1   g0357(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n550), .A2(new_n551), .A3(new_n554), .A4(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(KEYINPUT24), .ZN(new_n560));
  AND2_X1   g0360(.A1(new_n558), .A2(new_n554), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT24), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n561), .A2(new_n562), .A3(new_n551), .A4(new_n550), .ZN(new_n563));
  AND2_X1   g0363(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n545), .B1(new_n564), .B2(new_n288), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n541), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n533), .A2(new_n509), .A3(new_n535), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(G200), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n540), .A2(G190), .ZN(new_n569));
  INV_X1    g0369(.A(new_n545), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n560), .A2(new_n563), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n570), .B1(new_n571), .B2(new_n326), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n568), .A2(new_n569), .A3(new_n572), .ZN(new_n573));
  AND2_X1   g0373(.A1(new_n566), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n274), .A2(new_n210), .A3(G68), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT19), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n576), .B1(new_n282), .B2(new_n205), .ZN(new_n577));
  NAND3_X1  g0377(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT84), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n578), .A2(new_n579), .A3(new_n210), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n319), .A2(new_n205), .A3(new_n206), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n579), .B1(new_n578), .B2(new_n210), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n575), .B(new_n577), .C1(new_n582), .C2(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n288), .B1(new_n584), .B2(KEYINPUT85), .ZN(new_n585));
  OR2_X1    g0385(.A1(new_n582), .A2(new_n583), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT85), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n586), .A2(new_n587), .A3(new_n575), .A4(new_n577), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n324), .A2(new_n291), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n488), .A2(G87), .ZN(new_n591));
  AND3_X1   g0391(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n259), .A2(G274), .A3(new_n506), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n259), .A2(G250), .A3(new_n505), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n274), .A2(G244), .A3(G1698), .ZN(new_n596));
  NAND2_X1  g0396(.A1(G33), .A2(G116), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n596), .B(new_n597), .C1(new_n224), .C2(new_n271), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n595), .B1(new_n598), .B2(new_n278), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n341), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n600), .B1(G200), .B2(new_n599), .ZN(new_n601));
  AOI211_X1 g0401(.A(G179), .B(new_n595), .C1(new_n598), .C2(new_n278), .ZN(new_n602));
  INV_X1    g0402(.A(new_n599), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n602), .B1(new_n360), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n488), .A2(new_n323), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n589), .A2(new_n605), .A3(new_n590), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n592), .A2(new_n601), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n435), .A2(new_n441), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n608), .A2(G107), .B1(G77), .B2(new_n284), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n206), .A2(KEYINPUT6), .A3(G97), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(KEYINPUT81), .ZN(new_n611));
  OR2_X1    g0411(.A1(new_n610), .A2(KEYINPUT81), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT82), .ZN(new_n613));
  NAND2_X1  g0413(.A1(G97), .A2(G107), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n207), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT6), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n613), .B1(new_n207), .B2(new_n614), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n611), .B(new_n612), .C1(new_n617), .C2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(G20), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n609), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n326), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n292), .A2(G97), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n624), .B1(new_n487), .B2(new_n205), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n622), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n538), .B1(G257), .B2(new_n534), .ZN(new_n628));
  XOR2_X1   g0428(.A(KEYINPUT68), .B(G1698), .Z(new_n629));
  NAND4_X1  g0429(.A1(new_n629), .A2(KEYINPUT4), .A3(G244), .A4(new_n274), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n274), .A2(G250), .A3(G1698), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n630), .A2(new_n494), .A3(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT4), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n633), .B1(new_n271), .B2(new_n226), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT83), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  OAI211_X1 g0436(.A(KEYINPUT83), .B(new_n633), .C1(new_n271), .C2(new_n226), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n632), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n313), .B(new_n628), .C1(new_n638), .C2(new_n259), .ZN(new_n639));
  INV_X1    g0439(.A(new_n628), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n636), .A2(new_n637), .ZN(new_n641));
  INV_X1    g0441(.A(new_n632), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n640), .B1(new_n643), .B2(new_n278), .ZN(new_n644));
  OAI211_X1 g0444(.A(new_n627), .B(new_n639), .C1(G169), .C2(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n625), .B1(new_n621), .B2(new_n326), .ZN(new_n646));
  OAI211_X1 g0446(.A(G190), .B(new_n628), .C1(new_n638), .C2(new_n259), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n646), .B(new_n647), .C1(new_n644), .C2(new_n304), .ZN(new_n648));
  AND3_X1   g0448(.A1(new_n607), .A2(new_n645), .A3(new_n648), .ZN(new_n649));
  AND4_X1   g0449(.A1(new_n485), .A2(new_n522), .A3(new_n574), .A4(new_n649), .ZN(G372));
  NOR2_X1   g0450(.A1(new_n514), .A2(new_n518), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT91), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n541), .A2(new_n652), .A3(new_n565), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n652), .B1(new_n541), .B2(new_n565), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n651), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n592), .A2(new_n601), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT90), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n603), .A2(new_n657), .A3(new_n360), .ZN(new_n658));
  INV_X1    g0458(.A(new_n602), .ZN(new_n659));
  OAI21_X1  g0459(.A(KEYINPUT90), .B1(new_n599), .B2(G169), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n606), .A2(new_n658), .A3(new_n659), .A4(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n656), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  AND3_X1   g0463(.A1(new_n645), .A2(new_n573), .A3(new_n648), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n655), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n628), .B1(new_n638), .B2(new_n259), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n646), .B1(new_n360), .B2(new_n666), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n667), .A2(new_n656), .A3(new_n661), .A4(new_n639), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n661), .B1(new_n668), .B2(KEYINPUT26), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT26), .ZN(new_n670));
  INV_X1    g0470(.A(new_n645), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n670), .B1(new_n671), .B2(new_n607), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n484), .B1(new_n665), .B2(new_n673), .ZN(new_n674));
  AND3_X1   g0474(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n464), .B1(new_n462), .B2(new_n463), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n474), .B1(new_n677), .B2(new_n454), .ZN(new_n678));
  NOR4_X1   g0478(.A1(new_n472), .A2(new_n675), .A3(new_n676), .A4(KEYINPUT18), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NOR3_X1   g0481(.A1(new_n425), .A2(new_n398), .A3(new_n454), .ZN(new_n682));
  AOI21_X1  g0482(.A(KEYINPUT17), .B1(new_n480), .B2(new_n472), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n394), .B1(new_n388), .B2(new_n339), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n681), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n312), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n317), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n674), .A2(new_n688), .ZN(G369));
  OR2_X1    g0489(.A1(new_n653), .A2(new_n654), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n691));
  OR2_X1    g0491(.A1(new_n691), .A2(KEYINPUT27), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(KEYINPUT27), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n692), .A2(G213), .A3(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(G343), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n690), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n565), .A2(new_n696), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n566), .A2(new_n573), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(KEYINPUT92), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT92), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n566), .A2(new_n573), .A3(new_n698), .A4(new_n701), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n541), .A2(new_n565), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n703), .A2(KEYINPUT93), .A3(new_n696), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT93), .ZN(new_n705));
  INV_X1    g0505(.A(new_n696), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n705), .B1(new_n566), .B2(new_n706), .ZN(new_n707));
  AOI22_X1  g0507(.A1(new_n700), .A2(new_n702), .B1(new_n704), .B2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n706), .B1(new_n514), .B2(new_n518), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n697), .B1(new_n709), .B2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(G330), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n498), .A2(new_n696), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n522), .A2(new_n714), .ZN(new_n715));
  OAI211_X1 g0515(.A(new_n498), .B(new_n696), .C1(new_n514), .C2(new_n518), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n713), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n709), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n712), .A2(new_n718), .ZN(G399));
  INV_X1    g0519(.A(new_n213), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(G41), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n581), .A2(G116), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n722), .A2(G1), .A3(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n724), .B1(new_n221), .B2(new_n722), .ZN(new_n725));
  XNOR2_X1  g0525(.A(new_n725), .B(KEYINPUT28), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n663), .A2(new_n573), .A3(new_n645), .A4(new_n648), .ZN(new_n727));
  NOR3_X1   g0527(.A1(new_n703), .A2(new_n514), .A3(new_n518), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n661), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n668), .A2(new_n670), .ZN(new_n730));
  AOI21_X1  g0530(.A(KEYINPUT26), .B1(new_n671), .B2(new_n607), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n706), .B1(new_n729), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(KEYINPUT29), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT30), .ZN(new_n735));
  NOR3_X1   g0535(.A1(new_n603), .A2(new_n537), .A3(new_n539), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(new_n644), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n516), .A2(KEYINPUT94), .A3(G179), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n503), .A2(new_n510), .A3(G179), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT94), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n735), .B1(new_n737), .B2(new_n742), .ZN(new_n743));
  AND2_X1   g0543(.A1(new_n738), .A2(new_n741), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n530), .B1(new_n526), .B2(new_n524), .ZN(new_n745));
  OAI211_X1 g0545(.A(new_n599), .B(new_n535), .C1(new_n745), .C2(new_n259), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n666), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n744), .A2(new_n747), .A3(KEYINPUT30), .ZN(new_n748));
  NOR3_X1   g0548(.A1(new_n516), .A2(G179), .A3(new_n599), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n749), .A2(new_n666), .A3(new_n567), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n743), .A2(new_n748), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(new_n696), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT31), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND4_X1  g0554(.A1(new_n649), .A2(new_n522), .A3(new_n574), .A4(new_n706), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n751), .A2(KEYINPUT31), .A3(new_n696), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n754), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G330), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n696), .B1(new_n665), .B2(new_n673), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT29), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n734), .A2(new_n758), .A3(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n726), .B1(new_n763), .B2(G1), .ZN(G364));
  NAND3_X1  g0564(.A1(new_n715), .A2(new_n713), .A3(new_n716), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n290), .A2(G20), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n209), .B1(new_n766), .B2(G45), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n721), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n765), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n717), .A2(KEYINPUT95), .ZN(new_n772));
  INV_X1    g0572(.A(KEYINPUT95), .ZN(new_n773));
  AOI211_X1 g0573(.A(new_n773), .B(new_n713), .C1(new_n715), .C2(new_n716), .ZN(new_n774));
  NOR3_X1   g0574(.A1(new_n771), .A2(new_n772), .A3(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(G13), .A2(G33), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(G20), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n715), .A2(new_n716), .A3(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n351), .B1(G20), .B2(new_n360), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n210), .A2(G179), .ZN(new_n782));
  NOR2_X1   g0582(.A1(G190), .A2(G200), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n784), .B(KEYINPUT97), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n782), .A2(new_n341), .A3(G200), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  AOI22_X1  g0587(.A1(new_n785), .A2(G329), .B1(G283), .B2(new_n787), .ZN(new_n788));
  XOR2_X1   g0588(.A(new_n788), .B(KEYINPUT98), .Z(new_n789));
  NAND3_X1  g0589(.A1(new_n782), .A2(G190), .A3(G200), .ZN(new_n790));
  INV_X1    g0590(.A(G303), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n331), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  XOR2_X1   g0592(.A(new_n792), .B(KEYINPUT96), .Z(new_n793));
  NOR2_X1   g0593(.A1(new_n210), .A2(new_n313), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n794), .A2(G190), .A3(new_n304), .ZN(new_n795));
  INV_X1    g0595(.A(G322), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n794), .A2(new_n783), .ZN(new_n797));
  INV_X1    g0597(.A(G311), .ZN(new_n798));
  OAI22_X1  g0598(.A1(new_n795), .A2(new_n796), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n794), .A2(new_n341), .A3(G200), .ZN(new_n800));
  XOR2_X1   g0600(.A(KEYINPUT33), .B(G317), .Z(new_n801));
  NAND3_X1  g0601(.A1(new_n794), .A2(G190), .A3(G200), .ZN(new_n802));
  INV_X1    g0602(.A(G326), .ZN(new_n803));
  OAI22_X1  g0603(.A1(new_n800), .A2(new_n801), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NOR3_X1   g0604(.A1(new_n341), .A2(G179), .A3(G200), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n805), .A2(new_n210), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n799), .B(new_n804), .C1(G294), .C2(new_n807), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n789), .A2(new_n793), .A3(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(G159), .ZN(new_n810));
  NOR3_X1   g0610(.A1(new_n784), .A2(KEYINPUT32), .A3(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n800), .ZN(new_n812));
  AOI22_X1  g0612(.A1(G68), .A2(new_n812), .B1(new_n787), .B2(G107), .ZN(new_n813));
  INV_X1    g0613(.A(new_n790), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(G87), .ZN(new_n815));
  OAI211_X1 g0615(.A(new_n813), .B(new_n815), .C1(new_n205), .C2(new_n806), .ZN(new_n816));
  OAI21_X1  g0616(.A(KEYINPUT32), .B1(new_n784), .B2(new_n810), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n817), .B1(new_n202), .B2(new_n802), .ZN(new_n818));
  OAI221_X1 g0618(.A(new_n274), .B1(new_n797), .B2(new_n225), .C1(new_n426), .C2(new_n795), .ZN(new_n819));
  OR4_X1    g0619(.A1(new_n811), .A2(new_n816), .A3(new_n818), .A4(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n781), .B1(new_n809), .B2(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n778), .A2(new_n780), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n213), .A2(G355), .A3(new_n274), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n720), .A2(new_n274), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n824), .B1(G45), .B2(new_n221), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n253), .A2(new_n256), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n823), .B1(G116), .B2(new_n213), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n770), .B(new_n821), .C1(new_n822), .C2(new_n827), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n828), .B(KEYINPUT99), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n775), .B1(new_n779), .B2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(G396));
  NAND2_X1  g0631(.A1(new_n329), .A2(new_n696), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n339), .A2(new_n342), .A3(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT101), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND4_X1  g0635(.A1(new_n339), .A2(new_n342), .A3(KEYINPUT101), .A4(new_n832), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n759), .A2(new_n837), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n835), .B(new_n836), .C1(new_n339), .C2(new_n706), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n838), .B1(new_n759), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n769), .B1(new_n840), .B2(new_n758), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n841), .B1(new_n758), .B2(new_n840), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n780), .A2(new_n776), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n769), .B1(G77), .B2(new_n844), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n806), .A2(new_n205), .ZN(new_n846));
  OAI22_X1  g0646(.A1(new_n802), .A2(new_n791), .B1(new_n790), .B2(new_n206), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n846), .B(new_n847), .C1(G87), .C2(new_n787), .ZN(new_n848));
  AND2_X1   g0648(.A1(new_n800), .A2(KEYINPUT100), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n800), .A2(KEYINPUT100), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(G283), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n785), .A2(G311), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n331), .B1(new_n795), .B2(new_n529), .ZN(new_n855));
  INV_X1    g0655(.A(new_n797), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n855), .B1(G116), .B2(new_n856), .ZN(new_n857));
  NAND4_X1  g0657(.A1(new_n848), .A2(new_n853), .A3(new_n854), .A4(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n787), .A2(G68), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n859), .B1(new_n202), .B2(new_n790), .ZN(new_n860));
  AOI211_X1 g0660(.A(new_n331), .B(new_n860), .C1(G58), .C2(new_n807), .ZN(new_n861));
  INV_X1    g0661(.A(new_n795), .ZN(new_n862));
  AOI22_X1  g0662(.A1(new_n862), .A2(G143), .B1(new_n856), .B2(G159), .ZN(new_n863));
  INV_X1    g0663(.A(G137), .ZN(new_n864));
  OAI221_X1 g0664(.A(new_n863), .B1(new_n864), .B2(new_n802), .C1(new_n283), .C2(new_n800), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT34), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(G132), .ZN(new_n868));
  INV_X1    g0668(.A(new_n785), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n861), .B(new_n867), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n865), .A2(new_n866), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n858), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n845), .B1(new_n872), .B2(new_n780), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n873), .B1(new_n839), .B2(new_n777), .ZN(new_n874));
  AND2_X1   g0674(.A1(new_n842), .A2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(G384));
  NOR2_X1   g0676(.A1(new_n766), .A2(new_n209), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n446), .A2(new_n326), .ZN(new_n878));
  INV_X1    g0678(.A(new_n430), .ZN(new_n879));
  AOI21_X1  g0679(.A(KEYINPUT16), .B1(new_n470), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n453), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n881), .A2(new_n465), .A3(new_n461), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n472), .B1(new_n424), .B2(new_n423), .ZN(new_n883));
  INV_X1    g0683(.A(new_n694), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n882), .A2(new_n883), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(KEYINPUT37), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n454), .A2(new_n465), .A3(new_n461), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT37), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n454), .A2(new_n884), .ZN(new_n890));
  NAND4_X1  g0690(.A1(new_n883), .A2(new_n888), .A3(new_n889), .A4(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n887), .A2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n885), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n482), .A2(new_n893), .ZN(new_n894));
  AND3_X1   g0694(.A1(new_n892), .A2(new_n894), .A3(KEYINPUT38), .ZN(new_n895));
  INV_X1    g0695(.A(new_n890), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n482), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n883), .A2(new_n888), .A3(new_n890), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(KEYINPUT37), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n891), .ZN(new_n900));
  AOI21_X1  g0700(.A(KEYINPUT38), .B1(new_n897), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(KEYINPUT104), .B1(new_n895), .B2(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n892), .A2(new_n894), .A3(KEYINPUT38), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT104), .ZN(new_n904));
  AOI22_X1  g0704(.A1(new_n482), .A2(new_n896), .B1(new_n899), .B2(new_n891), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n903), .B(new_n904), .C1(KEYINPUT38), .C2(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n706), .B1(new_n380), .B2(new_n386), .ZN(new_n907));
  AOI211_X1 g0707(.A(new_n394), .B(new_n907), .C1(new_n367), .C2(new_n387), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n367), .A2(new_n907), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(KEYINPUT102), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT102), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n912), .B(new_n909), .C1(new_n396), .C2(new_n907), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n757), .A2(new_n911), .A3(new_n839), .A4(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT40), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n902), .A2(new_n906), .A3(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT38), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n885), .B1(new_n684), .B2(new_n680), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n480), .A2(new_n472), .B1(new_n881), .B2(new_n884), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n889), .B1(new_n920), .B2(new_n882), .ZN(new_n921));
  AND4_X1   g0721(.A1(new_n889), .A2(new_n883), .A3(new_n888), .A4(new_n890), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n918), .B1(new_n919), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n914), .B1(new_n924), .B2(new_n903), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n917), .B1(KEYINPUT40), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n485), .A2(new_n757), .ZN(new_n927));
  OR2_X1    g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n926), .A2(new_n927), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n928), .A2(G330), .A3(new_n929), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n930), .B(KEYINPUT105), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n339), .A2(new_n696), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n838), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n911), .A2(new_n913), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(KEYINPUT38), .B1(new_n892), .B2(new_n894), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n895), .A2(new_n938), .ZN(new_n939));
  OAI22_X1  g0739(.A1(new_n937), .A2(new_n939), .B1(new_n680), .B2(new_n884), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n388), .A2(new_n696), .ZN(new_n941));
  OAI21_X1  g0741(.A(KEYINPUT39), .B1(new_n895), .B2(new_n938), .ZN(new_n942));
  XNOR2_X1  g0742(.A(KEYINPUT103), .B(KEYINPUT39), .ZN(new_n943));
  OAI211_X1 g0743(.A(new_n903), .B(new_n943), .C1(KEYINPUT38), .C2(new_n905), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n940), .B1(new_n941), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n484), .B1(new_n734), .B2(new_n761), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n947), .A2(new_n688), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n946), .B(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n877), .B1(new_n931), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n931), .B2(new_n949), .ZN(new_n951));
  AOI211_X1 g0751(.A(new_n490), .B(new_n218), .C1(new_n619), .C2(KEYINPUT35), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(KEYINPUT35), .B2(new_n619), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(KEYINPUT36), .ZN(new_n954));
  OAI21_X1  g0754(.A(G77), .B1(new_n426), .B2(new_n223), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n249), .B1(new_n221), .B2(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n956), .A2(G1), .A3(new_n290), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n951), .A2(new_n954), .A3(new_n957), .ZN(G367));
  OAI21_X1  g0758(.A(new_n822), .B1(new_n213), .B2(new_n324), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n959), .B1(new_n824), .B2(new_n238), .ZN(new_n960));
  INV_X1    g0760(.A(new_n784), .ZN(new_n961));
  AOI22_X1  g0761(.A1(G50), .A2(new_n856), .B1(new_n961), .B2(G137), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n962), .B(new_n274), .C1(new_n283), .C2(new_n795), .ZN(new_n963));
  INV_X1    g0763(.A(new_n802), .ZN(new_n964));
  AOI22_X1  g0764(.A1(G143), .A2(new_n964), .B1(new_n787), .B2(G77), .ZN(new_n965));
  OAI221_X1 g0765(.A(new_n965), .B1(new_n426), .B2(new_n790), .C1(new_n223), .C2(new_n806), .ZN(new_n966));
  AOI211_X1 g0766(.A(new_n963), .B(new_n966), .C1(G159), .C2(new_n852), .ZN(new_n967));
  AOI22_X1  g0767(.A1(G107), .A2(new_n807), .B1(new_n964), .B2(G311), .ZN(new_n968));
  OAI221_X1 g0768(.A(new_n968), .B1(new_n205), .B2(new_n786), .C1(new_n851), .C2(new_n529), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT46), .ZN(new_n970));
  NOR3_X1   g0770(.A1(new_n790), .A2(new_n970), .A3(new_n490), .ZN(new_n971));
  AOI22_X1  g0771(.A1(G283), .A2(new_n856), .B1(new_n961), .B2(G317), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n274), .B1(new_n862), .B2(G303), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n970), .B1(new_n790), .B2(new_n490), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n972), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  NOR3_X1   g0775(.A1(new_n969), .A2(new_n971), .A3(new_n975), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n967), .A2(new_n976), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n977), .B(KEYINPUT47), .Z(new_n978));
  AOI211_X1 g0778(.A(new_n770), .B(new_n960), .C1(new_n978), .C2(new_n780), .ZN(new_n979));
  OR2_X1    g0779(.A1(new_n592), .A2(new_n706), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n663), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(new_n661), .B2(new_n980), .ZN(new_n982));
  INV_X1    g0782(.A(new_n778), .ZN(new_n983));
  OR2_X1    g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n979), .A2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT110), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT44), .ZN(new_n987));
  OAI211_X1 g0787(.A(new_n645), .B(new_n648), .C1(new_n646), .C2(new_n706), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n645), .B2(new_n706), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT106), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n987), .B1(new_n712), .B2(new_n990), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n708), .A2(new_n710), .B1(new_n690), .B2(new_n696), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT106), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n989), .B(new_n993), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n992), .A2(new_n994), .A3(KEYINPUT44), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n991), .A2(new_n995), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n712), .A2(KEYINPUT45), .A3(new_n990), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT45), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(new_n992), .B2(new_n994), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  AND3_X1   g0800(.A1(new_n996), .A2(new_n1000), .A3(new_n718), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n718), .B1(new_n996), .B2(new_n1000), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n709), .A2(new_n711), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n708), .A2(new_n710), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n772), .A2(new_n774), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1004), .A2(new_n717), .A3(new_n1005), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1008), .A2(KEYINPUT109), .A3(new_n1009), .ZN(new_n1010));
  OR2_X1    g0810(.A1(new_n1009), .A2(KEYINPUT109), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n762), .B1(new_n1003), .B2(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(KEYINPUT108), .B(KEYINPUT41), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n721), .B(new_n1014), .Z(new_n1015));
  OAI21_X1  g0815(.A(new_n986), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n996), .A2(new_n1000), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n718), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n762), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n996), .A2(new_n1000), .A3(new_n718), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1019), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1022), .A2(new_n763), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1015), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1023), .A2(KEYINPUT110), .A3(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n768), .B1(new_n1016), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1018), .A2(new_n990), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT107), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n982), .A2(KEYINPUT43), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1028), .B(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n982), .A2(KEYINPUT43), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n990), .A2(new_n709), .A3(new_n711), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1032), .A2(KEYINPUT42), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n671), .B1(new_n990), .B2(new_n703), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1033), .B1(new_n1034), .B2(new_n696), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n1032), .A2(KEYINPUT42), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1031), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1030), .B(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n1038), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n985), .B1(new_n1026), .B2(new_n1039), .ZN(G387));
  NOR2_X1   g0840(.A1(new_n1020), .A2(new_n722), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1041), .B1(new_n763), .B2(new_n1012), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n708), .A2(new_n778), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n723), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1044), .A2(new_n213), .A3(new_n274), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1045), .B1(G107), .B2(new_n213), .ZN(new_n1046));
  AOI211_X1 g0846(.A(G45), .B(new_n1044), .C1(G68), .C2(G77), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n281), .A2(G50), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT50), .ZN(new_n1049));
  AOI211_X1 g0849(.A(new_n720), .B(new_n274), .C1(new_n1047), .C2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n244), .A2(G45), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1046), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n822), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n769), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n331), .B1(new_n961), .B2(G150), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n1055), .B1(new_n225), .B2(new_n790), .C1(new_n205), .C2(new_n786), .ZN(new_n1056));
  XOR2_X1   g0856(.A(new_n1056), .B(KEYINPUT111), .Z(new_n1057));
  AOI22_X1  g0857(.A1(new_n862), .A2(G50), .B1(new_n856), .B2(G68), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(new_n281), .B2(new_n800), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n806), .A2(new_n324), .B1(new_n802), .B2(new_n810), .ZN(new_n1060));
  NOR3_X1   g0860(.A1(new_n1057), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT112), .Z(new_n1062));
  AOI21_X1  g0862(.A(new_n274), .B1(new_n961), .B2(G326), .ZN(new_n1063));
  INV_X1    g0863(.A(G283), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n806), .A2(new_n1064), .B1(new_n790), .B2(new_n529), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n862), .A2(G317), .B1(new_n856), .B2(G303), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n1066), .B1(new_n796), .B2(new_n802), .C1(new_n851), .C2(new_n798), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT48), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1065), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n1068), .B2(new_n1067), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT49), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n1063), .B1(new_n490), .B2(new_n786), .C1(new_n1070), .C2(new_n1071), .ZN(new_n1072));
  AND2_X1   g0872(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1062), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1054), .B1(new_n1074), .B2(new_n780), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n1012), .A2(new_n768), .B1(new_n1043), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1042), .A2(new_n1076), .ZN(G393));
  NAND2_X1  g0877(.A1(new_n824), .A2(new_n248), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1053), .B1(G97), .B2(new_n720), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n770), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n806), .A2(new_n490), .B1(new_n797), .B2(new_n529), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n862), .A2(G311), .B1(new_n964), .B2(G317), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT52), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n1081), .B(new_n1083), .C1(G303), .C2(new_n852), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n331), .B1(new_n784), .B2(new_n796), .C1(new_n206), .C2(new_n786), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1085), .B1(G283), .B2(new_n814), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1086), .B(KEYINPUT113), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n795), .A2(new_n810), .B1(new_n802), .B2(new_n283), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1088), .B(KEYINPUT51), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n331), .B1(new_n961), .B2(G143), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(new_n281), .B2(new_n797), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n807), .A2(G77), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n1092), .B1(new_n223), .B2(new_n790), .C1(new_n319), .C2(new_n786), .ZN(new_n1093));
  AOI211_X1 g0893(.A(new_n1091), .B(new_n1093), .C1(G50), .C2(new_n852), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n1084), .A2(new_n1087), .B1(new_n1089), .B2(new_n1094), .ZN(new_n1095));
  OAI221_X1 g0895(.A(new_n1080), .B1(new_n781), .B2(new_n1095), .C1(new_n990), .C2(new_n983), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1096), .B1(new_n1097), .B2(new_n767), .ZN(new_n1098));
  OR2_X1    g0898(.A1(new_n1003), .A2(new_n1020), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n722), .B1(new_n1003), .B2(new_n1020), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1098), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(G390));
  AOI21_X1  g0902(.A(new_n932), .B1(new_n759), .B2(new_n837), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n1103), .A2(new_n935), .B1(new_n388), .B2(new_n696), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1104), .A2(new_n942), .A3(new_n944), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n706), .B(new_n837), .C1(new_n729), .C2(new_n732), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(new_n933), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n941), .B1(new_n1107), .B2(new_n936), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1108), .A2(new_n902), .A3(new_n906), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1105), .A2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n757), .A2(G330), .A3(new_n839), .ZN(new_n1111));
  OR3_X1    g0911(.A1(new_n1111), .A2(KEYINPUT114), .A3(new_n935), .ZN(new_n1112));
  OAI21_X1  g0912(.A(KEYINPUT114), .B1(new_n1111), .B2(new_n935), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1110), .A2(new_n1115), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n1105), .B(new_n1109), .C1(new_n935), .C2(new_n1111), .ZN(new_n1117));
  AND2_X1   g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT116), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n839), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT115), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1120), .B1(new_n758), .B2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n757), .A2(KEYINPUT115), .A3(G330), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n936), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n933), .B(new_n1106), .C1(new_n1111), .C2(new_n935), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1111), .A2(new_n935), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1114), .A2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1126), .B1(new_n1128), .B2(new_n934), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n484), .A2(new_n758), .ZN(new_n1130));
  NOR3_X1   g0930(.A1(new_n947), .A2(new_n688), .A3(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1119), .B1(new_n1129), .B2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n722), .B1(new_n1118), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n1135), .B(new_n1119), .C1(new_n1132), .C2(new_n1129), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1118), .A2(new_n768), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n964), .A2(G283), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n1092), .A2(new_n1139), .A3(new_n815), .A4(new_n859), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n274), .B1(new_n862), .B2(G116), .ZN(new_n1141));
  OAI221_X1 g0941(.A(new_n1141), .B1(new_n205), .B2(new_n797), .C1(new_n869), .C2(new_n529), .ZN(new_n1142));
  AOI211_X1 g0942(.A(new_n1140), .B(new_n1142), .C1(G107), .C2(new_n852), .ZN(new_n1143));
  INV_X1    g0943(.A(G125), .ZN(new_n1144));
  OAI221_X1 g0944(.A(new_n274), .B1(new_n202), .B2(new_n786), .C1(new_n869), .C2(new_n1144), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1145), .B(KEYINPUT117), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n814), .A2(G150), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1147), .B(KEYINPUT53), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(KEYINPUT54), .B(G143), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n862), .A2(G132), .B1(new_n856), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(G128), .ZN(new_n1152));
  OAI221_X1 g0952(.A(new_n1151), .B1(new_n1152), .B2(new_n802), .C1(new_n810), .C2(new_n806), .ZN(new_n1153));
  AOI211_X1 g0953(.A(new_n1148), .B(new_n1153), .C1(G137), .C2(new_n852), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1143), .B1(new_n1146), .B2(new_n1154), .ZN(new_n1155));
  OAI221_X1 g0955(.A(new_n769), .B1(new_n450), .B2(new_n844), .C1(new_n1155), .C2(new_n781), .ZN(new_n1156));
  XOR2_X1   g0956(.A(new_n1156), .B(KEYINPUT118), .Z(new_n1157));
  OAI21_X1  g0957(.A(new_n1157), .B1(new_n945), .B2(new_n777), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1137), .A2(new_n1138), .A3(new_n1158), .ZN(G378));
  AND4_X1   g0959(.A1(new_n757), .A2(new_n911), .A3(new_n839), .A4(new_n913), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1160), .B1(new_n895), .B2(new_n938), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n713), .B1(new_n1161), .B2(new_n915), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n299), .A2(new_n694), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1165), .B1(new_n687), .B2(new_n316), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  NOR3_X1   g0967(.A1(new_n687), .A2(new_n316), .A3(new_n1165), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1164), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1168), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1170), .A2(new_n1166), .A3(new_n1163), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1169), .A2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  AND3_X1   g0973(.A1(new_n1162), .A2(new_n917), .A3(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1173), .B1(new_n1162), .B2(new_n917), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n946), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  AND3_X1   g0976(.A1(new_n902), .A2(new_n906), .A3(new_n916), .ZN(new_n1177));
  OAI21_X1  g0977(.A(G330), .B1(new_n925), .B2(KEYINPUT40), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1172), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n945), .A2(new_n941), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1103), .A2(new_n935), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n924), .A2(new_n903), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n1181), .A2(new_n1182), .B1(new_n681), .B2(new_n694), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1180), .A2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1162), .A2(new_n917), .A3(new_n1173), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1179), .A2(new_n1184), .A3(new_n1185), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1176), .A2(KEYINPUT122), .A3(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT122), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n946), .B(new_n1188), .C1(new_n1174), .C2(new_n1175), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n1112), .A2(new_n1113), .B1(new_n935), .B2(new_n1111), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n1190), .A2(new_n1103), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1116), .A2(new_n1191), .A3(new_n1117), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1192), .A2(new_n1131), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1187), .A2(new_n1189), .A3(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT57), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1195), .B1(new_n1176), .B2(new_n1186), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n722), .B1(new_n1197), .B2(new_n1193), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1196), .A2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1187), .A2(new_n768), .A3(new_n1189), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n806), .A2(new_n223), .B1(new_n790), .B2(new_n225), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n274), .A2(G41), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1202), .B1(new_n324), .B2(new_n797), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n1201), .B(new_n1203), .C1(G107), .C2(new_n862), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n786), .A2(new_n426), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n800), .A2(new_n205), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n1205), .B(new_n1206), .C1(G116), .C2(new_n964), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1204), .B(new_n1207), .C1(new_n1064), .C2(new_n869), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(new_n1208), .B(KEYINPUT119), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT58), .ZN(new_n1210));
  AND2_X1   g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(G33), .A2(G41), .ZN(new_n1212));
  NOR3_X1   g1012(.A1(new_n1202), .A2(G50), .A3(new_n1212), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n1144), .A2(new_n802), .B1(new_n800), .B2(new_n868), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(G150), .B2(new_n807), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n862), .A2(G128), .B1(new_n856), .B2(G137), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n1215), .B(new_n1216), .C1(new_n790), .C2(new_n1149), .ZN(new_n1217));
  OR2_X1    g1017(.A1(new_n1217), .A2(KEYINPUT59), .ZN(new_n1218));
  INV_X1    g1018(.A(G124), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n1212), .B1(new_n784), .B2(new_n1219), .C1(new_n810), .C2(new_n786), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(new_n1217), .B2(KEYINPUT59), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1213), .B1(new_n1218), .B2(new_n1221), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1222), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n780), .B1(new_n1211), .B2(new_n1223), .ZN(new_n1224));
  XNOR2_X1  g1024(.A(new_n1224), .B(KEYINPUT120), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n770), .B1(new_n202), .B2(new_n843), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n1225), .B(new_n1226), .C1(new_n1172), .C2(new_n777), .ZN(new_n1227));
  XNOR2_X1  g1027(.A(new_n1227), .B(KEYINPUT121), .ZN(new_n1228));
  AND2_X1   g1028(.A1(new_n1200), .A2(new_n1228), .ZN(new_n1229));
  AND2_X1   g1029(.A1(new_n1199), .A2(new_n1229), .ZN(new_n1230));
  AND2_X1   g1030(.A1(new_n1230), .A2(KEYINPUT123), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1230), .A2(KEYINPUT123), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1231), .A2(new_n1232), .ZN(G375));
  NOR2_X1   g1033(.A1(new_n1129), .A2(new_n1132), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1191), .A2(new_n1131), .ZN(new_n1235));
  OR3_X1    g1035(.A1(new_n1234), .A2(new_n1235), .A3(new_n1015), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n935), .A2(new_n776), .ZN(new_n1237));
  XOR2_X1   g1037(.A(new_n1237), .B(KEYINPUT124), .Z(new_n1238));
  OAI21_X1  g1038(.A(new_n769), .B1(G68), .B2(new_n844), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT125), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n274), .B1(new_n787), .B2(G77), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(new_n852), .A2(G116), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n785), .A2(G303), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n795), .A2(new_n1064), .B1(new_n797), .B2(new_n206), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n802), .A2(new_n529), .B1(new_n790), .B2(new_n205), .ZN(new_n1245));
  AOI211_X1 g1045(.A(new_n1244), .B(new_n1245), .C1(new_n323), .C2(new_n807), .ZN(new_n1246));
  OR2_X1    g1046(.A1(new_n1241), .A2(new_n1240), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1242), .A2(new_n1243), .A3(new_n1246), .A4(new_n1247), .ZN(new_n1248));
  OAI22_X1  g1048(.A1(new_n795), .A2(new_n864), .B1(new_n802), .B2(new_n868), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1249), .B1(new_n852), .B2(new_n1150), .ZN(new_n1250));
  XOR2_X1   g1050(.A(new_n1250), .B(KEYINPUT126), .Z(new_n1251));
  AOI211_X1 g1051(.A(new_n331), .B(new_n1205), .C1(G150), .C2(new_n856), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n807), .A2(G50), .B1(new_n814), .B2(G159), .ZN(new_n1253));
  OAI211_X1 g1053(.A(new_n1252), .B(new_n1253), .C1(new_n1152), .C2(new_n869), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1248), .B1(new_n1251), .B2(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1239), .B1(new_n1255), .B2(new_n780), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(new_n1191), .A2(new_n768), .B1(new_n1238), .B2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1236), .A2(new_n1257), .ZN(G381));
  NOR4_X1   g1058(.A1(G390), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1138), .A2(new_n1158), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1260), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1259), .A2(new_n1261), .A3(new_n1257), .A4(new_n1236), .ZN(new_n1262));
  OR3_X1    g1062(.A1(G375), .A2(G387), .A3(new_n1262), .ZN(G407));
  OAI21_X1  g1063(.A(new_n1261), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1264));
  OAI211_X1 g1064(.A(G407), .B(G213), .C1(G343), .C2(new_n1264), .ZN(G409));
  XNOR2_X1  g1065(.A(G393), .B(new_n830), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(KEYINPUT110), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1268));
  AOI211_X1 g1068(.A(new_n986), .B(new_n1015), .C1(new_n1022), .C2(new_n763), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n767), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(new_n1038), .ZN(new_n1271));
  AOI21_X1  g1071(.A(G390), .B1(new_n1271), .B2(new_n985), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n985), .ZN(new_n1273));
  AOI211_X1 g1073(.A(new_n1273), .B(new_n1101), .C1(new_n1270), .C2(new_n1038), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1267), .B1(new_n1272), .B2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(G387), .A2(new_n1101), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1271), .A2(new_n985), .A3(G390), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1276), .A2(new_n1266), .A3(new_n1277), .ZN(new_n1278));
  AND2_X1   g1078(.A1(new_n1275), .A2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT61), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n695), .A2(G213), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1199), .A2(G378), .A3(new_n1229), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1176), .A2(new_n1186), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(new_n768), .ZN(new_n1285));
  OAI211_X1 g1085(.A(new_n1228), .B(new_n1285), .C1(new_n1194), .C2(new_n1015), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(new_n1261), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1282), .B1(new_n1283), .B2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1191), .A2(new_n1131), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1235), .B1(KEYINPUT60), .B2(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1129), .A2(new_n1132), .A3(KEYINPUT60), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(new_n721), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1257), .B1(new_n1290), .B2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(new_n875), .ZN(new_n1294));
  OAI211_X1 g1094(.A(G384), .B(new_n1257), .C1(new_n1290), .C2(new_n1292), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1296), .A2(G2897), .A3(new_n1282), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1282), .A2(G2897), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1294), .A2(new_n1295), .A3(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1297), .A2(new_n1299), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1280), .B1(new_n1288), .B2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT62), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1296), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1302), .B1(new_n1288), .B2(new_n1303), .ZN(new_n1304));
  NOR2_X1   g1104(.A1(new_n1301), .A2(new_n1304), .ZN(new_n1305));
  AOI211_X1 g1105(.A(new_n1282), .B(new_n1296), .C1(new_n1283), .C2(new_n1287), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(new_n1302), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1279), .B1(new_n1305), .B2(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1288), .A2(KEYINPUT63), .A3(new_n1303), .ZN(new_n1309));
  OAI211_X1 g1109(.A(new_n1309), .B(new_n1280), .C1(new_n1288), .C2(new_n1300), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1279), .B1(new_n1306), .B2(KEYINPUT63), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  OAI21_X1  g1112(.A(KEYINPUT127), .B1(new_n1308), .B2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT127), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1275), .A2(new_n1278), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1288), .A2(new_n1303), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT63), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1315), .B1(new_n1316), .B2(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1301), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1318), .A2(new_n1319), .A3(new_n1309), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(new_n1316), .A2(KEYINPUT62), .ZN(new_n1321));
  NOR3_X1   g1121(.A1(new_n1321), .A2(new_n1301), .A3(new_n1304), .ZN(new_n1322));
  OAI211_X1 g1122(.A(new_n1314), .B(new_n1320), .C1(new_n1322), .C2(new_n1279), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1313), .A2(new_n1323), .ZN(G405));
  XNOR2_X1  g1124(.A(new_n1315), .B(new_n1296), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1264), .B1(new_n1261), .B2(new_n1230), .ZN(new_n1326));
  XNOR2_X1  g1126(.A(new_n1325), .B(new_n1326), .ZN(G402));
endmodule


