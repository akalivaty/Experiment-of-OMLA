

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591;

  XNOR2_X1 U327 ( .A(n366), .B(n365), .ZN(n561) );
  XNOR2_X1 U328 ( .A(n384), .B(KEYINPUT65), .ZN(n385) );
  XNOR2_X1 U329 ( .A(n386), .B(n385), .ZN(n387) );
  INV_X1 U330 ( .A(n407), .ZN(n354) );
  XNOR2_X1 U331 ( .A(KEYINPUT121), .B(KEYINPUT54), .ZN(n413) );
  XNOR2_X1 U332 ( .A(n355), .B(n354), .ZN(n356) );
  XNOR2_X1 U333 ( .A(n414), .B(n413), .ZN(n573) );
  XNOR2_X1 U334 ( .A(n357), .B(n356), .ZN(n361) );
  NOR2_X1 U335 ( .A1(n501), .A2(n458), .ZN(n570) );
  XOR2_X1 U336 ( .A(n310), .B(n309), .Z(n535) );
  XNOR2_X1 U337 ( .A(n459), .B(G190GAT), .ZN(n460) );
  XNOR2_X1 U338 ( .A(n461), .B(n460), .ZN(G1351GAT) );
  XOR2_X1 U339 ( .A(G43GAT), .B(G134GAT), .Z(n350) );
  XNOR2_X1 U340 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n295) );
  XNOR2_X1 U341 ( .A(n295), .B(KEYINPUT81), .ZN(n450) );
  XNOR2_X1 U342 ( .A(n350), .B(n450), .ZN(n296) );
  XOR2_X1 U343 ( .A(G15GAT), .B(G127GAT), .Z(n373) );
  XNOR2_X1 U344 ( .A(n296), .B(n373), .ZN(n301) );
  XNOR2_X1 U345 ( .A(G99GAT), .B(G71GAT), .ZN(n297) );
  XNOR2_X1 U346 ( .A(n297), .B(G120GAT), .ZN(n323) );
  XOR2_X1 U347 ( .A(n323), .B(KEYINPUT20), .Z(n299) );
  NAND2_X1 U348 ( .A1(G227GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U349 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U350 ( .A(n301), .B(n300), .Z(n310) );
  XNOR2_X1 U351 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n302) );
  XNOR2_X1 U352 ( .A(n302), .B(KEYINPUT17), .ZN(n303) );
  XOR2_X1 U353 ( .A(n303), .B(KEYINPUT82), .Z(n305) );
  XNOR2_X1 U354 ( .A(G169GAT), .B(G183GAT), .ZN(n304) );
  XNOR2_X1 U355 ( .A(n305), .B(n304), .ZN(n403) );
  XOR2_X1 U356 ( .A(KEYINPUT84), .B(G176GAT), .Z(n307) );
  XNOR2_X1 U357 ( .A(G190GAT), .B(KEYINPUT83), .ZN(n306) );
  XNOR2_X1 U358 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U359 ( .A(n403), .B(n308), .ZN(n309) );
  INV_X1 U360 ( .A(n535), .ZN(n501) );
  XOR2_X1 U361 ( .A(KEYINPUT71), .B(KEYINPUT32), .Z(n312) );
  XNOR2_X1 U362 ( .A(KEYINPUT13), .B(KEYINPUT73), .ZN(n311) );
  XNOR2_X1 U363 ( .A(n312), .B(n311), .ZN(n327) );
  XOR2_X1 U364 ( .A(G85GAT), .B(G57GAT), .Z(n434) );
  XOR2_X1 U365 ( .A(G64GAT), .B(G92GAT), .Z(n314) );
  XNOR2_X1 U366 ( .A(G176GAT), .B(G204GAT), .ZN(n313) );
  XNOR2_X1 U367 ( .A(n314), .B(n313), .ZN(n401) );
  XOR2_X1 U368 ( .A(n434), .B(n401), .Z(n316) );
  NAND2_X1 U369 ( .A1(G230GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U370 ( .A(n316), .B(n315), .ZN(n320) );
  XOR2_X1 U371 ( .A(KEYINPUT31), .B(KEYINPUT70), .Z(n318) );
  XNOR2_X1 U372 ( .A(KEYINPUT33), .B(KEYINPUT74), .ZN(n317) );
  XNOR2_X1 U373 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U374 ( .A(n320), .B(n319), .Z(n325) );
  XOR2_X1 U375 ( .A(G78GAT), .B(G148GAT), .Z(n322) );
  XNOR2_X1 U376 ( .A(G106GAT), .B(KEYINPUT72), .ZN(n321) );
  XNOR2_X1 U377 ( .A(n322), .B(n321), .ZN(n429) );
  XNOR2_X1 U378 ( .A(n323), .B(n429), .ZN(n324) );
  XNOR2_X1 U379 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U380 ( .A(n327), .B(n326), .ZN(n580) );
  XOR2_X1 U381 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n329) );
  XNOR2_X1 U382 ( .A(G1GAT), .B(KEYINPUT67), .ZN(n328) );
  XNOR2_X1 U383 ( .A(n329), .B(n328), .ZN(n337) );
  XOR2_X1 U384 ( .A(KEYINPUT68), .B(KEYINPUT69), .Z(n335) );
  XOR2_X1 U385 ( .A(G8GAT), .B(G197GAT), .Z(n331) );
  XNOR2_X1 U386 ( .A(G141GAT), .B(G22GAT), .ZN(n330) );
  XNOR2_X1 U387 ( .A(n331), .B(n330), .ZN(n333) );
  XNOR2_X1 U388 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n332) );
  XNOR2_X1 U389 ( .A(n332), .B(KEYINPUT7), .ZN(n353) );
  XNOR2_X1 U390 ( .A(n333), .B(n353), .ZN(n334) );
  XNOR2_X1 U391 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U392 ( .A(n337), .B(n336), .ZN(n345) );
  NAND2_X1 U393 ( .A1(G229GAT), .A2(G233GAT), .ZN(n343) );
  XOR2_X1 U394 ( .A(G15GAT), .B(G113GAT), .Z(n339) );
  XNOR2_X1 U395 ( .A(G169GAT), .B(G43GAT), .ZN(n338) );
  XNOR2_X1 U396 ( .A(n339), .B(n338), .ZN(n341) );
  XOR2_X1 U397 ( .A(G50GAT), .B(G36GAT), .Z(n340) );
  XNOR2_X1 U398 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U399 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U400 ( .A(n345), .B(n344), .Z(n508) );
  INV_X1 U401 ( .A(n508), .ZN(n576) );
  XOR2_X1 U402 ( .A(KEYINPUT77), .B(KEYINPUT64), .Z(n347) );
  XNOR2_X1 U403 ( .A(G85GAT), .B(KEYINPUT66), .ZN(n346) );
  XNOR2_X1 U404 ( .A(n347), .B(n346), .ZN(n349) );
  INV_X1 U405 ( .A(G92GAT), .ZN(n348) );
  XNOR2_X1 U406 ( .A(n349), .B(n348), .ZN(n352) );
  XNOR2_X1 U407 ( .A(n350), .B(G218GAT), .ZN(n351) );
  XNOR2_X1 U408 ( .A(n352), .B(n351), .ZN(n357) );
  XOR2_X1 U409 ( .A(G50GAT), .B(G162GAT), .Z(n416) );
  XNOR2_X1 U410 ( .A(n353), .B(n416), .ZN(n355) );
  XOR2_X1 U411 ( .A(G36GAT), .B(G190GAT), .Z(n407) );
  XOR2_X1 U412 ( .A(KEYINPUT11), .B(G106GAT), .Z(n359) );
  NAND2_X1 U413 ( .A1(G232GAT), .A2(G233GAT), .ZN(n358) );
  XNOR2_X1 U414 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U415 ( .A(n361), .B(n360), .ZN(n366) );
  XOR2_X1 U416 ( .A(KEYINPUT9), .B(KEYINPUT10), .Z(n363) );
  XNOR2_X1 U417 ( .A(KEYINPUT75), .B(KEYINPUT76), .ZN(n362) );
  XNOR2_X1 U418 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U419 ( .A(G99GAT), .B(n364), .ZN(n365) );
  XOR2_X1 U420 ( .A(KEYINPUT36), .B(n561), .Z(n588) );
  XOR2_X1 U421 ( .A(G8GAT), .B(KEYINPUT78), .Z(n402) );
  XOR2_X1 U422 ( .A(G22GAT), .B(G155GAT), .Z(n420) );
  XOR2_X1 U423 ( .A(n402), .B(n420), .Z(n368) );
  XNOR2_X1 U424 ( .A(G183GAT), .B(G71GAT), .ZN(n367) );
  XNOR2_X1 U425 ( .A(n368), .B(n367), .ZN(n372) );
  XOR2_X1 U426 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n370) );
  NAND2_X1 U427 ( .A1(G231GAT), .A2(G233GAT), .ZN(n369) );
  XNOR2_X1 U428 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U429 ( .A(n372), .B(n371), .Z(n375) );
  XNOR2_X1 U430 ( .A(n373), .B(KEYINPUT79), .ZN(n374) );
  XNOR2_X1 U431 ( .A(n375), .B(n374), .ZN(n383) );
  XOR2_X1 U432 ( .A(KEYINPUT13), .B(G64GAT), .Z(n377) );
  XNOR2_X1 U433 ( .A(G78GAT), .B(G211GAT), .ZN(n376) );
  XNOR2_X1 U434 ( .A(n377), .B(n376), .ZN(n381) );
  XOR2_X1 U435 ( .A(G57GAT), .B(KEYINPUT15), .Z(n379) );
  XNOR2_X1 U436 ( .A(G1GAT), .B(KEYINPUT80), .ZN(n378) );
  XNOR2_X1 U437 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U438 ( .A(n381), .B(n380), .Z(n382) );
  XOR2_X1 U439 ( .A(n383), .B(n382), .Z(n584) );
  INV_X1 U440 ( .A(n584), .ZN(n477) );
  OR2_X1 U441 ( .A1(n588), .A2(n477), .ZN(n386) );
  INV_X1 U442 ( .A(KEYINPUT45), .ZN(n384) );
  NOR2_X1 U443 ( .A1(n576), .A2(n387), .ZN(n388) );
  NAND2_X1 U444 ( .A1(n580), .A2(n388), .ZN(n397) );
  XNOR2_X1 U445 ( .A(KEYINPUT41), .B(n580), .ZN(n553) );
  NAND2_X1 U446 ( .A1(n553), .A2(n576), .ZN(n389) );
  XNOR2_X1 U447 ( .A(n389), .B(KEYINPUT46), .ZN(n390) );
  NAND2_X1 U448 ( .A1(n390), .A2(n477), .ZN(n391) );
  XNOR2_X1 U449 ( .A(KEYINPUT113), .B(n391), .ZN(n393) );
  INV_X1 U450 ( .A(n561), .ZN(n392) );
  NAND2_X1 U451 ( .A1(n393), .A2(n392), .ZN(n395) );
  XOR2_X1 U452 ( .A(KEYINPUT47), .B(KEYINPUT114), .Z(n394) );
  XNOR2_X1 U453 ( .A(n395), .B(n394), .ZN(n396) );
  NAND2_X1 U454 ( .A1(n397), .A2(n396), .ZN(n398) );
  XNOR2_X1 U455 ( .A(n398), .B(KEYINPUT48), .ZN(n549) );
  XOR2_X1 U456 ( .A(G211GAT), .B(KEYINPUT21), .Z(n400) );
  XNOR2_X1 U457 ( .A(G197GAT), .B(G218GAT), .ZN(n399) );
  XNOR2_X1 U458 ( .A(n400), .B(n399), .ZN(n415) );
  XOR2_X1 U459 ( .A(n415), .B(n401), .Z(n411) );
  XOR2_X1 U460 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n405) );
  XNOR2_X1 U461 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U462 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U463 ( .A(n407), .B(n406), .Z(n409) );
  NAND2_X1 U464 ( .A1(G226GAT), .A2(G233GAT), .ZN(n408) );
  XNOR2_X1 U465 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U466 ( .A(n411), .B(n410), .ZN(n465) );
  INV_X1 U467 ( .A(n465), .ZN(n527) );
  INV_X1 U468 ( .A(n527), .ZN(n499) );
  XOR2_X1 U469 ( .A(KEYINPUT120), .B(n499), .Z(n412) );
  NAND2_X1 U470 ( .A1(n549), .A2(n412), .ZN(n414) );
  XOR2_X1 U471 ( .A(n416), .B(n415), .Z(n418) );
  NAND2_X1 U472 ( .A1(G228GAT), .A2(G233GAT), .ZN(n417) );
  XNOR2_X1 U473 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U474 ( .A(n419), .B(G204GAT), .Z(n422) );
  XNOR2_X1 U475 ( .A(n420), .B(KEYINPUT86), .ZN(n421) );
  XNOR2_X1 U476 ( .A(n422), .B(n421), .ZN(n426) );
  XOR2_X1 U477 ( .A(KEYINPUT22), .B(KEYINPUT88), .Z(n424) );
  XNOR2_X1 U478 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n423) );
  XNOR2_X1 U479 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U480 ( .A(n426), .B(n425), .ZN(n431) );
  XOR2_X1 U481 ( .A(KEYINPUT2), .B(KEYINPUT87), .Z(n428) );
  XNOR2_X1 U482 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n427) );
  XNOR2_X1 U483 ( .A(n428), .B(n427), .ZN(n449) );
  XOR2_X1 U484 ( .A(n449), .B(n429), .Z(n430) );
  XNOR2_X1 U485 ( .A(n431), .B(n430), .ZN(n469) );
  XOR2_X1 U486 ( .A(G148GAT), .B(G127GAT), .Z(n433) );
  XNOR2_X1 U487 ( .A(G120GAT), .B(G134GAT), .ZN(n432) );
  XNOR2_X1 U488 ( .A(n433), .B(n432), .ZN(n435) );
  XOR2_X1 U489 ( .A(n435), .B(n434), .Z(n437) );
  XNOR2_X1 U490 ( .A(G29GAT), .B(G162GAT), .ZN(n436) );
  XNOR2_X1 U491 ( .A(n437), .B(n436), .ZN(n441) );
  XOR2_X1 U492 ( .A(KEYINPUT1), .B(KEYINPUT92), .Z(n439) );
  XNOR2_X1 U493 ( .A(KEYINPUT93), .B(KEYINPUT89), .ZN(n438) );
  XNOR2_X1 U494 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U495 ( .A(n441), .B(n440), .ZN(n445) );
  XOR2_X1 U496 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n443) );
  XNOR2_X1 U497 ( .A(G1GAT), .B(G155GAT), .ZN(n442) );
  XNOR2_X1 U498 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U499 ( .A(n445), .B(n444), .ZN(n454) );
  XOR2_X1 U500 ( .A(KEYINPUT90), .B(KEYINPUT91), .Z(n447) );
  NAND2_X1 U501 ( .A1(G225GAT), .A2(G233GAT), .ZN(n446) );
  XNOR2_X1 U502 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U503 ( .A(n448), .B(KEYINPUT6), .Z(n452) );
  XNOR2_X1 U504 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U505 ( .A(n452), .B(n451), .ZN(n453) );
  XOR2_X1 U506 ( .A(n454), .B(n453), .Z(n524) );
  NOR2_X1 U507 ( .A1(n469), .A2(n524), .ZN(n455) );
  AND2_X1 U508 ( .A1(n573), .A2(n455), .ZN(n457) );
  XNOR2_X1 U509 ( .A(KEYINPUT55), .B(KEYINPUT122), .ZN(n456) );
  XNOR2_X1 U510 ( .A(n457), .B(n456), .ZN(n458) );
  NAND2_X1 U511 ( .A1(n570), .A2(n561), .ZN(n461) );
  XOR2_X1 U512 ( .A(KEYINPUT125), .B(KEYINPUT58), .Z(n459) );
  XNOR2_X1 U513 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n483) );
  XNOR2_X1 U514 ( .A(n469), .B(KEYINPUT28), .ZN(n530) );
  INV_X1 U515 ( .A(n530), .ZN(n505) );
  INV_X1 U516 ( .A(n524), .ZN(n572) );
  XNOR2_X1 U517 ( .A(n465), .B(KEYINPUT27), .ZN(n471) );
  NOR2_X1 U518 ( .A1(n572), .A2(n471), .ZN(n462) );
  XNOR2_X1 U519 ( .A(n462), .B(KEYINPUT96), .ZN(n548) );
  NAND2_X1 U520 ( .A1(n505), .A2(n548), .ZN(n537) );
  XOR2_X1 U521 ( .A(KEYINPUT85), .B(n535), .Z(n463) );
  NOR2_X1 U522 ( .A1(n537), .A2(n463), .ZN(n476) );
  XNOR2_X1 U523 ( .A(KEYINPUT25), .B(KEYINPUT98), .ZN(n464) );
  XNOR2_X1 U524 ( .A(n464), .B(KEYINPUT97), .ZN(n468) );
  NOR2_X1 U525 ( .A1(n501), .A2(n465), .ZN(n466) );
  NOR2_X1 U526 ( .A1(n469), .A2(n466), .ZN(n467) );
  XNOR2_X1 U527 ( .A(n468), .B(n467), .ZN(n473) );
  NAND2_X1 U528 ( .A1(n469), .A2(n501), .ZN(n470) );
  XNOR2_X1 U529 ( .A(n470), .B(KEYINPUT26), .ZN(n575) );
  NOR2_X1 U530 ( .A1(n575), .A2(n471), .ZN(n472) );
  NOR2_X1 U531 ( .A1(n473), .A2(n472), .ZN(n474) );
  NOR2_X1 U532 ( .A1(n524), .A2(n474), .ZN(n475) );
  NOR2_X1 U533 ( .A1(n476), .A2(n475), .ZN(n490) );
  NOR2_X1 U534 ( .A1(n561), .A2(n477), .ZN(n478) );
  XOR2_X1 U535 ( .A(KEYINPUT16), .B(n478), .Z(n479) );
  NOR2_X1 U536 ( .A1(n490), .A2(n479), .ZN(n480) );
  XNOR2_X1 U537 ( .A(KEYINPUT99), .B(n480), .ZN(n509) );
  NAND2_X1 U538 ( .A1(n576), .A2(n580), .ZN(n494) );
  NOR2_X1 U539 ( .A1(n509), .A2(n494), .ZN(n481) );
  XNOR2_X1 U540 ( .A(n481), .B(KEYINPUT100), .ZN(n487) );
  NAND2_X1 U541 ( .A1(n524), .A2(n487), .ZN(n482) );
  XNOR2_X1 U542 ( .A(n483), .B(n482), .ZN(G1324GAT) );
  NAND2_X1 U543 ( .A1(n487), .A2(n527), .ZN(n484) );
  XNOR2_X1 U544 ( .A(n484), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U545 ( .A(G15GAT), .B(KEYINPUT35), .Z(n486) );
  NAND2_X1 U546 ( .A1(n487), .A2(n535), .ZN(n485) );
  XNOR2_X1 U547 ( .A(n486), .B(n485), .ZN(G1326GAT) );
  XOR2_X1 U548 ( .A(G22GAT), .B(KEYINPUT101), .Z(n489) );
  NAND2_X1 U549 ( .A1(n487), .A2(n530), .ZN(n488) );
  XNOR2_X1 U550 ( .A(n489), .B(n488), .ZN(G1327GAT) );
  NOR2_X1 U551 ( .A1(n584), .A2(n490), .ZN(n491) );
  XOR2_X1 U552 ( .A(KEYINPUT102), .B(n491), .Z(n492) );
  NOR2_X1 U553 ( .A1(n588), .A2(n492), .ZN(n493) );
  XNOR2_X1 U554 ( .A(KEYINPUT37), .B(n493), .ZN(n521) );
  NOR2_X1 U555 ( .A1(n521), .A2(n494), .ZN(n495) );
  XOR2_X1 U556 ( .A(KEYINPUT38), .B(n495), .Z(n504) );
  NOR2_X1 U557 ( .A1(n504), .A2(n572), .ZN(n498) );
  XOR2_X1 U558 ( .A(G29GAT), .B(KEYINPUT39), .Z(n496) );
  XNOR2_X1 U559 ( .A(KEYINPUT103), .B(n496), .ZN(n497) );
  XNOR2_X1 U560 ( .A(n498), .B(n497), .ZN(G1328GAT) );
  NOR2_X1 U561 ( .A1(n504), .A2(n499), .ZN(n500) );
  XOR2_X1 U562 ( .A(G36GAT), .B(n500), .Z(G1329GAT) );
  NOR2_X1 U563 ( .A1(n501), .A2(n504), .ZN(n502) );
  XOR2_X1 U564 ( .A(KEYINPUT40), .B(n502), .Z(n503) );
  XNOR2_X1 U565 ( .A(G43GAT), .B(n503), .ZN(G1330GAT) );
  NOR2_X1 U566 ( .A1(n505), .A2(n504), .ZN(n506) );
  XOR2_X1 U567 ( .A(KEYINPUT104), .B(n506), .Z(n507) );
  XNOR2_X1 U568 ( .A(G50GAT), .B(n507), .ZN(G1331GAT) );
  XOR2_X1 U569 ( .A(KEYINPUT42), .B(KEYINPUT107), .Z(n512) );
  XOR2_X1 U570 ( .A(n553), .B(KEYINPUT105), .Z(n567) );
  NAND2_X1 U571 ( .A1(n508), .A2(n567), .ZN(n522) );
  NOR2_X1 U572 ( .A1(n509), .A2(n522), .ZN(n510) );
  XNOR2_X1 U573 ( .A(n510), .B(KEYINPUT106), .ZN(n518) );
  NAND2_X1 U574 ( .A1(n524), .A2(n518), .ZN(n511) );
  XNOR2_X1 U575 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U576 ( .A(G57GAT), .B(n513), .ZN(G1332GAT) );
  NAND2_X1 U577 ( .A1(n518), .A2(n527), .ZN(n514) );
  XNOR2_X1 U578 ( .A(n514), .B(KEYINPUT108), .ZN(n515) );
  XNOR2_X1 U579 ( .A(G64GAT), .B(n515), .ZN(G1333GAT) );
  XOR2_X1 U580 ( .A(G71GAT), .B(KEYINPUT109), .Z(n517) );
  NAND2_X1 U581 ( .A1(n518), .A2(n535), .ZN(n516) );
  XNOR2_X1 U582 ( .A(n517), .B(n516), .ZN(G1334GAT) );
  XOR2_X1 U583 ( .A(G78GAT), .B(KEYINPUT43), .Z(n520) );
  NAND2_X1 U584 ( .A1(n518), .A2(n530), .ZN(n519) );
  XNOR2_X1 U585 ( .A(n520), .B(n519), .ZN(G1335GAT) );
  XOR2_X1 U586 ( .A(G85GAT), .B(KEYINPUT111), .Z(n526) );
  NOR2_X1 U587 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U588 ( .A(n523), .B(KEYINPUT110), .ZN(n531) );
  NAND2_X1 U589 ( .A1(n524), .A2(n531), .ZN(n525) );
  XNOR2_X1 U590 ( .A(n526), .B(n525), .ZN(G1336GAT) );
  NAND2_X1 U591 ( .A1(n531), .A2(n527), .ZN(n528) );
  XNOR2_X1 U592 ( .A(n528), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U593 ( .A1(n535), .A2(n531), .ZN(n529) );
  XNOR2_X1 U594 ( .A(G99GAT), .B(n529), .ZN(G1338GAT) );
  XOR2_X1 U595 ( .A(KEYINPUT112), .B(KEYINPUT44), .Z(n533) );
  NAND2_X1 U596 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U597 ( .A(n533), .B(n532), .ZN(n534) );
  XOR2_X1 U598 ( .A(G106GAT), .B(n534), .Z(G1339GAT) );
  XOR2_X1 U599 ( .A(G113GAT), .B(KEYINPUT115), .Z(n539) );
  NAND2_X1 U600 ( .A1(n549), .A2(n535), .ZN(n536) );
  NOR2_X1 U601 ( .A1(n537), .A2(n536), .ZN(n545) );
  NAND2_X1 U602 ( .A1(n545), .A2(n576), .ZN(n538) );
  XNOR2_X1 U603 ( .A(n539), .B(n538), .ZN(G1340GAT) );
  XOR2_X1 U604 ( .A(G120GAT), .B(KEYINPUT49), .Z(n541) );
  NAND2_X1 U605 ( .A1(n545), .A2(n567), .ZN(n540) );
  XNOR2_X1 U606 ( .A(n541), .B(n540), .ZN(G1341GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n543) );
  NAND2_X1 U608 ( .A1(n545), .A2(n584), .ZN(n542) );
  XNOR2_X1 U609 ( .A(n543), .B(n542), .ZN(n544) );
  XOR2_X1 U610 ( .A(G127GAT), .B(n544), .Z(G1342GAT) );
  XOR2_X1 U611 ( .A(G134GAT), .B(KEYINPUT51), .Z(n547) );
  NAND2_X1 U612 ( .A1(n545), .A2(n561), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n547), .B(n546), .ZN(G1343GAT) );
  XOR2_X1 U614 ( .A(G141GAT), .B(KEYINPUT117), .Z(n552) );
  NAND2_X1 U615 ( .A1(n549), .A2(n548), .ZN(n550) );
  NOR2_X1 U616 ( .A1(n575), .A2(n550), .ZN(n560) );
  NAND2_X1 U617 ( .A1(n560), .A2(n576), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n552), .B(n551), .ZN(G1344GAT) );
  XNOR2_X1 U619 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n557) );
  XOR2_X1 U620 ( .A(KEYINPUT118), .B(KEYINPUT53), .Z(n555) );
  NAND2_X1 U621 ( .A1(n560), .A2(n553), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n557), .B(n556), .ZN(G1345GAT) );
  XOR2_X1 U624 ( .A(G155GAT), .B(KEYINPUT119), .Z(n559) );
  NAND2_X1 U625 ( .A1(n560), .A2(n584), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(G1346GAT) );
  NAND2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U629 ( .A1(n570), .A2(n576), .ZN(n563) );
  XNOR2_X1 U630 ( .A(G169GAT), .B(n563), .ZN(G1348GAT) );
  XOR2_X1 U631 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n565) );
  XNOR2_X1 U632 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n564) );
  XNOR2_X1 U633 ( .A(n565), .B(n564), .ZN(n566) );
  XOR2_X1 U634 ( .A(KEYINPUT56), .B(n566), .Z(n569) );
  NAND2_X1 U635 ( .A1(n567), .A2(n570), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n569), .B(n568), .ZN(G1349GAT) );
  NAND2_X1 U637 ( .A1(n570), .A2(n584), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n571), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U639 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n578) );
  NAND2_X1 U640 ( .A1(n573), .A2(n572), .ZN(n574) );
  NOR2_X1 U641 ( .A1(n575), .A2(n574), .ZN(n585) );
  NAND2_X1 U642 ( .A1(n585), .A2(n576), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U644 ( .A(G197GAT), .B(n579), .ZN(G1352GAT) );
  XOR2_X1 U645 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n582) );
  INV_X1 U646 ( .A(n585), .ZN(n587) );
  OR2_X1 U647 ( .A1(n587), .A2(n580), .ZN(n581) );
  XNOR2_X1 U648 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U649 ( .A(G204GAT), .B(n583), .ZN(G1353GAT) );
  NAND2_X1 U650 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n586), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U652 ( .A1(n588), .A2(n587), .ZN(n590) );
  XNOR2_X1 U653 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n589) );
  XNOR2_X1 U654 ( .A(n590), .B(n589), .ZN(n591) );
  XNOR2_X1 U655 ( .A(G218GAT), .B(n591), .ZN(G1355GAT) );
endmodule

