

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U555 ( .A(n671), .B(n670), .ZN(n673) );
  NOR2_X1 U556 ( .A1(n742), .A2(n741), .ZN(n744) );
  NOR2_X1 U557 ( .A1(n804), .A2(n696), .ZN(n697) );
  XNOR2_X1 U558 ( .A(n774), .B(KEYINPUT100), .ZN(n776) );
  XNOR2_X1 U559 ( .A(G299), .B(G290), .ZN(n674) );
  XOR2_X1 U560 ( .A(KEYINPUT96), .B(KEYINPUT30), .Z(n521) );
  NOR2_X1 U561 ( .A1(n980), .A2(n705), .ZN(n711) );
  INV_X1 U562 ( .A(KEYINPUT31), .ZN(n737) );
  XNOR2_X1 U563 ( .A(n738), .B(n737), .ZN(n739) );
  INV_X1 U564 ( .A(KEYINPUT97), .ZN(n743) );
  XNOR2_X1 U565 ( .A(n748), .B(KEYINPUT98), .ZN(n782) );
  XNOR2_X1 U566 ( .A(n679), .B(KEYINPUT19), .ZN(n670) );
  INV_X1 U567 ( .A(n1002), .ZN(n775) );
  NAND2_X1 U568 ( .A1(G8), .A2(n749), .ZN(n786) );
  AND2_X1 U569 ( .A1(n776), .A2(n775), .ZN(n777) );
  XNOR2_X1 U570 ( .A(n675), .B(n674), .ZN(n898) );
  AND2_X1 U571 ( .A1(G2104), .A2(G2105), .ZN(n884) );
  XNOR2_X1 U572 ( .A(n899), .B(G286), .ZN(n900) );
  XOR2_X1 U573 ( .A(KEYINPUT65), .B(n536), .Z(n661) );
  AND2_X1 U574 ( .A1(n842), .A2(n841), .ZN(n843) );
  XNOR2_X1 U575 ( .A(n901), .B(n900), .ZN(n902) );
  NAND2_X1 U576 ( .A1(n884), .A2(G114), .ZN(n522) );
  XNOR2_X1 U577 ( .A(n522), .B(KEYINPUT88), .ZN(n525) );
  INV_X1 U578 ( .A(G2105), .ZN(n527) );
  AND2_X1 U579 ( .A1(G2104), .A2(n527), .ZN(n523) );
  XNOR2_X1 U580 ( .A(n523), .B(KEYINPUT66), .ZN(n629) );
  NAND2_X1 U581 ( .A1(G102), .A2(n629), .ZN(n524) );
  NAND2_X1 U582 ( .A1(n525), .A2(n524), .ZN(n531) );
  NOR2_X1 U583 ( .A1(G2104), .A2(G2105), .ZN(n526) );
  XOR2_X1 U584 ( .A(KEYINPUT17), .B(n526), .Z(n589) );
  NAND2_X1 U585 ( .A1(G138), .A2(n589), .ZN(n529) );
  NOR2_X1 U586 ( .A1(G2104), .A2(n527), .ZN(n885) );
  NAND2_X1 U587 ( .A1(G126), .A2(n885), .ZN(n528) );
  NAND2_X1 U588 ( .A1(n529), .A2(n528), .ZN(n530) );
  NOR2_X1 U589 ( .A1(n531), .A2(n530), .ZN(G164) );
  NOR2_X1 U590 ( .A1(G651), .A2(G543), .ZN(n652) );
  NAND2_X1 U591 ( .A1(n652), .A2(G89), .ZN(n532) );
  XNOR2_X1 U592 ( .A(n532), .B(KEYINPUT4), .ZN(n534) );
  XOR2_X1 U593 ( .A(G543), .B(KEYINPUT0), .Z(n666) );
  INV_X1 U594 ( .A(G651), .ZN(n538) );
  NOR2_X1 U595 ( .A1(n666), .A2(n538), .ZN(n655) );
  NAND2_X1 U596 ( .A1(G76), .A2(n655), .ZN(n533) );
  NAND2_X1 U597 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U598 ( .A(n535), .B(KEYINPUT5), .ZN(n545) );
  NOR2_X1 U599 ( .A1(G651), .A2(n666), .ZN(n536) );
  NAND2_X1 U600 ( .A1(n661), .A2(G51), .ZN(n537) );
  XNOR2_X1 U601 ( .A(n537), .B(KEYINPUT76), .ZN(n542) );
  NOR2_X1 U602 ( .A1(G543), .A2(n538), .ZN(n540) );
  XNOR2_X1 U603 ( .A(KEYINPUT67), .B(KEYINPUT1), .ZN(n539) );
  XNOR2_X1 U604 ( .A(n540), .B(n539), .ZN(n665) );
  NAND2_X1 U605 ( .A1(G63), .A2(n665), .ZN(n541) );
  NAND2_X1 U606 ( .A1(n542), .A2(n541), .ZN(n543) );
  XOR2_X1 U607 ( .A(KEYINPUT6), .B(n543), .Z(n544) );
  NAND2_X1 U608 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U609 ( .A(n546), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U610 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U611 ( .A1(G65), .A2(n665), .ZN(n548) );
  NAND2_X1 U612 ( .A1(G53), .A2(n661), .ZN(n547) );
  NAND2_X1 U613 ( .A1(n548), .A2(n547), .ZN(n552) );
  NAND2_X1 U614 ( .A1(G91), .A2(n652), .ZN(n550) );
  NAND2_X1 U615 ( .A1(G78), .A2(n655), .ZN(n549) );
  NAND2_X1 U616 ( .A1(n550), .A2(n549), .ZN(n551) );
  NOR2_X1 U617 ( .A1(n552), .A2(n551), .ZN(n979) );
  INV_X1 U618 ( .A(n979), .ZN(G299) );
  NAND2_X1 U619 ( .A1(G85), .A2(n652), .ZN(n554) );
  NAND2_X1 U620 ( .A1(G72), .A2(n655), .ZN(n553) );
  NAND2_X1 U621 ( .A1(n554), .A2(n553), .ZN(n558) );
  NAND2_X1 U622 ( .A1(G60), .A2(n665), .ZN(n556) );
  NAND2_X1 U623 ( .A1(G47), .A2(n661), .ZN(n555) );
  NAND2_X1 U624 ( .A1(n556), .A2(n555), .ZN(n557) );
  OR2_X1 U625 ( .A1(n558), .A2(n557), .ZN(G290) );
  NAND2_X1 U626 ( .A1(G64), .A2(n665), .ZN(n560) );
  NAND2_X1 U627 ( .A1(G52), .A2(n661), .ZN(n559) );
  NAND2_X1 U628 ( .A1(n560), .A2(n559), .ZN(n565) );
  NAND2_X1 U629 ( .A1(G90), .A2(n652), .ZN(n562) );
  NAND2_X1 U630 ( .A1(G77), .A2(n655), .ZN(n561) );
  NAND2_X1 U631 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U632 ( .A(KEYINPUT9), .B(n563), .Z(n564) );
  NOR2_X1 U633 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U634 ( .A(KEYINPUT68), .B(n566), .ZN(G171) );
  INV_X1 U635 ( .A(G171), .ZN(G301) );
  XOR2_X1 U636 ( .A(G2446), .B(KEYINPUT106), .Z(n568) );
  XNOR2_X1 U637 ( .A(G2451), .B(G2430), .ZN(n567) );
  XNOR2_X1 U638 ( .A(n568), .B(n567), .ZN(n569) );
  XOR2_X1 U639 ( .A(n569), .B(G2427), .Z(n571) );
  XNOR2_X1 U640 ( .A(G1341), .B(G1348), .ZN(n570) );
  XNOR2_X1 U641 ( .A(n571), .B(n570), .ZN(n575) );
  XOR2_X1 U642 ( .A(G2443), .B(G2435), .Z(n573) );
  XNOR2_X1 U643 ( .A(G2438), .B(G2454), .ZN(n572) );
  XNOR2_X1 U644 ( .A(n573), .B(n572), .ZN(n574) );
  XOR2_X1 U645 ( .A(n575), .B(n574), .Z(n576) );
  AND2_X1 U646 ( .A1(G14), .A2(n576), .ZN(G401) );
  INV_X1 U647 ( .A(G57), .ZN(G237) );
  INV_X1 U648 ( .A(G132), .ZN(G219) );
  NAND2_X1 U649 ( .A1(G62), .A2(n665), .ZN(n578) );
  NAND2_X1 U650 ( .A1(G50), .A2(n661), .ZN(n577) );
  NAND2_X1 U651 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U652 ( .A(KEYINPUT82), .B(n579), .ZN(n582) );
  NAND2_X1 U653 ( .A1(G75), .A2(n655), .ZN(n580) );
  XNOR2_X1 U654 ( .A(KEYINPUT83), .B(n580), .ZN(n581) );
  NOR2_X1 U655 ( .A1(n582), .A2(n581), .ZN(n584) );
  NAND2_X1 U656 ( .A1(n652), .A2(G88), .ZN(n583) );
  NAND2_X1 U657 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U658 ( .A(KEYINPUT84), .B(n585), .ZN(G303) );
  INV_X1 U659 ( .A(G303), .ZN(G166) );
  NAND2_X1 U660 ( .A1(n884), .A2(G113), .ZN(n588) );
  NAND2_X1 U661 ( .A1(n629), .A2(G101), .ZN(n586) );
  XOR2_X1 U662 ( .A(KEYINPUT23), .B(n586), .Z(n587) );
  NAND2_X1 U663 ( .A1(n588), .A2(n587), .ZN(n593) );
  BUF_X1 U664 ( .A(n589), .Z(n880) );
  NAND2_X1 U665 ( .A1(G137), .A2(n880), .ZN(n591) );
  NAND2_X1 U666 ( .A1(G125), .A2(n885), .ZN(n590) );
  NAND2_X1 U667 ( .A1(n591), .A2(n590), .ZN(n592) );
  NOR2_X1 U668 ( .A1(n593), .A2(n592), .ZN(G160) );
  NAND2_X1 U669 ( .A1(G94), .A2(G452), .ZN(n594) );
  XNOR2_X1 U670 ( .A(n594), .B(KEYINPUT69), .ZN(G173) );
  XOR2_X1 U671 ( .A(KEYINPUT10), .B(KEYINPUT71), .Z(n596) );
  NAND2_X1 U672 ( .A1(G7), .A2(G661), .ZN(n595) );
  XNOR2_X1 U673 ( .A(n596), .B(n595), .ZN(G223) );
  INV_X1 U674 ( .A(G223), .ZN(n844) );
  NAND2_X1 U675 ( .A1(n844), .A2(G567), .ZN(n597) );
  XOR2_X1 U676 ( .A(KEYINPUT11), .B(n597), .Z(G234) );
  XOR2_X1 U677 ( .A(KEYINPUT72), .B(KEYINPUT14), .Z(n599) );
  NAND2_X1 U678 ( .A1(G56), .A2(n665), .ZN(n598) );
  XNOR2_X1 U679 ( .A(n599), .B(n598), .ZN(n605) );
  NAND2_X1 U680 ( .A1(n652), .A2(G81), .ZN(n600) );
  XNOR2_X1 U681 ( .A(n600), .B(KEYINPUT12), .ZN(n602) );
  NAND2_X1 U682 ( .A1(G68), .A2(n655), .ZN(n601) );
  NAND2_X1 U683 ( .A1(n602), .A2(n601), .ZN(n603) );
  XOR2_X1 U684 ( .A(KEYINPUT13), .B(n603), .Z(n604) );
  NOR2_X1 U685 ( .A1(n605), .A2(n604), .ZN(n607) );
  NAND2_X1 U686 ( .A1(n661), .A2(G43), .ZN(n606) );
  NAND2_X1 U687 ( .A1(n607), .A2(n606), .ZN(n980) );
  INV_X1 U688 ( .A(G860), .ZN(n643) );
  OR2_X1 U689 ( .A1(n980), .A2(n643), .ZN(G153) );
  NAND2_X1 U690 ( .A1(G79), .A2(n655), .ZN(n609) );
  NAND2_X1 U691 ( .A1(G54), .A2(n661), .ZN(n608) );
  NAND2_X1 U692 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U693 ( .A(KEYINPUT74), .B(n610), .ZN(n613) );
  NAND2_X1 U694 ( .A1(G92), .A2(n652), .ZN(n611) );
  XNOR2_X1 U695 ( .A(KEYINPUT73), .B(n611), .ZN(n612) );
  NOR2_X1 U696 ( .A1(n613), .A2(n612), .ZN(n615) );
  NAND2_X1 U697 ( .A1(n665), .A2(G66), .ZN(n614) );
  NAND2_X1 U698 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U699 ( .A(KEYINPUT15), .B(n616), .ZN(n995) );
  NOR2_X1 U700 ( .A1(n995), .A2(G868), .ZN(n617) );
  XNOR2_X1 U701 ( .A(n617), .B(KEYINPUT75), .ZN(n619) );
  NAND2_X1 U702 ( .A1(G868), .A2(G301), .ZN(n618) );
  NAND2_X1 U703 ( .A1(n619), .A2(n618), .ZN(G284) );
  NOR2_X1 U704 ( .A1(G868), .A2(G299), .ZN(n621) );
  INV_X1 U705 ( .A(G868), .ZN(n678) );
  NOR2_X1 U706 ( .A1(G286), .A2(n678), .ZN(n620) );
  NOR2_X1 U707 ( .A1(n621), .A2(n620), .ZN(G297) );
  NAND2_X1 U708 ( .A1(G559), .A2(n643), .ZN(n622) );
  XOR2_X1 U709 ( .A(KEYINPUT77), .B(n622), .Z(n623) );
  NAND2_X1 U710 ( .A1(n623), .A2(n995), .ZN(n624) );
  XNOR2_X1 U711 ( .A(n624), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U712 ( .A1(n995), .A2(G868), .ZN(n625) );
  NOR2_X1 U713 ( .A1(G559), .A2(n625), .ZN(n626) );
  XNOR2_X1 U714 ( .A(n626), .B(KEYINPUT78), .ZN(n628) );
  NOR2_X1 U715 ( .A1(n980), .A2(G868), .ZN(n627) );
  NOR2_X1 U716 ( .A1(n628), .A2(n627), .ZN(G282) );
  INV_X1 U717 ( .A(n629), .ZN(n630) );
  INV_X1 U718 ( .A(n630), .ZN(n881) );
  NAND2_X1 U719 ( .A1(G99), .A2(n881), .ZN(n631) );
  XOR2_X1 U720 ( .A(KEYINPUT79), .B(n631), .Z(n633) );
  NAND2_X1 U721 ( .A1(n884), .A2(G111), .ZN(n632) );
  NAND2_X1 U722 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U723 ( .A(KEYINPUT80), .B(n634), .ZN(n639) );
  NAND2_X1 U724 ( .A1(G123), .A2(n885), .ZN(n635) );
  XNOR2_X1 U725 ( .A(n635), .B(KEYINPUT18), .ZN(n637) );
  NAND2_X1 U726 ( .A1(n880), .A2(G135), .ZN(n636) );
  NAND2_X1 U727 ( .A1(n637), .A2(n636), .ZN(n638) );
  NOR2_X1 U728 ( .A1(n639), .A2(n638), .ZN(n949) );
  XNOR2_X1 U729 ( .A(n949), .B(G2096), .ZN(n641) );
  INV_X1 U730 ( .A(G2100), .ZN(n640) );
  NAND2_X1 U731 ( .A1(n641), .A2(n640), .ZN(G156) );
  NAND2_X1 U732 ( .A1(G559), .A2(n995), .ZN(n642) );
  XOR2_X1 U733 ( .A(n980), .B(n642), .Z(n676) );
  NAND2_X1 U734 ( .A1(n643), .A2(n676), .ZN(n651) );
  NAND2_X1 U735 ( .A1(G93), .A2(n652), .ZN(n645) );
  NAND2_X1 U736 ( .A1(G80), .A2(n655), .ZN(n644) );
  NAND2_X1 U737 ( .A1(n645), .A2(n644), .ZN(n648) );
  NAND2_X1 U738 ( .A1(G55), .A2(n661), .ZN(n646) );
  XNOR2_X1 U739 ( .A(KEYINPUT81), .B(n646), .ZN(n647) );
  NOR2_X1 U740 ( .A1(n648), .A2(n647), .ZN(n650) );
  NAND2_X1 U741 ( .A1(n665), .A2(G67), .ZN(n649) );
  NAND2_X1 U742 ( .A1(n650), .A2(n649), .ZN(n679) );
  XNOR2_X1 U743 ( .A(n651), .B(n679), .ZN(G145) );
  NAND2_X1 U744 ( .A1(G61), .A2(n665), .ZN(n654) );
  NAND2_X1 U745 ( .A1(G86), .A2(n652), .ZN(n653) );
  NAND2_X1 U746 ( .A1(n654), .A2(n653), .ZN(n658) );
  NAND2_X1 U747 ( .A1(n655), .A2(G73), .ZN(n656) );
  XOR2_X1 U748 ( .A(KEYINPUT2), .B(n656), .Z(n657) );
  NOR2_X1 U749 ( .A1(n658), .A2(n657), .ZN(n660) );
  NAND2_X1 U750 ( .A1(n661), .A2(G48), .ZN(n659) );
  NAND2_X1 U751 ( .A1(n660), .A2(n659), .ZN(G305) );
  NAND2_X1 U752 ( .A1(G49), .A2(n661), .ZN(n663) );
  NAND2_X1 U753 ( .A1(G74), .A2(G651), .ZN(n662) );
  NAND2_X1 U754 ( .A1(n663), .A2(n662), .ZN(n664) );
  NOR2_X1 U755 ( .A1(n665), .A2(n664), .ZN(n668) );
  NAND2_X1 U756 ( .A1(n666), .A2(G87), .ZN(n667) );
  NAND2_X1 U757 ( .A1(n668), .A2(n667), .ZN(G288) );
  XNOR2_X1 U758 ( .A(G303), .B(G305), .ZN(n671) );
  XNOR2_X1 U759 ( .A(G288), .B(KEYINPUT85), .ZN(n672) );
  XNOR2_X1 U760 ( .A(n673), .B(n672), .ZN(n675) );
  XOR2_X1 U761 ( .A(n898), .B(n676), .Z(n677) );
  NOR2_X1 U762 ( .A1(n678), .A2(n677), .ZN(n681) );
  NOR2_X1 U763 ( .A1(G868), .A2(n679), .ZN(n680) );
  NOR2_X1 U764 ( .A1(n681), .A2(n680), .ZN(G295) );
  NAND2_X1 U765 ( .A1(G2078), .A2(G2084), .ZN(n683) );
  XOR2_X1 U766 ( .A(KEYINPUT86), .B(KEYINPUT20), .Z(n682) );
  XNOR2_X1 U767 ( .A(n683), .B(n682), .ZN(n684) );
  NAND2_X1 U768 ( .A1(G2090), .A2(n684), .ZN(n685) );
  XNOR2_X1 U769 ( .A(KEYINPUT21), .B(n685), .ZN(n686) );
  NAND2_X1 U770 ( .A1(n686), .A2(G2072), .ZN(G158) );
  XOR2_X1 U771 ( .A(KEYINPUT70), .B(G82), .Z(G220) );
  XNOR2_X1 U772 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U773 ( .A1(G220), .A2(G219), .ZN(n688) );
  XNOR2_X1 U774 ( .A(KEYINPUT22), .B(KEYINPUT87), .ZN(n687) );
  XNOR2_X1 U775 ( .A(n688), .B(n687), .ZN(n689) );
  NOR2_X1 U776 ( .A1(n689), .A2(G218), .ZN(n690) );
  NAND2_X1 U777 ( .A1(G96), .A2(n690), .ZN(n850) );
  NAND2_X1 U778 ( .A1(n850), .A2(G2106), .ZN(n694) );
  NAND2_X1 U779 ( .A1(G69), .A2(G120), .ZN(n691) );
  NOR2_X1 U780 ( .A1(G237), .A2(n691), .ZN(n692) );
  NAND2_X1 U781 ( .A1(G108), .A2(n692), .ZN(n851) );
  NAND2_X1 U782 ( .A1(n851), .A2(G567), .ZN(n693) );
  NAND2_X1 U783 ( .A1(n694), .A2(n693), .ZN(n852) );
  NAND2_X1 U784 ( .A1(G483), .A2(G661), .ZN(n695) );
  NOR2_X1 U785 ( .A1(n852), .A2(n695), .ZN(n849) );
  NAND2_X1 U786 ( .A1(n849), .A2(G36), .ZN(G176) );
  NAND2_X1 U787 ( .A1(G160), .A2(G40), .ZN(n804) );
  NOR2_X1 U788 ( .A1(G164), .A2(G1384), .ZN(n805) );
  INV_X1 U789 ( .A(n805), .ZN(n696) );
  XNOR2_X1 U790 ( .A(KEYINPUT64), .B(n697), .ZN(n725) );
  INV_X1 U791 ( .A(n725), .ZN(n749) );
  NOR2_X1 U792 ( .A1(G1981), .A2(G305), .ZN(n698) );
  XOR2_X1 U793 ( .A(n698), .B(KEYINPUT24), .Z(n699) );
  NOR2_X1 U794 ( .A1(n786), .A2(n699), .ZN(n778) );
  XOR2_X1 U795 ( .A(G1996), .B(KEYINPUT94), .Z(n928) );
  INV_X1 U796 ( .A(n928), .ZN(n700) );
  AND2_X1 U797 ( .A1(n725), .A2(n700), .ZN(n702) );
  INV_X1 U798 ( .A(KEYINPUT26), .ZN(n701) );
  XNOR2_X1 U799 ( .A(n702), .B(n701), .ZN(n704) );
  NAND2_X1 U800 ( .A1(n749), .A2(G1341), .ZN(n703) );
  NAND2_X1 U801 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U802 ( .A1(n995), .A2(n711), .ZN(n710) );
  AND2_X1 U803 ( .A1(n749), .A2(G1348), .ZN(n706) );
  XNOR2_X1 U804 ( .A(n706), .B(KEYINPUT95), .ZN(n708) );
  NAND2_X1 U805 ( .A1(n725), .A2(G2067), .ZN(n707) );
  NAND2_X1 U806 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U807 ( .A1(n710), .A2(n709), .ZN(n713) );
  OR2_X1 U808 ( .A1(n995), .A2(n711), .ZN(n712) );
  NAND2_X1 U809 ( .A1(n713), .A2(n712), .ZN(n718) );
  NAND2_X1 U810 ( .A1(G2072), .A2(n725), .ZN(n714) );
  XNOR2_X1 U811 ( .A(n714), .B(KEYINPUT27), .ZN(n716) );
  INV_X1 U812 ( .A(G1956), .ZN(n1011) );
  NOR2_X1 U813 ( .A1(n725), .A2(n1011), .ZN(n715) );
  NOR2_X1 U814 ( .A1(n716), .A2(n715), .ZN(n719) );
  NAND2_X1 U815 ( .A1(n979), .A2(n719), .ZN(n717) );
  NAND2_X1 U816 ( .A1(n718), .A2(n717), .ZN(n722) );
  NOR2_X1 U817 ( .A1(n979), .A2(n719), .ZN(n720) );
  XOR2_X1 U818 ( .A(n720), .B(KEYINPUT28), .Z(n721) );
  NAND2_X1 U819 ( .A1(n722), .A2(n721), .ZN(n723) );
  XOR2_X1 U820 ( .A(KEYINPUT29), .B(n723), .Z(n730) );
  XOR2_X1 U821 ( .A(G2078), .B(KEYINPUT25), .Z(n724) );
  XNOR2_X1 U822 ( .A(KEYINPUT92), .B(n724), .ZN(n927) );
  NAND2_X1 U823 ( .A1(n725), .A2(n927), .ZN(n727) );
  NAND2_X1 U824 ( .A1(n749), .A2(G1961), .ZN(n726) );
  NAND2_X1 U825 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U826 ( .A(n728), .B(KEYINPUT93), .ZN(n731) );
  NAND2_X1 U827 ( .A1(n731), .A2(G171), .ZN(n729) );
  NAND2_X1 U828 ( .A1(n730), .A2(n729), .ZN(n740) );
  NOR2_X1 U829 ( .A1(n731), .A2(G171), .ZN(n736) );
  NOR2_X1 U830 ( .A1(n749), .A2(G2084), .ZN(n745) );
  NOR2_X1 U831 ( .A1(G1966), .A2(n786), .ZN(n741) );
  NOR2_X1 U832 ( .A1(n745), .A2(n741), .ZN(n732) );
  AND2_X1 U833 ( .A1(n732), .A2(G8), .ZN(n733) );
  XNOR2_X1 U834 ( .A(n733), .B(n521), .ZN(n734) );
  NOR2_X1 U835 ( .A1(G168), .A2(n734), .ZN(n735) );
  NOR2_X1 U836 ( .A1(n736), .A2(n735), .ZN(n738) );
  NAND2_X1 U837 ( .A1(n740), .A2(n739), .ZN(n753) );
  INV_X1 U838 ( .A(n753), .ZN(n742) );
  XNOR2_X1 U839 ( .A(n744), .B(n743), .ZN(n747) );
  NAND2_X1 U840 ( .A1(G8), .A2(n745), .ZN(n746) );
  NAND2_X1 U841 ( .A1(n747), .A2(n746), .ZN(n748) );
  XOR2_X1 U842 ( .A(KEYINPUT99), .B(KEYINPUT32), .Z(n758) );
  NOR2_X1 U843 ( .A1(n749), .A2(G2090), .ZN(n751) );
  NOR2_X1 U844 ( .A1(G1971), .A2(n786), .ZN(n750) );
  NOR2_X1 U845 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U846 ( .A1(G303), .A2(n752), .ZN(n755) );
  NAND2_X1 U847 ( .A1(G286), .A2(n753), .ZN(n754) );
  NAND2_X1 U848 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U849 ( .A1(G8), .A2(n756), .ZN(n757) );
  XNOR2_X1 U850 ( .A(n758), .B(n757), .ZN(n781) );
  NOR2_X1 U851 ( .A1(G1976), .A2(G288), .ZN(n987) );
  INV_X1 U852 ( .A(n786), .ZN(n761) );
  NAND2_X1 U853 ( .A1(n987), .A2(n761), .ZN(n759) );
  NAND2_X1 U854 ( .A1(n759), .A2(KEYINPUT33), .ZN(n768) );
  INV_X1 U855 ( .A(n768), .ZN(n764) );
  INV_X1 U856 ( .A(KEYINPUT33), .ZN(n760) );
  NAND2_X1 U857 ( .A1(G1976), .A2(G288), .ZN(n988) );
  AND2_X1 U858 ( .A1(n760), .A2(n988), .ZN(n762) );
  AND2_X1 U859 ( .A1(n762), .A2(n761), .ZN(n763) );
  OR2_X1 U860 ( .A1(n764), .A2(n763), .ZN(n766) );
  AND2_X1 U861 ( .A1(n781), .A2(n766), .ZN(n765) );
  NAND2_X1 U862 ( .A1(n782), .A2(n765), .ZN(n773) );
  INV_X1 U863 ( .A(n766), .ZN(n771) );
  NOR2_X1 U864 ( .A1(G303), .A2(G1971), .ZN(n767) );
  NOR2_X1 U865 ( .A1(n987), .A2(n767), .ZN(n769) );
  AND2_X1 U866 ( .A1(n769), .A2(n768), .ZN(n770) );
  OR2_X1 U867 ( .A1(n771), .A2(n770), .ZN(n772) );
  NAND2_X1 U868 ( .A1(n773), .A2(n772), .ZN(n774) );
  XNOR2_X1 U869 ( .A(G1981), .B(G305), .ZN(n1002) );
  NOR2_X1 U870 ( .A1(n778), .A2(n777), .ZN(n830) );
  NAND2_X1 U871 ( .A1(G8), .A2(G166), .ZN(n779) );
  NOR2_X1 U872 ( .A1(G2090), .A2(n779), .ZN(n780) );
  XNOR2_X1 U873 ( .A(n780), .B(KEYINPUT101), .ZN(n784) );
  NAND2_X1 U874 ( .A1(n782), .A2(n781), .ZN(n783) );
  NAND2_X1 U875 ( .A1(n784), .A2(n783), .ZN(n785) );
  XNOR2_X1 U876 ( .A(n785), .B(KEYINPUT102), .ZN(n787) );
  NAND2_X1 U877 ( .A1(n787), .A2(n786), .ZN(n828) );
  NAND2_X1 U878 ( .A1(n881), .A2(G105), .ZN(n788) );
  XOR2_X1 U879 ( .A(KEYINPUT38), .B(n788), .Z(n793) );
  NAND2_X1 U880 ( .A1(G117), .A2(n884), .ZN(n790) );
  NAND2_X1 U881 ( .A1(G129), .A2(n885), .ZN(n789) );
  NAND2_X1 U882 ( .A1(n790), .A2(n789), .ZN(n791) );
  XOR2_X1 U883 ( .A(KEYINPUT91), .B(n791), .Z(n792) );
  NOR2_X1 U884 ( .A1(n793), .A2(n792), .ZN(n795) );
  NAND2_X1 U885 ( .A1(n880), .A2(G141), .ZN(n794) );
  NAND2_X1 U886 ( .A1(n795), .A2(n794), .ZN(n891) );
  NOR2_X1 U887 ( .A1(G1996), .A2(n891), .ZN(n964) );
  NAND2_X1 U888 ( .A1(n880), .A2(G131), .ZN(n797) );
  NAND2_X1 U889 ( .A1(G95), .A2(n881), .ZN(n796) );
  NAND2_X1 U890 ( .A1(n797), .A2(n796), .ZN(n801) );
  NAND2_X1 U891 ( .A1(G107), .A2(n884), .ZN(n799) );
  NAND2_X1 U892 ( .A1(G119), .A2(n885), .ZN(n798) );
  NAND2_X1 U893 ( .A1(n799), .A2(n798), .ZN(n800) );
  NOR2_X1 U894 ( .A1(n801), .A2(n800), .ZN(n876) );
  INV_X1 U895 ( .A(G1991), .ZN(n932) );
  NOR2_X1 U896 ( .A1(n876), .A2(n932), .ZN(n803) );
  AND2_X1 U897 ( .A1(n891), .A2(G1996), .ZN(n802) );
  NOR2_X1 U898 ( .A1(n803), .A2(n802), .ZN(n958) );
  NOR2_X1 U899 ( .A1(n805), .A2(n804), .ZN(n836) );
  INV_X1 U900 ( .A(n836), .ZN(n806) );
  NOR2_X1 U901 ( .A1(n958), .A2(n806), .ZN(n832) );
  NOR2_X1 U902 ( .A1(G1986), .A2(G290), .ZN(n808) );
  AND2_X1 U903 ( .A1(n932), .A2(n876), .ZN(n807) );
  XOR2_X1 U904 ( .A(KEYINPUT103), .B(n807), .Z(n960) );
  NOR2_X1 U905 ( .A1(n808), .A2(n960), .ZN(n809) );
  NOR2_X1 U906 ( .A1(n832), .A2(n809), .ZN(n810) );
  XNOR2_X1 U907 ( .A(n810), .B(KEYINPUT104), .ZN(n811) );
  NOR2_X1 U908 ( .A1(n964), .A2(n811), .ZN(n812) );
  XNOR2_X1 U909 ( .A(n812), .B(KEYINPUT39), .ZN(n823) );
  NAND2_X1 U910 ( .A1(n880), .A2(G140), .ZN(n814) );
  NAND2_X1 U911 ( .A1(G104), .A2(n881), .ZN(n813) );
  NAND2_X1 U912 ( .A1(n814), .A2(n813), .ZN(n815) );
  XNOR2_X1 U913 ( .A(KEYINPUT34), .B(n815), .ZN(n820) );
  NAND2_X1 U914 ( .A1(G116), .A2(n884), .ZN(n817) );
  NAND2_X1 U915 ( .A1(G128), .A2(n885), .ZN(n816) );
  NAND2_X1 U916 ( .A1(n817), .A2(n816), .ZN(n818) );
  XOR2_X1 U917 ( .A(KEYINPUT35), .B(n818), .Z(n819) );
  NOR2_X1 U918 ( .A1(n820), .A2(n819), .ZN(n821) );
  XOR2_X1 U919 ( .A(KEYINPUT36), .B(n821), .Z(n877) );
  XOR2_X1 U920 ( .A(G2067), .B(KEYINPUT37), .Z(n824) );
  AND2_X1 U921 ( .A1(n877), .A2(n824), .ZN(n950) );
  NAND2_X1 U922 ( .A1(n950), .A2(n836), .ZN(n822) );
  XNOR2_X1 U923 ( .A(n822), .B(KEYINPUT90), .ZN(n833) );
  NAND2_X1 U924 ( .A1(n823), .A2(n833), .ZN(n826) );
  NOR2_X1 U925 ( .A1(n824), .A2(n877), .ZN(n825) );
  XNOR2_X1 U926 ( .A(n825), .B(KEYINPUT105), .ZN(n967) );
  NAND2_X1 U927 ( .A1(n826), .A2(n967), .ZN(n827) );
  NAND2_X1 U928 ( .A1(n827), .A2(n836), .ZN(n831) );
  AND2_X1 U929 ( .A1(n828), .A2(n831), .ZN(n829) );
  NAND2_X1 U930 ( .A1(n830), .A2(n829), .ZN(n842) );
  INV_X1 U931 ( .A(n831), .ZN(n840) );
  INV_X1 U932 ( .A(n832), .ZN(n834) );
  NAND2_X1 U933 ( .A1(n834), .A2(n833), .ZN(n838) );
  XOR2_X1 U934 ( .A(G1986), .B(KEYINPUT89), .Z(n835) );
  XNOR2_X1 U935 ( .A(G290), .B(n835), .ZN(n982) );
  AND2_X1 U936 ( .A1(n982), .A2(n836), .ZN(n837) );
  NOR2_X1 U937 ( .A1(n838), .A2(n837), .ZN(n839) );
  OR2_X1 U938 ( .A1(n840), .A2(n839), .ZN(n841) );
  XNOR2_X1 U939 ( .A(n843), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U940 ( .A1(G2106), .A2(n844), .ZN(G217) );
  NAND2_X1 U941 ( .A1(G15), .A2(G2), .ZN(n845) );
  XNOR2_X1 U942 ( .A(KEYINPUT107), .B(n845), .ZN(n846) );
  NAND2_X1 U943 ( .A1(n846), .A2(G661), .ZN(n847) );
  XNOR2_X1 U944 ( .A(KEYINPUT108), .B(n847), .ZN(G259) );
  NAND2_X1 U945 ( .A1(G3), .A2(G1), .ZN(n848) );
  NAND2_X1 U946 ( .A1(n849), .A2(n848), .ZN(G188) );
  NOR2_X1 U947 ( .A1(n851), .A2(n850), .ZN(G325) );
  XNOR2_X1 U948 ( .A(KEYINPUT109), .B(G325), .ZN(G261) );
  INV_X1 U950 ( .A(G120), .ZN(G236) );
  INV_X1 U951 ( .A(G96), .ZN(G221) );
  INV_X1 U952 ( .A(G69), .ZN(G235) );
  INV_X1 U953 ( .A(n852), .ZN(G319) );
  XOR2_X1 U954 ( .A(KEYINPUT110), .B(KEYINPUT44), .Z(n854) );
  NAND2_X1 U955 ( .A1(G124), .A2(n885), .ZN(n853) );
  XNOR2_X1 U956 ( .A(n854), .B(n853), .ZN(n857) );
  NAND2_X1 U957 ( .A1(n880), .A2(G136), .ZN(n855) );
  XNOR2_X1 U958 ( .A(KEYINPUT111), .B(n855), .ZN(n856) );
  NOR2_X1 U959 ( .A1(n857), .A2(n856), .ZN(n858) );
  XNOR2_X1 U960 ( .A(n858), .B(KEYINPUT112), .ZN(n860) );
  NAND2_X1 U961 ( .A1(G112), .A2(n884), .ZN(n859) );
  NAND2_X1 U962 ( .A1(n860), .A2(n859), .ZN(n863) );
  NAND2_X1 U963 ( .A1(G100), .A2(n881), .ZN(n861) );
  XNOR2_X1 U964 ( .A(KEYINPUT113), .B(n861), .ZN(n862) );
  NOR2_X1 U965 ( .A1(n863), .A2(n862), .ZN(G162) );
  XOR2_X1 U966 ( .A(KEYINPUT48), .B(KEYINPUT115), .Z(n874) );
  NAND2_X1 U967 ( .A1(G118), .A2(n884), .ZN(n865) );
  NAND2_X1 U968 ( .A1(G130), .A2(n885), .ZN(n864) );
  NAND2_X1 U969 ( .A1(n865), .A2(n864), .ZN(n871) );
  NAND2_X1 U970 ( .A1(n880), .A2(G142), .ZN(n867) );
  NAND2_X1 U971 ( .A1(G106), .A2(n881), .ZN(n866) );
  NAND2_X1 U972 ( .A1(n867), .A2(n866), .ZN(n868) );
  XOR2_X1 U973 ( .A(KEYINPUT45), .B(n868), .Z(n869) );
  XNOR2_X1 U974 ( .A(KEYINPUT114), .B(n869), .ZN(n870) );
  NOR2_X1 U975 ( .A1(n871), .A2(n870), .ZN(n872) );
  XNOR2_X1 U976 ( .A(n872), .B(KEYINPUT46), .ZN(n873) );
  XNOR2_X1 U977 ( .A(n874), .B(n873), .ZN(n875) );
  XOR2_X1 U978 ( .A(n875), .B(n949), .Z(n879) );
  XNOR2_X1 U979 ( .A(n877), .B(n876), .ZN(n878) );
  XNOR2_X1 U980 ( .A(n879), .B(n878), .ZN(n896) );
  NAND2_X1 U981 ( .A1(n880), .A2(G139), .ZN(n883) );
  NAND2_X1 U982 ( .A1(G103), .A2(n881), .ZN(n882) );
  NAND2_X1 U983 ( .A1(n883), .A2(n882), .ZN(n890) );
  NAND2_X1 U984 ( .A1(G115), .A2(n884), .ZN(n887) );
  NAND2_X1 U985 ( .A1(G127), .A2(n885), .ZN(n886) );
  NAND2_X1 U986 ( .A1(n887), .A2(n886), .ZN(n888) );
  XOR2_X1 U987 ( .A(KEYINPUT47), .B(n888), .Z(n889) );
  NOR2_X1 U988 ( .A1(n890), .A2(n889), .ZN(n951) );
  XNOR2_X1 U989 ( .A(n951), .B(n891), .ZN(n893) );
  XNOR2_X1 U990 ( .A(G164), .B(G160), .ZN(n892) );
  XNOR2_X1 U991 ( .A(n893), .B(n892), .ZN(n894) );
  XOR2_X1 U992 ( .A(G162), .B(n894), .Z(n895) );
  XNOR2_X1 U993 ( .A(n896), .B(n895), .ZN(n897) );
  NOR2_X1 U994 ( .A1(G37), .A2(n897), .ZN(G395) );
  XNOR2_X1 U995 ( .A(n980), .B(n898), .ZN(n901) );
  XNOR2_X1 U996 ( .A(G301), .B(n995), .ZN(n899) );
  NOR2_X1 U997 ( .A1(G37), .A2(n902), .ZN(G397) );
  XOR2_X1 U998 ( .A(G2100), .B(G2096), .Z(n904) );
  XNOR2_X1 U999 ( .A(KEYINPUT42), .B(G2678), .ZN(n903) );
  XNOR2_X1 U1000 ( .A(n904), .B(n903), .ZN(n908) );
  XOR2_X1 U1001 ( .A(KEYINPUT43), .B(G2072), .Z(n906) );
  XNOR2_X1 U1002 ( .A(G2067), .B(G2090), .ZN(n905) );
  XNOR2_X1 U1003 ( .A(n906), .B(n905), .ZN(n907) );
  XOR2_X1 U1004 ( .A(n908), .B(n907), .Z(n910) );
  XNOR2_X1 U1005 ( .A(G2078), .B(G2084), .ZN(n909) );
  XNOR2_X1 U1006 ( .A(n910), .B(n909), .ZN(G227) );
  XOR2_X1 U1007 ( .A(G1976), .B(G1956), .Z(n912) );
  XNOR2_X1 U1008 ( .A(G1986), .B(G1971), .ZN(n911) );
  XNOR2_X1 U1009 ( .A(n912), .B(n911), .ZN(n913) );
  XOR2_X1 U1010 ( .A(n913), .B(G2474), .Z(n915) );
  XNOR2_X1 U1011 ( .A(G1966), .B(G1981), .ZN(n914) );
  XNOR2_X1 U1012 ( .A(n915), .B(n914), .ZN(n919) );
  XOR2_X1 U1013 ( .A(KEYINPUT41), .B(G1961), .Z(n917) );
  XNOR2_X1 U1014 ( .A(G1996), .B(G1991), .ZN(n916) );
  XNOR2_X1 U1015 ( .A(n917), .B(n916), .ZN(n918) );
  XNOR2_X1 U1016 ( .A(n919), .B(n918), .ZN(G229) );
  NOR2_X1 U1017 ( .A1(G395), .A2(G397), .ZN(n920) );
  XOR2_X1 U1018 ( .A(KEYINPUT116), .B(n920), .Z(n921) );
  NOR2_X1 U1019 ( .A1(G401), .A2(n921), .ZN(n922) );
  NAND2_X1 U1020 ( .A1(G319), .A2(n922), .ZN(n925) );
  NOR2_X1 U1021 ( .A1(G227), .A2(G229), .ZN(n923) );
  XNOR2_X1 U1022 ( .A(KEYINPUT49), .B(n923), .ZN(n924) );
  NOR2_X1 U1023 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1024 ( .A(KEYINPUT117), .B(n926), .ZN(G225) );
  INV_X1 U1025 ( .A(G225), .ZN(G308) );
  INV_X1 U1026 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1027 ( .A(G2090), .B(G35), .ZN(n942) );
  XOR2_X1 U1028 ( .A(n927), .B(G27), .Z(n930) );
  XNOR2_X1 U1029 ( .A(n928), .B(G32), .ZN(n929) );
  NAND2_X1 U1030 ( .A1(n930), .A2(n929), .ZN(n939) );
  XNOR2_X1 U1031 ( .A(KEYINPUT119), .B(G2067), .ZN(n931) );
  XNOR2_X1 U1032 ( .A(n931), .B(G26), .ZN(n937) );
  XNOR2_X1 U1033 ( .A(G25), .B(n932), .ZN(n933) );
  NAND2_X1 U1034 ( .A1(n933), .A2(G28), .ZN(n935) );
  XNOR2_X1 U1035 ( .A(G33), .B(G2072), .ZN(n934) );
  NOR2_X1 U1036 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1037 ( .A1(n937), .A2(n936), .ZN(n938) );
  NOR2_X1 U1038 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1039 ( .A(KEYINPUT53), .B(n940), .ZN(n941) );
  NOR2_X1 U1040 ( .A1(n942), .A2(n941), .ZN(n945) );
  XOR2_X1 U1041 ( .A(G2084), .B(G34), .Z(n943) );
  XNOR2_X1 U1042 ( .A(KEYINPUT54), .B(n943), .ZN(n944) );
  NAND2_X1 U1043 ( .A1(n945), .A2(n944), .ZN(n948) );
  NOR2_X1 U1044 ( .A1(G29), .A2(KEYINPUT55), .ZN(n946) );
  NAND2_X1 U1045 ( .A1(n948), .A2(n946), .ZN(n947) );
  NAND2_X1 U1046 ( .A1(G11), .A2(n947), .ZN(n978) );
  INV_X1 U1047 ( .A(KEYINPUT55), .ZN(n972) );
  OR2_X1 U1048 ( .A1(n972), .A2(n948), .ZN(n976) );
  NOR2_X1 U1049 ( .A1(n950), .A2(n949), .ZN(n962) );
  XOR2_X1 U1050 ( .A(G2072), .B(n951), .Z(n953) );
  XOR2_X1 U1051 ( .A(G164), .B(G2078), .Z(n952) );
  NOR2_X1 U1052 ( .A1(n953), .A2(n952), .ZN(n954) );
  XOR2_X1 U1053 ( .A(KEYINPUT50), .B(n954), .Z(n956) );
  XOR2_X1 U1054 ( .A(G160), .B(G2084), .Z(n955) );
  NOR2_X1 U1055 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1056 ( .A1(n958), .A2(n957), .ZN(n959) );
  NOR2_X1 U1057 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1058 ( .A1(n962), .A2(n961), .ZN(n970) );
  XOR2_X1 U1059 ( .A(G2090), .B(G162), .Z(n963) );
  NOR2_X1 U1060 ( .A1(n964), .A2(n963), .ZN(n965) );
  XOR2_X1 U1061 ( .A(KEYINPUT118), .B(n965), .Z(n966) );
  XNOR2_X1 U1062 ( .A(n966), .B(KEYINPUT51), .ZN(n968) );
  NAND2_X1 U1063 ( .A1(n968), .A2(n967), .ZN(n969) );
  NOR2_X1 U1064 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1065 ( .A(n971), .B(KEYINPUT52), .ZN(n973) );
  NAND2_X1 U1066 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1067 ( .A1(G29), .A2(n974), .ZN(n975) );
  NAND2_X1 U1068 ( .A1(n976), .A2(n975), .ZN(n977) );
  NOR2_X1 U1069 ( .A1(n978), .A2(n977), .ZN(n1037) );
  XNOR2_X1 U1070 ( .A(G16), .B(KEYINPUT56), .ZN(n1007) );
  XNOR2_X1 U1071 ( .A(n979), .B(G1956), .ZN(n984) );
  XNOR2_X1 U1072 ( .A(G1341), .B(n980), .ZN(n981) );
  NOR2_X1 U1073 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1074 ( .A1(n984), .A2(n983), .ZN(n986) );
  XNOR2_X1 U1075 ( .A(G1961), .B(G301), .ZN(n985) );
  NOR2_X1 U1076 ( .A1(n986), .A2(n985), .ZN(n999) );
  INV_X1 U1077 ( .A(n987), .ZN(n989) );
  NAND2_X1 U1078 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1079 ( .A(KEYINPUT120), .B(n990), .ZN(n993) );
  XOR2_X1 U1080 ( .A(G1971), .B(G303), .Z(n991) );
  XNOR2_X1 U1081 ( .A(KEYINPUT121), .B(n991), .ZN(n992) );
  NOR2_X1 U1082 ( .A1(n993), .A2(n992), .ZN(n994) );
  XOR2_X1 U1083 ( .A(KEYINPUT122), .B(n994), .Z(n997) );
  XOR2_X1 U1084 ( .A(n995), .B(G1348), .Z(n996) );
  NOR2_X1 U1085 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1086 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1087 ( .A(KEYINPUT123), .B(n1000), .ZN(n1005) );
  XOR2_X1 U1088 ( .A(G168), .B(G1966), .Z(n1001) );
  NOR2_X1 U1089 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XOR2_X1 U1090 ( .A(KEYINPUT57), .B(n1003), .Z(n1004) );
  NAND2_X1 U1091 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1092 ( .A1(n1007), .A2(n1006), .ZN(n1034) );
  INV_X1 U1093 ( .A(G16), .ZN(n1032) );
  XNOR2_X1 U1094 ( .A(G1961), .B(G5), .ZN(n1009) );
  XNOR2_X1 U1095 ( .A(G1966), .B(G21), .ZN(n1008) );
  NOR2_X1 U1096 ( .A1(n1009), .A2(n1008), .ZN(n1022) );
  XNOR2_X1 U1097 ( .A(KEYINPUT60), .B(KEYINPUT125), .ZN(n1020) );
  XNOR2_X1 U1098 ( .A(KEYINPUT59), .B(G1348), .ZN(n1010) );
  XNOR2_X1 U1099 ( .A(n1010), .B(G4), .ZN(n1018) );
  XNOR2_X1 U1100 ( .A(G20), .B(n1011), .ZN(n1015) );
  XNOR2_X1 U1101 ( .A(G1341), .B(G19), .ZN(n1013) );
  XNOR2_X1 U1102 ( .A(G1981), .B(G6), .ZN(n1012) );
  NOR2_X1 U1103 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XOR2_X1 U1105 ( .A(KEYINPUT124), .B(n1016), .Z(n1017) );
  NAND2_X1 U1106 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1107 ( .A(n1020), .B(n1019), .ZN(n1021) );
  NAND2_X1 U1108 ( .A1(n1022), .A2(n1021), .ZN(n1029) );
  XNOR2_X1 U1109 ( .A(G1971), .B(G22), .ZN(n1024) );
  XNOR2_X1 U1110 ( .A(G23), .B(G1976), .ZN(n1023) );
  NOR2_X1 U1111 ( .A1(n1024), .A2(n1023), .ZN(n1026) );
  XOR2_X1 U1112 ( .A(G1986), .B(G24), .Z(n1025) );
  NAND2_X1 U1113 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1114 ( .A(KEYINPUT58), .B(n1027), .ZN(n1028) );
  NOR2_X1 U1115 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XNOR2_X1 U1116 ( .A(KEYINPUT61), .B(n1030), .ZN(n1031) );
  NAND2_X1 U1117 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NAND2_X1 U1118 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  XOR2_X1 U1119 ( .A(KEYINPUT126), .B(n1035), .Z(n1036) );
  NAND2_X1 U1120 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  XNOR2_X1 U1121 ( .A(n1038), .B(KEYINPUT127), .ZN(n1039) );
  XNOR2_X1 U1122 ( .A(KEYINPUT62), .B(n1039), .ZN(G311) );
  INV_X1 U1123 ( .A(G311), .ZN(G150) );
endmodule

