//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 1 1 0 1 1 0 0 1 0 1 1 0 1 1 0 1 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 1 0 1 0 0 0 1 1 0 0 0 1 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:21 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n738, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n763, new_n764,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n995, new_n996, new_n997, new_n998, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032;
  NOR2_X1   g000(.A1(G237), .A2(G953), .ZN(new_n187));
  NAND3_X1  g001(.A1(new_n187), .A2(G143), .A3(G214), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  AOI21_X1  g003(.A(G143), .B1(new_n187), .B2(G214), .ZN(new_n190));
  OAI21_X1  g004(.A(G131), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT17), .ZN(new_n192));
  INV_X1    g006(.A(G237), .ZN(new_n193));
  INV_X1    g007(.A(G953), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n193), .A2(new_n194), .A3(G214), .ZN(new_n195));
  INV_X1    g009(.A(G143), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G131), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n197), .A2(new_n198), .A3(new_n188), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n191), .A2(new_n192), .A3(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G146), .ZN(new_n201));
  INV_X1    g015(.A(G140), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G125), .ZN(new_n203));
  INV_X1    g017(.A(G125), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G140), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT16), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR3_X1   g022(.A1(new_n204), .A2(KEYINPUT16), .A3(G140), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n201), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(new_n209), .ZN(new_n211));
  OAI211_X1 g025(.A(new_n211), .B(G146), .C1(new_n206), .C2(new_n207), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n197), .A2(new_n188), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n213), .A2(KEYINPUT17), .A3(G131), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n200), .A2(new_n210), .A3(new_n212), .A4(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT76), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n204), .A2(G140), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n202), .A2(G125), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n203), .A2(new_n205), .A3(KEYINPUT76), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n219), .A2(new_n201), .A3(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(KEYINPUT77), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT77), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n219), .A2(new_n223), .A3(new_n201), .A4(new_n220), .ZN(new_n224));
  AOI22_X1  g038(.A1(new_n222), .A2(new_n224), .B1(G146), .B2(new_n206), .ZN(new_n225));
  AND2_X1   g039(.A1(KEYINPUT18), .A2(G131), .ZN(new_n226));
  XNOR2_X1  g040(.A(new_n213), .B(new_n226), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n215), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  XNOR2_X1  g042(.A(G113), .B(G122), .ZN(new_n229));
  OR2_X1    g043(.A1(new_n229), .A2(G104), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(G104), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n228), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT89), .ZN(new_n234));
  XNOR2_X1  g048(.A(new_n232), .B(new_n234), .ZN(new_n235));
  OAI211_X1 g049(.A(new_n235), .B(new_n215), .C1(new_n225), .C2(new_n227), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n233), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G902), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G475), .ZN(new_n240));
  INV_X1    g054(.A(G122), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G116), .ZN(new_n242));
  INV_X1    g056(.A(G116), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G122), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G107), .ZN(new_n246));
  INV_X1    g060(.A(G107), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n242), .A2(new_n244), .A3(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT13), .ZN(new_n250));
  INV_X1    g064(.A(G128), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n250), .B1(new_n251), .B2(G143), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(G143), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n196), .A2(G128), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n255), .A2(new_n250), .ZN(new_n256));
  OAI21_X1  g070(.A(G134), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(G134), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n255), .A2(new_n253), .A3(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n249), .A2(new_n257), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n255), .A2(new_n253), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G134), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(new_n259), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n243), .A2(KEYINPUT14), .A3(G122), .ZN(new_n264));
  OAI211_X1 g078(.A(G107), .B(new_n264), .C1(new_n245), .C2(KEYINPUT14), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n263), .A2(new_n248), .A3(new_n265), .ZN(new_n266));
  XNOR2_X1  g080(.A(KEYINPUT9), .B(G234), .ZN(new_n267));
  INV_X1    g081(.A(G217), .ZN(new_n268));
  NOR3_X1   g082(.A1(new_n267), .A2(new_n268), .A3(G953), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n260), .A2(new_n266), .A3(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n270), .B1(new_n260), .B2(new_n266), .ZN(new_n273));
  NOR3_X1   g087(.A1(new_n272), .A2(new_n273), .A3(G902), .ZN(new_n274));
  INV_X1    g088(.A(G478), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n275), .A2(KEYINPUT15), .ZN(new_n276));
  XNOR2_X1  g090(.A(new_n274), .B(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT20), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n191), .A2(new_n199), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT19), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n219), .A2(new_n280), .A3(new_n220), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n206), .A2(KEYINPUT19), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  OAI211_X1 g097(.A(new_n212), .B(new_n279), .C1(new_n283), .C2(G146), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n284), .B1(new_n225), .B2(new_n227), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(new_n232), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(new_n236), .ZN(new_n287));
  NOR2_X1   g101(.A1(G475), .A2(G902), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n278), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n288), .ZN(new_n290));
  AOI211_X1 g104(.A(KEYINPUT20), .B(new_n290), .C1(new_n286), .C2(new_n236), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n240), .B(new_n277), .C1(new_n289), .C2(new_n291), .ZN(new_n292));
  AND2_X1   g106(.A1(new_n194), .A2(G952), .ZN(new_n293));
  INV_X1    g107(.A(G234), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n293), .B1(new_n294), .B2(new_n193), .ZN(new_n295));
  AOI211_X1 g109(.A(new_n238), .B(new_n194), .C1(G234), .C2(G237), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  XNOR2_X1  g111(.A(KEYINPUT21), .B(G898), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n295), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(KEYINPUT90), .B1(new_n292), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n206), .A2(G146), .ZN(new_n303));
  AND2_X1   g117(.A1(new_n221), .A2(KEYINPUT77), .ZN(new_n304));
  INV_X1    g118(.A(new_n224), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n303), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(new_n227), .ZN(new_n307));
  AND3_X1   g121(.A1(new_n210), .A2(new_n212), .A3(new_n214), .ZN(new_n308));
  AOI22_X1  g122(.A1(new_n306), .A2(new_n307), .B1(new_n200), .B2(new_n308), .ZN(new_n309));
  AOI22_X1  g123(.A1(new_n309), .A2(new_n235), .B1(new_n285), .B2(new_n232), .ZN(new_n310));
  OAI21_X1  g124(.A(KEYINPUT20), .B1(new_n310), .B2(new_n290), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n287), .A2(new_n278), .A3(new_n288), .ZN(new_n312));
  AOI22_X1  g126(.A1(new_n311), .A2(new_n312), .B1(G475), .B2(new_n239), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT90), .ZN(new_n314));
  NAND4_X1  g128(.A1(new_n313), .A2(new_n314), .A3(new_n300), .A4(new_n277), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n302), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g130(.A(G214), .B1(G237), .B2(G902), .ZN(new_n317));
  XOR2_X1   g131(.A(new_n317), .B(KEYINPUT83), .Z(new_n318));
  INV_X1    g132(.A(G104), .ZN(new_n319));
  OAI21_X1  g133(.A(KEYINPUT3), .B1(new_n319), .B2(G107), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT3), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n321), .A2(new_n247), .A3(G104), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n247), .A2(G104), .ZN(new_n324));
  OAI21_X1  g138(.A(G101), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(KEYINPUT80), .A2(G101), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  NOR2_X1   g141(.A1(KEYINPUT80), .A2(G101), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n319), .A2(G107), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n329), .A2(new_n320), .A3(new_n322), .A4(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n325), .A2(new_n331), .A3(KEYINPUT4), .ZN(new_n332));
  INV_X1    g146(.A(G113), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(KEYINPUT2), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT2), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(G113), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(KEYINPUT67), .B1(new_n243), .B2(G119), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT67), .ZN(new_n340));
  INV_X1    g154(.A(G119), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n340), .A2(new_n341), .A3(G116), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n243), .A2(G119), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n339), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n338), .A2(new_n344), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n337), .A2(new_n339), .A3(new_n342), .A4(new_n343), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT4), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n348), .B(G101), .C1(new_n323), .C2(new_n324), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n332), .A2(new_n347), .A3(new_n349), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n319), .A2(G107), .ZN(new_n351));
  OAI21_X1  g165(.A(G101), .B1(new_n351), .B2(new_n324), .ZN(new_n352));
  OR2_X1    g166(.A1(KEYINPUT80), .A2(G101), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n353), .A2(new_n330), .A3(new_n326), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n352), .B1(new_n323), .B2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n243), .A2(G119), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT5), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n333), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n359), .B1(new_n344), .B2(new_n358), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n356), .A2(new_n346), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n350), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(KEYINPUT84), .ZN(new_n363));
  XNOR2_X1  g177(.A(G110), .B(G122), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT84), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n350), .A2(new_n361), .A3(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n363), .A2(new_n365), .A3(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT6), .ZN(new_n369));
  INV_X1    g183(.A(new_n362), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n369), .B1(new_n370), .B2(new_n364), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n368), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n201), .A2(G143), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT65), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n374), .B1(new_n196), .B2(G146), .ZN(new_n375));
  NOR3_X1   g189(.A1(new_n201), .A2(KEYINPUT65), .A3(G143), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n373), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(KEYINPUT0), .A2(G128), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n196), .A2(G146), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT64), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n380), .B1(new_n201), .B2(G143), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n196), .A2(KEYINPUT64), .A3(G146), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n379), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n378), .ZN(new_n384));
  NOR2_X1   g198(.A1(KEYINPUT0), .A2(G128), .ZN(new_n385));
  OR2_X1    g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  OAI22_X1  g200(.A1(new_n377), .A2(new_n378), .B1(new_n383), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(G125), .ZN(new_n388));
  OAI21_X1  g202(.A(KEYINPUT1), .B1(new_n196), .B2(G146), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(KEYINPUT66), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT66), .ZN(new_n391));
  OAI211_X1 g205(.A(new_n391), .B(KEYINPUT1), .C1(new_n196), .C2(G146), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n390), .A2(G128), .A3(new_n392), .ZN(new_n393));
  AND3_X1   g207(.A1(new_n196), .A2(KEYINPUT64), .A3(G146), .ZN(new_n394));
  AOI21_X1  g208(.A(KEYINPUT64), .B1(new_n196), .B2(G146), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n373), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n393), .A2(new_n396), .ZN(new_n397));
  OAI21_X1  g211(.A(KEYINPUT65), .B1(new_n201), .B2(G143), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n374), .A2(new_n196), .A3(G146), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n379), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n251), .A2(KEYINPUT1), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n397), .A2(new_n204), .A3(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT86), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n388), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n404), .B1(new_n388), .B2(new_n403), .ZN(new_n407));
  INV_X1    g221(.A(G224), .ZN(new_n408));
  OAI22_X1  g222(.A1(new_n406), .A2(new_n407), .B1(new_n408), .B2(G953), .ZN(new_n409));
  INV_X1    g223(.A(new_n407), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n408), .A2(G953), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n410), .A2(new_n411), .A3(new_n405), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n409), .A2(new_n412), .ZN(new_n413));
  XOR2_X1   g227(.A(KEYINPUT85), .B(KEYINPUT6), .Z(new_n414));
  NAND4_X1  g228(.A1(new_n363), .A2(new_n365), .A3(new_n367), .A4(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n372), .A2(new_n413), .A3(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT7), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n411), .A2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT87), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n397), .A2(new_n419), .A3(new_n204), .A4(new_n402), .ZN(new_n420));
  AND2_X1   g234(.A1(new_n420), .A2(new_n388), .ZN(new_n421));
  AOI22_X1  g235(.A1(new_n393), .A2(new_n396), .B1(new_n400), .B2(new_n401), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n419), .B1(new_n422), .B2(new_n204), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n418), .B1(new_n421), .B2(new_n424), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n364), .B(KEYINPUT8), .ZN(new_n426));
  AND4_X1   g240(.A1(new_n346), .A2(new_n360), .A3(new_n331), .A4(new_n352), .ZN(new_n427));
  AOI22_X1  g241(.A1(new_n360), .A2(new_n346), .B1(new_n331), .B2(new_n352), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n426), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n388), .A2(new_n403), .A3(new_n418), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(KEYINPUT88), .B1(new_n425), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n420), .A2(new_n388), .ZN(new_n433));
  OAI22_X1  g247(.A1(new_n433), .A2(new_n423), .B1(new_n417), .B2(new_n411), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT88), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n434), .A2(new_n435), .A3(new_n430), .A4(new_n429), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n370), .A2(new_n364), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n432), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n416), .A2(new_n438), .A3(new_n238), .ZN(new_n439));
  OAI21_X1  g253(.A(G210), .B1(G237), .B2(G902), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n416), .A2(new_n438), .A3(new_n238), .A4(new_n440), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n318), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(G469), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT1), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n446), .B1(G143), .B2(new_n201), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT81), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n251), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n389), .A2(KEYINPUT81), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n400), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n402), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n356), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT10), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT11), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n456), .B1(new_n258), .B2(G137), .ZN(new_n457));
  INV_X1    g271(.A(G137), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n458), .A2(KEYINPUT11), .A3(G134), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n258), .A2(G137), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n457), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(G131), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n457), .A2(new_n459), .A3(new_n198), .A4(new_n460), .ZN(new_n463));
  AND2_X1   g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n392), .A2(G128), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n391), .B1(new_n373), .B2(KEYINPUT1), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n402), .B1(new_n467), .B2(new_n383), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n468), .A2(KEYINPUT10), .A3(new_n356), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n384), .A2(new_n385), .ZN(new_n470));
  AOI22_X1  g284(.A1(new_n396), .A2(new_n470), .B1(new_n400), .B2(new_n384), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n332), .A2(new_n471), .A3(new_n349), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n455), .A2(new_n464), .A3(new_n469), .A4(new_n472), .ZN(new_n473));
  XNOR2_X1  g287(.A(G110), .B(G140), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n194), .A2(G227), .ZN(new_n475));
  XOR2_X1   g289(.A(new_n474), .B(new_n475), .Z(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n473), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT82), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n355), .A2(new_n402), .ZN(new_n480));
  INV_X1    g294(.A(new_n465), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n383), .B1(new_n481), .B2(new_n390), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n479), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n397), .A2(KEYINPUT82), .A3(new_n355), .A4(new_n402), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n483), .A2(new_n484), .A3(new_n453), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n462), .A2(new_n463), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT12), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n485), .A2(KEYINPUT12), .A3(new_n486), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n478), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n469), .A2(new_n472), .ZN(new_n492));
  INV_X1    g306(.A(new_n450), .ZN(new_n493));
  OAI21_X1  g307(.A(G128), .B1(new_n389), .B2(KEYINPUT81), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n377), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n355), .B1(new_n495), .B2(new_n402), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n496), .A2(KEYINPUT10), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n486), .B1(new_n492), .B2(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n477), .B1(new_n498), .B2(new_n473), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n445), .B(new_n238), .C1(new_n491), .C2(new_n499), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n492), .A2(new_n497), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n476), .B1(new_n501), .B2(new_n464), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(new_n498), .ZN(new_n503));
  INV_X1    g317(.A(new_n473), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n504), .B1(new_n489), .B2(new_n490), .ZN(new_n505));
  OAI211_X1 g319(.A(G469), .B(new_n503), .C1(new_n505), .C2(new_n477), .ZN(new_n506));
  NAND2_X1  g320(.A1(G469), .A2(G902), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n500), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  OAI21_X1  g322(.A(G221), .B1(new_n267), .B2(G902), .ZN(new_n509));
  AND2_X1   g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AND3_X1   g324(.A1(new_n316), .A2(new_n444), .A3(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT28), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT68), .ZN(new_n513));
  INV_X1    g327(.A(new_n460), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n258), .A2(G137), .ZN(new_n515));
  OAI21_X1  g329(.A(G131), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n463), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n513), .B1(new_n422), .B2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n517), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n468), .A2(KEYINPUT68), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n347), .B1(new_n471), .B2(new_n486), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n518), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n471), .A2(new_n486), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n518), .A2(new_n520), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(new_n347), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT74), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n523), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n525), .A2(KEYINPUT74), .A3(new_n347), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n512), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  OAI22_X1  g344(.A1(new_n422), .A2(new_n517), .B1(new_n464), .B2(new_n387), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n512), .B1(new_n531), .B2(new_n347), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n187), .A2(G210), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n533), .B(KEYINPUT27), .ZN(new_n534));
  XNOR2_X1  g348(.A(KEYINPUT26), .B(G101), .ZN(new_n535));
  XNOR2_X1  g349(.A(new_n534), .B(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n532), .A2(KEYINPUT29), .A3(new_n536), .ZN(new_n537));
  OAI211_X1 g351(.A(KEYINPUT75), .B(new_n238), .C1(new_n530), .C2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT75), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n526), .A2(new_n527), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n540), .A2(new_n522), .A3(new_n529), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n537), .B1(new_n541), .B2(KEYINPUT28), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n539), .B1(new_n542), .B2(G902), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT73), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT69), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT30), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n546), .B1(new_n471), .B2(new_n486), .ZN(new_n547));
  AND3_X1   g361(.A1(new_n518), .A2(new_n520), .A3(new_n547), .ZN(new_n548));
  AOI22_X1  g362(.A1(new_n468), .A2(new_n519), .B1(new_n471), .B2(new_n486), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n347), .B1(new_n549), .B2(KEYINPUT30), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n545), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(new_n347), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n552), .B1(new_n531), .B2(new_n546), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n518), .A2(new_n520), .A3(new_n547), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n553), .A2(KEYINPUT69), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n523), .B1(new_n551), .B2(new_n555), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n544), .B1(new_n556), .B2(new_n536), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n464), .A2(new_n387), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n517), .B1(new_n397), .B2(new_n402), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n546), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  AND4_X1   g374(.A1(KEYINPUT69), .A2(new_n554), .A3(new_n560), .A4(new_n347), .ZN(new_n561));
  AOI21_X1  g375(.A(KEYINPUT69), .B1(new_n553), .B2(new_n554), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n522), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n536), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n563), .A2(KEYINPUT73), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n557), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT29), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n347), .B1(new_n558), .B2(new_n559), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n522), .A2(new_n568), .ZN(new_n569));
  XOR2_X1   g383(.A(KEYINPUT71), .B(KEYINPUT28), .Z(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(KEYINPUT72), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT72), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n569), .A2(new_n574), .A3(new_n571), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n573), .A2(new_n575), .A3(new_n532), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n567), .B1(new_n576), .B2(new_n564), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n538), .B(new_n543), .C1(new_n566), .C2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(G472), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT32), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT31), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n522), .A2(new_n536), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n581), .B(new_n583), .C1(new_n561), .C2(new_n562), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(KEYINPUT70), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n582), .B1(new_n551), .B2(new_n555), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT70), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n586), .A2(new_n587), .A3(new_n581), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n583), .B1(new_n561), .B2(new_n562), .ZN(new_n590));
  AOI22_X1  g404(.A1(new_n576), .A2(new_n564), .B1(new_n590), .B2(KEYINPUT31), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NOR2_X1   g406(.A1(G472), .A2(G902), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n580), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n593), .ZN(new_n595));
  AOI211_X1 g409(.A(KEYINPUT32), .B(new_n595), .C1(new_n589), .C2(new_n591), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n579), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n268), .B1(G234), .B2(new_n238), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT25), .ZN(new_n600));
  XOR2_X1   g414(.A(G119), .B(G128), .Z(new_n601));
  XNOR2_X1  g415(.A(KEYINPUT24), .B(G110), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT23), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n604), .B1(new_n341), .B2(G128), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n251), .A2(KEYINPUT23), .A3(G119), .ZN(new_n606));
  OAI211_X1 g420(.A(new_n605), .B(new_n606), .C1(G119), .C2(new_n251), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n603), .B1(new_n607), .B2(G110), .ZN(new_n608));
  OAI211_X1 g422(.A(new_n212), .B(new_n608), .C1(new_n304), .C2(new_n305), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n210), .A2(new_n212), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n607), .A2(G110), .ZN(new_n611));
  OAI211_X1 g425(.A(new_n610), .B(new_n611), .C1(new_n601), .C2(new_n602), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n194), .A2(G221), .A3(G234), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(KEYINPUT78), .ZN(new_n614));
  XNOR2_X1  g428(.A(KEYINPUT22), .B(G137), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(new_n616));
  AND3_X1   g430(.A1(new_n609), .A2(new_n612), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n616), .B1(new_n609), .B2(new_n612), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n600), .B1(new_n619), .B2(G902), .ZN(new_n620));
  OAI211_X1 g434(.A(KEYINPUT25), .B(new_n238), .C1(new_n617), .C2(new_n618), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n599), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NOR3_X1   g436(.A1(new_n619), .A2(G902), .A3(new_n598), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AND3_X1   g438(.A1(new_n597), .A2(KEYINPUT79), .A3(new_n624), .ZN(new_n625));
  AOI21_X1  g439(.A(KEYINPUT79), .B1(new_n597), .B2(new_n624), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n511), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  XOR2_X1   g441(.A(new_n627), .B(new_n329), .Z(G3));
  INV_X1    g442(.A(new_n317), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n629), .B1(new_n442), .B2(new_n443), .ZN(new_n630));
  INV_X1    g444(.A(G475), .ZN(new_n631));
  AOI21_X1  g445(.A(G902), .B1(new_n233), .B2(new_n236), .ZN(new_n632));
  OAI22_X1  g446(.A1(new_n289), .A2(new_n291), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g447(.A(KEYINPUT93), .B1(new_n274), .B2(G478), .ZN(new_n634));
  INV_X1    g448(.A(new_n273), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n635), .A2(new_n238), .A3(new_n271), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT93), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n636), .A2(new_n637), .A3(new_n275), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT33), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n635), .A2(new_n640), .A3(new_n271), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT91), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n260), .A2(new_n266), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT92), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n644), .A2(new_n645), .A3(new_n270), .ZN(new_n646));
  OAI211_X1 g460(.A(new_n260), .B(new_n266), .C1(KEYINPUT92), .C2(new_n269), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n646), .A2(KEYINPUT33), .A3(new_n647), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n635), .A2(KEYINPUT91), .A3(new_n640), .A4(new_n271), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n275), .A2(G902), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n643), .A2(new_n648), .A3(new_n649), .A4(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n639), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n633), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n653), .A2(new_n301), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n630), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(KEYINPUT94), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT94), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n630), .A2(new_n654), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n592), .A2(new_n593), .ZN(new_n660));
  INV_X1    g474(.A(G472), .ZN(new_n661));
  AOI21_X1  g475(.A(G902), .B1(new_n589), .B2(new_n591), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n660), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n510), .A2(new_n624), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n659), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(KEYINPUT95), .ZN(new_n667));
  XNOR2_X1  g481(.A(KEYINPUT34), .B(G104), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G6));
  INV_X1    g483(.A(new_n630), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n636), .B(new_n276), .ZN(new_n671));
  OAI211_X1 g485(.A(new_n240), .B(new_n671), .C1(new_n289), .C2(new_n291), .ZN(new_n672));
  NOR3_X1   g486(.A1(new_n670), .A2(new_n301), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n665), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(KEYINPUT97), .B(G107), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(KEYINPUT96), .B(KEYINPUT35), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G9));
  NAND2_X1  g492(.A1(new_n609), .A2(new_n612), .ZN(new_n679));
  OR2_X1    g493(.A1(new_n616), .A2(KEYINPUT36), .ZN(new_n680));
  XOR2_X1   g494(.A(new_n679), .B(new_n680), .Z(new_n681));
  AND3_X1   g495(.A1(new_n681), .A2(new_n238), .A3(new_n599), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n622), .A2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n316), .A2(new_n510), .A3(new_n444), .A4(new_n684), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n685), .A2(new_n663), .ZN(new_n686));
  XNOR2_X1  g500(.A(KEYINPUT37), .B(G110), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G12));
  NAND2_X1  g502(.A1(new_n508), .A2(new_n509), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n689), .A2(new_n683), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n295), .B(KEYINPUT98), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(G900), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n692), .B1(new_n693), .B2(new_n296), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  AND4_X1   g509(.A1(new_n671), .A2(new_n630), .A3(new_n313), .A4(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n597), .A2(new_n690), .A3(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(KEYINPUT99), .B(G128), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(G30));
  NOR3_X1   g513(.A1(new_n313), .A2(new_n277), .A3(new_n629), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(new_n683), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n442), .A2(new_n443), .ZN(new_n702));
  XOR2_X1   g516(.A(new_n702), .B(KEYINPUT38), .Z(new_n703));
  INV_X1    g517(.A(KEYINPUT40), .ZN(new_n704));
  XOR2_X1   g518(.A(new_n694), .B(KEYINPUT39), .Z(new_n705));
  AND2_X1   g519(.A1(new_n510), .A2(new_n705), .ZN(new_n706));
  AOI211_X1 g520(.A(new_n701), .B(new_n703), .C1(new_n704), .C2(new_n706), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n556), .A2(new_n564), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n238), .B1(new_n541), .B2(new_n536), .ZN(new_n709));
  OAI21_X1  g523(.A(G472), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(KEYINPUT100), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n711), .B1(new_n594), .B2(new_n596), .ZN(new_n712));
  OAI211_X1 g526(.A(new_n707), .B(new_n712), .C1(new_n704), .C2(new_n706), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G143), .ZN(G45));
  INV_X1    g528(.A(new_n653), .ZN(new_n715));
  AND3_X1   g529(.A1(new_n630), .A2(new_n715), .A3(new_n695), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n597), .A2(new_n690), .A3(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G146), .ZN(G48));
  NAND2_X1  g532(.A1(new_n500), .A2(new_n509), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT102), .ZN(new_n720));
  INV_X1    g534(.A(new_n490), .ZN(new_n721));
  AOI21_X1  g535(.A(KEYINPUT12), .B1(new_n485), .B2(new_n486), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n502), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(new_n499), .ZN(new_n724));
  AOI21_X1  g538(.A(G902), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  OAI21_X1  g539(.A(G469), .B1(new_n725), .B2(KEYINPUT101), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n238), .B1(new_n491), .B2(new_n499), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT101), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n720), .B1(new_n726), .B2(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n445), .B1(new_n727), .B2(new_n728), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n725), .A2(KEYINPUT101), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n731), .A2(KEYINPUT102), .A3(new_n732), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n719), .B1(new_n730), .B2(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n659), .A2(new_n597), .A3(new_n624), .A4(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(KEYINPUT41), .B(G113), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n735), .B(new_n736), .ZN(G15));
  NAND4_X1  g551(.A1(new_n597), .A2(new_n673), .A3(new_n624), .A4(new_n734), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G116), .ZN(G18));
  AOI21_X1  g553(.A(new_n683), .B1(new_n302), .B2(new_n315), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n597), .A2(new_n630), .A3(new_n740), .A4(new_n734), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G119), .ZN(G21));
  INV_X1    g556(.A(KEYINPUT104), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n702), .A2(new_n700), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n744), .A2(new_n301), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n734), .A2(new_n745), .ZN(new_n746));
  AOI22_X1  g560(.A1(new_n585), .A2(new_n588), .B1(KEYINPUT31), .B2(new_n590), .ZN(new_n747));
  INV_X1    g561(.A(new_n532), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n564), .B1(new_n530), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n593), .B(KEYINPUT103), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  OAI211_X1 g566(.A(new_n752), .B(new_n624), .C1(new_n661), .C2(new_n662), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n743), .B1(new_n746), .B2(new_n753), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n661), .B1(new_n592), .B2(new_n238), .ZN(new_n755));
  INV_X1    g569(.A(new_n751), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n756), .B1(new_n747), .B2(new_n749), .ZN(new_n757));
  INV_X1    g571(.A(new_n624), .ZN(new_n758));
  NOR3_X1   g572(.A1(new_n755), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n759), .A2(KEYINPUT104), .A3(new_n734), .A4(new_n745), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n754), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G122), .ZN(G24));
  NOR2_X1   g576(.A1(new_n755), .A2(new_n757), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n763), .A2(new_n716), .A3(new_n734), .A4(new_n684), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G125), .ZN(G27));
  INV_X1    g579(.A(KEYINPUT42), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n597), .A2(new_n624), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n442), .A2(new_n443), .A3(new_n317), .A4(new_n695), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n768), .A2(new_n689), .A3(new_n653), .ZN(new_n769));
  INV_X1    g583(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n766), .B1(new_n767), .B2(new_n770), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n597), .A2(new_n769), .A3(KEYINPUT42), .A4(new_n624), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G131), .ZN(G33));
  INV_X1    g588(.A(KEYINPUT105), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n775), .B1(new_n672), .B2(new_n694), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n313), .A2(KEYINPUT105), .A3(new_n671), .A4(new_n695), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NOR4_X1   g592(.A1(new_n778), .A2(new_n689), .A3(new_n702), .A4(new_n629), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n779), .A2(new_n597), .A3(new_n624), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G134), .ZN(G36));
  AND2_X1   g595(.A1(new_n639), .A2(new_n651), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n633), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(KEYINPUT43), .ZN(new_n784));
  AND3_X1   g598(.A1(new_n663), .A2(new_n684), .A3(new_n784), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n785), .A2(KEYINPUT44), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(KEYINPUT106), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n503), .B1(new_n505), .B2(new_n477), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT45), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n445), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n790), .B1(new_n789), .B2(new_n788), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(new_n507), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT46), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n791), .A2(KEYINPUT46), .A3(new_n507), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n794), .A2(new_n500), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(new_n509), .ZN(new_n797));
  INV_X1    g611(.A(new_n797), .ZN(new_n798));
  AOI211_X1 g612(.A(new_n702), .B(new_n629), .C1(new_n785), .C2(KEYINPUT44), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n787), .A2(new_n705), .A3(new_n798), .A4(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(G137), .ZN(G39));
  NAND2_X1  g615(.A1(new_n798), .A2(KEYINPUT47), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT47), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n797), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  NOR4_X1   g619(.A1(new_n597), .A2(new_n624), .A3(new_n653), .A4(new_n768), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(G140), .ZN(G42));
  INV_X1    g622(.A(new_n509), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n758), .A2(new_n318), .A3(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT107), .ZN(new_n811));
  OR2_X1    g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n810), .A2(new_n811), .ZN(new_n813));
  AND4_X1   g627(.A1(new_n703), .A2(new_n812), .A3(new_n783), .A4(new_n813), .ZN(new_n814));
  AOI22_X1  g628(.A1(new_n730), .A2(new_n733), .B1(new_n445), .B2(new_n725), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(KEYINPUT49), .ZN(new_n816));
  INV_X1    g630(.A(new_n712), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n814), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n683), .A2(new_n695), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n744), .A2(new_n819), .A3(new_n689), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n712), .A2(new_n820), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n697), .A2(new_n717), .A3(new_n821), .A4(new_n764), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n822), .B(KEYINPUT52), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n624), .A2(new_n508), .A3(new_n509), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n824), .B(new_n660), .C1(new_n661), .C2(new_n662), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n672), .A2(KEYINPUT109), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT109), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n313), .A2(new_n827), .A3(new_n671), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n313), .A2(new_n782), .A3(KEYINPUT108), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT108), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n830), .B1(new_n633), .B2(new_n652), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n826), .B(new_n828), .C1(new_n829), .C2(new_n831), .ZN(new_n832));
  AOI211_X1 g646(.A(new_n301), .B(new_n318), .C1(new_n442), .C2(new_n443), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OAI22_X1  g648(.A1(new_n825), .A2(new_n834), .B1(new_n685), .B2(new_n663), .ZN(new_n835));
  INV_X1    g649(.A(new_n734), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n836), .B1(new_n658), .B2(new_n656), .ZN(new_n837));
  INV_X1    g651(.A(new_n767), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n835), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n738), .A2(new_n741), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n839), .A2(new_n627), .A3(new_n840), .A4(new_n761), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT110), .ZN(new_n842));
  OR3_X1    g656(.A1(new_n768), .A2(new_n842), .A3(new_n292), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n842), .B1(new_n768), .B2(new_n292), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n597), .A2(new_n843), .A3(new_n690), .A4(new_n844), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n755), .A2(new_n757), .A3(new_n683), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(new_n769), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n845), .A2(new_n780), .A3(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(new_n773), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT53), .ZN(new_n851));
  NOR4_X1   g665(.A1(new_n823), .A2(new_n841), .A3(new_n850), .A4(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n841), .A2(new_n850), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n697), .A2(new_n764), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n717), .A2(new_n821), .ZN(new_n855));
  AOI21_X1  g669(.A(KEYINPUT52), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT52), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n822), .A2(new_n857), .ZN(new_n858));
  OAI21_X1  g672(.A(KEYINPUT111), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n854), .A2(new_n855), .A3(KEYINPUT52), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT111), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n822), .A2(new_n857), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n853), .A2(new_n859), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n852), .B1(new_n851), .B2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT54), .ZN(new_n866));
  OAI21_X1  g680(.A(KEYINPUT112), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n864), .A2(new_n851), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n860), .A2(new_n862), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n853), .A2(KEYINPUT53), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT112), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n871), .A2(new_n872), .A3(KEYINPUT54), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n867), .A2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(new_n834), .ZN(new_n875));
  AND4_X1   g689(.A1(new_n316), .A2(new_n510), .A3(new_n444), .A4(new_n684), .ZN(new_n876));
  INV_X1    g690(.A(new_n663), .ZN(new_n877));
  AOI22_X1  g691(.A1(new_n875), .A2(new_n665), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n878), .A2(new_n735), .A3(new_n738), .A4(new_n741), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n754), .A2(new_n760), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n848), .B1(new_n771), .B2(new_n772), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n869), .A2(new_n627), .A3(new_n881), .A4(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(new_n851), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n853), .A2(new_n859), .A3(KEYINPUT53), .A4(new_n863), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n884), .A2(new_n885), .A3(new_n866), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(KEYINPUT113), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n784), .A2(new_n692), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(KEYINPUT115), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(new_n759), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n703), .A2(new_n629), .A3(new_n734), .ZN(new_n892));
  OR2_X1    g706(.A1(new_n892), .A2(KEYINPUT118), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(KEYINPUT118), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n891), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT50), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n891), .A2(KEYINPUT50), .A3(new_n893), .A4(new_n894), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n890), .A2(new_n702), .A3(new_n629), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT116), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n509), .B1(new_n815), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n902), .B1(new_n901), .B2(new_n815), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n802), .A2(new_n804), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n900), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n702), .A2(new_n629), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n734), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n758), .A2(new_n295), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n907), .A2(new_n817), .A3(new_n908), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n909), .A2(new_n633), .A3(new_n652), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n889), .A2(new_n907), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n910), .B1(new_n846), .B2(new_n911), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n899), .A2(KEYINPUT51), .A3(new_n905), .A4(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n734), .A2(new_n630), .ZN(new_n914));
  OAI221_X1 g728(.A(new_n293), .B1(new_n909), .B2(new_n653), .C1(new_n890), .C2(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n911), .A2(new_n838), .ZN(new_n916));
  OR2_X1    g730(.A1(new_n916), .A2(KEYINPUT48), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(KEYINPUT48), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n915), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n913), .A2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(new_n905), .ZN(new_n921));
  OR2_X1    g735(.A1(new_n921), .A2(KEYINPUT117), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(KEYINPUT117), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n922), .A2(new_n923), .A3(new_n899), .A4(new_n912), .ZN(new_n924));
  XNOR2_X1  g738(.A(KEYINPUT114), .B(KEYINPUT51), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n920), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AND3_X1   g740(.A1(new_n874), .A2(new_n887), .A3(new_n926), .ZN(new_n927));
  NOR2_X1   g741(.A1(G952), .A2(G953), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n818), .B1(new_n927), .B2(new_n928), .ZN(G75));
  INV_X1    g743(.A(KEYINPUT56), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n884), .A2(new_n885), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(G902), .ZN(new_n932));
  INV_X1    g746(.A(G210), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n930), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n372), .A2(new_n415), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(new_n413), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT55), .ZN(new_n937));
  AND2_X1   g751(.A1(new_n934), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n934), .A2(new_n937), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n194), .A2(G952), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(G51));
  XNOR2_X1  g755(.A(new_n791), .B(KEYINPUT120), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n932), .A2(new_n942), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n507), .B(KEYINPUT57), .Z(new_n944));
  INV_X1    g758(.A(new_n886), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n866), .B1(new_n884), .B2(new_n885), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n944), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n723), .A2(new_n724), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT119), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n943), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n947), .A2(KEYINPUT119), .A3(new_n948), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n940), .B1(new_n951), .B2(new_n952), .ZN(G54));
  INV_X1    g767(.A(new_n940), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT58), .ZN(new_n955));
  NOR3_X1   g769(.A1(new_n932), .A2(new_n955), .A3(new_n631), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n954), .B1(new_n956), .B2(new_n287), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n957), .B1(new_n287), .B2(new_n956), .ZN(G60));
  NAND3_X1  g772(.A1(new_n643), .A2(new_n649), .A3(new_n648), .ZN(new_n959));
  XNOR2_X1  g773(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n275), .A2(new_n238), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n960), .B(new_n961), .Z(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n959), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n964), .B1(new_n945), .B2(new_n946), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(new_n954), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n872), .B1(new_n871), .B2(KEYINPUT54), .ZN(new_n967));
  AOI211_X1 g781(.A(KEYINPUT112), .B(new_n866), .C1(new_n868), .C2(new_n870), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT113), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n886), .B(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n962), .B1(new_n969), .B2(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n966), .B1(new_n972), .B2(new_n959), .ZN(G63));
  NAND2_X1  g787(.A1(G217), .A2(G902), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(KEYINPUT60), .ZN(new_n975));
  INV_X1    g789(.A(new_n975), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n681), .B(KEYINPUT123), .Z(new_n977));
  NAND4_X1  g791(.A1(new_n881), .A2(new_n882), .A3(KEYINPUT53), .A4(new_n627), .ZN(new_n978));
  AND3_X1   g792(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n861), .B1(new_n860), .B2(new_n862), .ZN(new_n980));
  NOR3_X1   g794(.A1(new_n978), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g795(.A(KEYINPUT53), .B1(new_n853), .B2(new_n869), .ZN(new_n982));
  OAI211_X1 g796(.A(new_n976), .B(new_n977), .C1(new_n981), .C2(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT124), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n931), .A2(KEYINPUT124), .A3(new_n976), .A4(new_n977), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n979), .A2(new_n980), .ZN(new_n987));
  INV_X1    g801(.A(new_n978), .ZN(new_n988));
  AOI22_X1  g802(.A1(new_n987), .A2(new_n988), .B1(new_n883), .B2(new_n851), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n619), .B1(new_n989), .B2(new_n975), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n985), .A2(new_n954), .A3(new_n986), .A4(new_n990), .ZN(new_n991));
  AND3_X1   g805(.A1(new_n991), .A2(KEYINPUT122), .A3(KEYINPUT61), .ZN(new_n992));
  AOI21_X1  g806(.A(KEYINPUT61), .B1(new_n991), .B2(KEYINPUT122), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n992), .A2(new_n993), .ZN(G66));
  AOI21_X1  g808(.A(new_n194), .B1(new_n299), .B2(G224), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n995), .B1(new_n841), .B2(new_n194), .ZN(new_n996));
  INV_X1    g810(.A(G898), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n935), .B1(new_n997), .B2(G953), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n996), .B(new_n998), .ZN(G69));
  NAND2_X1  g813(.A1(new_n554), .A2(new_n560), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n1000), .B(KEYINPUT125), .Z(new_n1001));
  XNOR2_X1  g815(.A(new_n1001), .B(new_n283), .ZN(new_n1002));
  INV_X1    g816(.A(new_n1002), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n1003), .B1(G900), .B2(G953), .ZN(new_n1004));
  AND2_X1   g818(.A1(new_n800), .A2(new_n807), .ZN(new_n1005));
  INV_X1    g819(.A(new_n705), .ZN(new_n1006));
  NOR3_X1   g820(.A1(new_n797), .A2(new_n1006), .A3(new_n744), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n838), .B1(new_n1007), .B2(new_n779), .ZN(new_n1008));
  AND3_X1   g822(.A1(new_n773), .A2(new_n717), .A3(new_n854), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n1005), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n1004), .B1(new_n1010), .B2(G953), .ZN(new_n1011));
  INV_X1    g825(.A(new_n1011), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n713), .A2(new_n717), .A3(new_n854), .ZN(new_n1013));
  OR2_X1    g827(.A1(new_n1013), .A2(KEYINPUT62), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1013), .A2(KEYINPUT62), .ZN(new_n1015));
  AND2_X1   g829(.A1(new_n706), .A2(new_n906), .ZN(new_n1016));
  XOR2_X1   g830(.A(new_n832), .B(KEYINPUT126), .Z(new_n1017));
  OAI211_X1 g831(.A(new_n1016), .B(new_n1017), .C1(new_n625), .C2(new_n626), .ZN(new_n1018));
  NAND4_X1  g832(.A1(new_n1005), .A2(new_n1014), .A3(new_n1015), .A4(new_n1018), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n1002), .B1(new_n1019), .B2(new_n194), .ZN(new_n1020));
  NOR2_X1   g834(.A1(new_n1012), .A2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n194), .B1(G227), .B2(G900), .ZN(new_n1022));
  INV_X1    g836(.A(KEYINPUT127), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n1022), .B1(new_n1011), .B2(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g838(.A(new_n1021), .B(new_n1024), .ZN(G72));
  NAND2_X1  g839(.A1(G472), .A2(G902), .ZN(new_n1026));
  XOR2_X1   g840(.A(new_n1026), .B(KEYINPUT63), .Z(new_n1027));
  OAI21_X1  g841(.A(new_n1027), .B1(new_n1019), .B2(new_n841), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n1028), .A2(new_n708), .ZN(new_n1029));
  OAI21_X1  g843(.A(new_n1027), .B1(new_n1010), .B2(new_n841), .ZN(new_n1030));
  NAND3_X1  g844(.A1(new_n1030), .A2(new_n564), .A3(new_n556), .ZN(new_n1031));
  OAI211_X1 g845(.A(new_n871), .B(new_n1027), .C1(new_n586), .C2(new_n566), .ZN(new_n1032));
  AND4_X1   g846(.A1(new_n954), .A2(new_n1029), .A3(new_n1031), .A4(new_n1032), .ZN(G57));
endmodule


