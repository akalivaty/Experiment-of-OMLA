//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 0 0 0 1 1 0 1 1 0 0 0 0 1 1 1 1 1 1 1 1 0 1 1 0 0 1 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 1 0 1 0 0 0 0 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:04 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n723, new_n724,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n788, new_n789, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n976, new_n977, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070;
  XNOR2_X1  g000(.A(G110), .B(G140), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G227), .ZN(new_n189));
  XOR2_X1   g003(.A(new_n187), .B(new_n189), .Z(new_n190));
  INV_X1    g004(.A(KEYINPUT10), .ZN(new_n191));
  INV_X1    g005(.A(G143), .ZN(new_n192));
  OAI21_X1  g006(.A(KEYINPUT66), .B1(new_n192), .B2(G146), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT66), .ZN(new_n194));
  INV_X1    g008(.A(G146), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n194), .A2(new_n195), .A3(G143), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n192), .A2(G146), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n193), .A2(new_n196), .A3(new_n197), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n192), .A2(G146), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT1), .ZN(new_n200));
  OAI21_X1  g014(.A(G128), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n198), .A2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n200), .A2(KEYINPUT67), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT67), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(KEYINPUT1), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n203), .A2(new_n205), .A3(G128), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n202), .B1(new_n198), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G104), .ZN(new_n208));
  OAI21_X1  g022(.A(KEYINPUT3), .B1(new_n208), .B2(G107), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT3), .ZN(new_n210));
  INV_X1    g024(.A(G107), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n210), .A2(new_n211), .A3(G104), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n208), .A2(G107), .ZN(new_n213));
  AND3_X1   g027(.A1(new_n209), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  AND2_X1   g028(.A1(KEYINPUT76), .A2(G101), .ZN(new_n215));
  NOR2_X1   g029(.A1(KEYINPUT76), .A2(G101), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n211), .A2(G104), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(new_n213), .ZN(new_n219));
  AOI22_X1  g033(.A1(new_n214), .A2(new_n217), .B1(G101), .B2(new_n219), .ZN(new_n220));
  AND3_X1   g034(.A1(new_n207), .A2(KEYINPUT78), .A3(new_n220), .ZN(new_n221));
  AOI21_X1  g035(.A(KEYINPUT78), .B1(new_n207), .B2(new_n220), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n191), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT11), .ZN(new_n224));
  INV_X1    g038(.A(G134), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n224), .B1(new_n225), .B2(G137), .ZN(new_n226));
  INV_X1    g040(.A(G137), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n227), .A2(KEYINPUT11), .A3(G134), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n225), .A2(G137), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n226), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G131), .ZN(new_n231));
  INV_X1    g045(.A(G131), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n226), .A2(new_n228), .A3(new_n232), .A4(new_n229), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n217), .A2(new_n209), .A3(new_n212), .A4(new_n213), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n219), .A2(G101), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(KEYINPUT79), .ZN(new_n239));
  INV_X1    g053(.A(G128), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n203), .A2(new_n205), .ZN(new_n241));
  INV_X1    g055(.A(new_n199), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n240), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  OAI21_X1  g057(.A(KEYINPUT65), .B1(new_n192), .B2(G146), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT65), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n245), .A2(new_n195), .A3(G143), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n244), .A2(new_n246), .A3(new_n197), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  OAI22_X1  g062(.A1(new_n243), .A2(new_n248), .B1(new_n198), .B2(new_n206), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT79), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n236), .A2(new_n250), .A3(new_n237), .ZN(new_n251));
  NAND4_X1  g065(.A1(new_n239), .A2(new_n249), .A3(KEYINPUT10), .A4(new_n251), .ZN(new_n252));
  NOR2_X1   g066(.A1(KEYINPUT0), .A2(G128), .ZN(new_n253));
  NAND2_X1  g067(.A1(KEYINPUT0), .A2(G128), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(KEYINPUT64), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT64), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n256), .A2(KEYINPUT0), .A3(G128), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n253), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(new_n247), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT71), .ZN(new_n260));
  INV_X1    g074(.A(new_n254), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n193), .A2(new_n196), .A3(new_n261), .A4(new_n197), .ZN(new_n262));
  AND3_X1   g076(.A1(new_n259), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n260), .B1(new_n259), .B2(new_n262), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n209), .A2(new_n212), .A3(new_n213), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT4), .ZN(new_n267));
  AND2_X1   g081(.A1(new_n267), .A2(G101), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(KEYINPUT77), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT77), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n266), .A2(new_n271), .A3(new_n268), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n267), .B1(new_n266), .B2(G101), .ZN(new_n273));
  AOI22_X1  g087(.A1(new_n270), .A2(new_n272), .B1(new_n273), .B2(new_n236), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n265), .A2(new_n274), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n223), .A2(new_n235), .A3(new_n252), .A4(new_n275), .ZN(new_n276));
  XNOR2_X1  g090(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n277));
  OAI21_X1  g091(.A(G128), .B1(new_n277), .B2(new_n199), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(new_n247), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n198), .A2(new_n206), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n238), .A2(new_n279), .A3(new_n281), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n282), .B1(new_n221), .B2(new_n222), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT12), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n284), .A2(KEYINPUT80), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n285), .A2(KEYINPUT12), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n234), .A2(KEYINPUT80), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  AND3_X1   g103(.A1(new_n283), .A2(new_n287), .A3(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n287), .B1(new_n283), .B2(new_n289), .ZN(new_n291));
  OAI211_X1 g105(.A(KEYINPUT81), .B(new_n276), .C1(new_n290), .C2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n249), .A2(new_n220), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n207), .A2(new_n220), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT78), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n207), .A2(KEYINPUT78), .A3(new_n220), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n294), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n286), .B1(new_n299), .B2(new_n288), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n283), .A2(new_n287), .A3(new_n289), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(KEYINPUT81), .B1(new_n302), .B2(new_n276), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n190), .B1(new_n293), .B2(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(KEYINPUT10), .B1(new_n297), .B2(new_n298), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n259), .A2(new_n262), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(KEYINPUT71), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n259), .A2(new_n260), .A3(new_n262), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n270), .A2(new_n272), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n273), .A2(new_n236), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n252), .B1(new_n309), .B2(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n234), .B1(new_n305), .B2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(new_n190), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n314), .A2(new_n315), .A3(new_n276), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n304), .A2(G469), .A3(new_n316), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n290), .A2(new_n291), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n276), .A2(new_n315), .ZN(new_n319));
  OAI21_X1  g133(.A(KEYINPUT82), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT82), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n302), .A2(new_n321), .A3(new_n315), .A4(new_n276), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n315), .B1(new_n314), .B2(new_n276), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n320), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(G469), .ZN(new_n326));
  INV_X1    g140(.A(G902), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n325), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n326), .A2(new_n327), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n317), .A2(new_n328), .A3(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(G214), .B1(G237), .B2(G902), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(G210), .B1(G237), .B2(G902), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(G125), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(KEYINPUT75), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT75), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(G125), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  OR3_X1    g154(.A1(new_n249), .A2(KEYINPUT85), .A3(new_n340), .ZN(new_n341));
  XNOR2_X1  g155(.A(KEYINPUT75), .B(G125), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n281), .A2(new_n279), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n306), .A2(new_n340), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n343), .A2(new_n344), .A3(KEYINPUT85), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n341), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n188), .A2(G224), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n346), .B(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT5), .ZN(new_n350));
  INV_X1    g164(.A(G119), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(KEYINPUT69), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT69), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(G119), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n352), .A2(new_n354), .A3(G116), .ZN(new_n355));
  INV_X1    g169(.A(G116), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(G119), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT70), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n355), .A2(KEYINPUT70), .A3(new_n357), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n350), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(G113), .B1(new_n355), .B2(KEYINPUT5), .ZN(new_n363));
  OAI21_X1  g177(.A(KEYINPUT83), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(G113), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(KEYINPUT2), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT2), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(G113), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n355), .A2(new_n357), .A3(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n251), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n250), .B1(new_n236), .B2(new_n237), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  AND3_X1   g187(.A1(new_n355), .A2(KEYINPUT70), .A3(new_n357), .ZN(new_n374));
  AOI21_X1  g188(.A(KEYINPUT70), .B1(new_n355), .B2(new_n357), .ZN(new_n375));
  OAI21_X1  g189(.A(KEYINPUT5), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT83), .ZN(new_n377));
  INV_X1    g191(.A(new_n363), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n376), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n364), .A2(new_n370), .A3(new_n373), .A4(new_n379), .ZN(new_n380));
  AND3_X1   g194(.A1(new_n366), .A2(new_n368), .A3(KEYINPUT68), .ZN(new_n381));
  AOI21_X1  g195(.A(KEYINPUT68), .B1(new_n366), .B2(new_n368), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n360), .A2(new_n361), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(new_n370), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(new_n274), .ZN(new_n386));
  XNOR2_X1  g200(.A(G110), .B(G122), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n380), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(KEYINPUT6), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n380), .A2(new_n386), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n387), .A2(KEYINPUT84), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n389), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n390), .A2(KEYINPUT6), .A3(new_n391), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n349), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n347), .A2(KEYINPUT7), .ZN(new_n396));
  AND2_X1   g210(.A1(new_n341), .A2(new_n345), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT7), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n398), .A2(KEYINPUT87), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n396), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n346), .A2(KEYINPUT87), .A3(KEYINPUT7), .A4(new_n347), .ZN(new_n401));
  XOR2_X1   g215(.A(new_n387), .B(KEYINPUT8), .Z(new_n402));
  INV_X1    g216(.A(KEYINPUT86), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n403), .B1(new_n358), .B2(new_n350), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n378), .ZN(new_n405));
  NOR3_X1   g219(.A1(new_n358), .A2(new_n403), .A3(new_n350), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n370), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n402), .B1(new_n407), .B2(new_n220), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n364), .A2(new_n370), .A3(new_n379), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n408), .B1(new_n409), .B2(new_n220), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n400), .A2(new_n388), .A3(new_n401), .A4(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(new_n327), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n335), .B1(new_n395), .B2(new_n412), .ZN(new_n413));
  AND2_X1   g227(.A1(new_n411), .A2(new_n327), .ZN(new_n414));
  AOI22_X1  g228(.A1(new_n388), .A2(KEYINPUT6), .B1(new_n390), .B2(new_n391), .ZN(new_n415));
  INV_X1    g229(.A(new_n394), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n348), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n414), .A2(new_n417), .A3(new_n334), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n333), .B1(new_n413), .B2(new_n418), .ZN(new_n419));
  XNOR2_X1  g233(.A(KEYINPUT9), .B(G234), .ZN(new_n420));
  OAI21_X1  g234(.A(G221), .B1(new_n420), .B2(G902), .ZN(new_n421));
  AND3_X1   g235(.A1(new_n331), .A2(new_n419), .A3(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(G217), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n423), .B1(G234), .B2(new_n327), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n351), .A2(new_n240), .ZN(new_n425));
  XNOR2_X1  g239(.A(KEYINPUT69), .B(G119), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n425), .B1(new_n426), .B2(new_n240), .ZN(new_n427));
  XNOR2_X1  g241(.A(KEYINPUT24), .B(G110), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  OAI211_X1 g244(.A(KEYINPUT23), .B(new_n425), .C1(new_n426), .C2(new_n240), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT23), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n432), .B1(new_n426), .B2(G128), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(G110), .ZN(new_n435));
  INV_X1    g249(.A(G140), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n436), .B1(new_n337), .B2(new_n339), .ZN(new_n437));
  NOR2_X1   g251(.A1(G125), .A2(G140), .ZN(new_n438));
  OAI21_X1  g252(.A(KEYINPUT16), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT16), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n340), .A2(new_n440), .A3(new_n436), .ZN(new_n441));
  AND3_X1   g255(.A1(new_n439), .A2(G146), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(G146), .B1(new_n439), .B2(new_n441), .ZN(new_n443));
  OAI211_X1 g257(.A(new_n430), .B(new_n435), .C1(new_n442), .C2(new_n443), .ZN(new_n444));
  OAI211_X1 g258(.A(new_n428), .B(new_n425), .C1(new_n426), .C2(new_n240), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n445), .B1(new_n434), .B2(G110), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n439), .A2(G146), .A3(new_n441), .ZN(new_n447));
  XNOR2_X1  g261(.A(G125), .B(G140), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(new_n195), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n446), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  XNOR2_X1  g264(.A(KEYINPUT22), .B(G137), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n451), .B(new_n452), .ZN(new_n453));
  AND3_X1   g267(.A1(new_n444), .A2(new_n450), .A3(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n453), .B1(new_n444), .B2(new_n450), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(KEYINPUT25), .B1(new_n456), .B2(new_n327), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT25), .ZN(new_n458));
  NOR4_X1   g272(.A1(new_n454), .A2(new_n455), .A3(new_n458), .A4(G902), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n424), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n456), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n424), .A2(G902), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n460), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT32), .ZN(new_n465));
  NOR2_X1   g279(.A1(G472), .A2(G902), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT31), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n307), .A2(new_n234), .A3(new_n308), .ZN(new_n469));
  INV_X1    g283(.A(new_n229), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n225), .A2(G137), .ZN(new_n471));
  OAI21_X1  g285(.A(G131), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n249), .A2(new_n233), .A3(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n469), .A2(KEYINPUT30), .A3(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT30), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n235), .A2(new_n306), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n472), .A2(new_n233), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n477), .B1(new_n281), .B2(new_n279), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n475), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n474), .A2(new_n385), .A3(new_n479), .ZN(new_n480));
  NOR2_X1   g294(.A1(G237), .A2(G953), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(G210), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n482), .B(KEYINPUT27), .ZN(new_n483));
  XNOR2_X1  g297(.A(KEYINPUT26), .B(G101), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n483), .B(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n385), .A2(KEYINPUT72), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT72), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n384), .A2(new_n487), .A3(new_n370), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n486), .A2(new_n469), .A3(new_n473), .A4(new_n488), .ZN(new_n489));
  AND4_X1   g303(.A1(new_n468), .A2(new_n480), .A3(new_n485), .A4(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n485), .ZN(new_n491));
  AND3_X1   g305(.A1(new_n384), .A2(new_n487), .A3(new_n370), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n487), .B1(new_n384), .B2(new_n370), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n478), .B1(new_n265), .B2(new_n234), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n491), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n468), .B1(new_n496), .B2(new_n480), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n490), .A2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT28), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n473), .B1(new_n235), .B2(new_n306), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(new_n385), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n499), .B1(new_n489), .B2(new_n501), .ZN(new_n502));
  AOI21_X1  g316(.A(KEYINPUT28), .B1(new_n494), .B2(new_n495), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n491), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n467), .B1(new_n498), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n465), .B1(new_n505), .B2(KEYINPUT73), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n480), .A2(new_n485), .A3(new_n489), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(KEYINPUT31), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n496), .A2(new_n468), .A3(new_n480), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n504), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(new_n466), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT73), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n511), .A2(new_n512), .A3(KEYINPUT32), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n506), .A2(new_n513), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n502), .A2(new_n503), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT74), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n515), .A2(new_n516), .A3(new_n485), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n489), .A2(new_n499), .ZN(new_n518));
  AOI22_X1  g332(.A1(new_n494), .A2(new_n495), .B1(new_n385), .B2(new_n500), .ZN(new_n519));
  OAI211_X1 g333(.A(new_n485), .B(new_n518), .C1(new_n519), .C2(new_n499), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(KEYINPUT74), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n480), .A2(new_n489), .ZN(new_n522));
  AOI21_X1  g336(.A(KEYINPUT29), .B1(new_n522), .B2(new_n491), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n517), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  AOI22_X1  g338(.A1(new_n486), .A2(new_n488), .B1(new_n469), .B2(new_n473), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(new_n489), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n503), .B1(new_n527), .B2(KEYINPUT28), .ZN(new_n528));
  AND2_X1   g342(.A1(new_n485), .A2(KEYINPUT29), .ZN(new_n529));
  AOI21_X1  g343(.A(G902), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n524), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(G472), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n464), .B1(new_n514), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n439), .A2(new_n441), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(new_n195), .ZN(new_n535));
  AND2_X1   g349(.A1(KEYINPUT88), .A2(G143), .ZN(new_n536));
  NOR2_X1   g350(.A1(KEYINPUT88), .A2(G143), .ZN(new_n537));
  OAI211_X1 g351(.A(G214), .B(new_n481), .C1(new_n536), .C2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(G237), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n539), .A2(new_n188), .A3(G214), .ZN(new_n540));
  NAND2_X1  g354(.A1(KEYINPUT88), .A2(G143), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n538), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(G131), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT17), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n538), .A2(new_n232), .A3(new_n542), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n232), .B1(new_n538), .B2(new_n542), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(KEYINPUT17), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n535), .A2(new_n547), .A3(new_n447), .A4(new_n549), .ZN(new_n550));
  XOR2_X1   g364(.A(G113), .B(G122), .Z(new_n551));
  XOR2_X1   g365(.A(KEYINPUT91), .B(G104), .Z(new_n552));
  XOR2_X1   g366(.A(new_n551), .B(new_n552), .Z(new_n553));
  INV_X1    g367(.A(new_n438), .ZN(new_n554));
  OAI211_X1 g368(.A(G146), .B(new_n554), .C1(new_n342), .C2(new_n436), .ZN(new_n555));
  AOI22_X1  g369(.A1(new_n548), .A2(KEYINPUT18), .B1(new_n555), .B2(new_n449), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT18), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n538), .B(new_n542), .C1(new_n557), .C2(new_n232), .ZN(new_n558));
  AND2_X1   g372(.A1(new_n558), .A2(KEYINPUT89), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n558), .A2(KEYINPUT89), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n556), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  AND3_X1   g375(.A1(new_n550), .A2(new_n553), .A3(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT90), .ZN(new_n563));
  INV_X1    g377(.A(new_n546), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n563), .B1(new_n564), .B2(new_n548), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n544), .A2(KEYINPUT90), .A3(new_n546), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT19), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n448), .A2(new_n567), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n554), .B1(new_n342), .B2(new_n436), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n195), .B(new_n568), .C1(new_n569), .C2(new_n567), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n565), .A2(new_n566), .A3(new_n447), .A4(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n553), .B1(new_n571), .B2(new_n561), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n562), .A2(new_n572), .ZN(new_n573));
  NOR2_X1   g387(.A1(G475), .A2(G902), .ZN(new_n574));
  XOR2_X1   g388(.A(new_n574), .B(KEYINPUT92), .Z(new_n575));
  OAI21_X1  g389(.A(KEYINPUT20), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT20), .ZN(new_n577));
  INV_X1    g391(.A(new_n575), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n577), .B(new_n578), .C1(new_n562), .C2(new_n572), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n553), .B1(new_n550), .B2(new_n561), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n327), .B1(new_n562), .B2(new_n580), .ZN(new_n581));
  AOI22_X1  g395(.A1(new_n576), .A2(new_n579), .B1(G475), .B2(new_n581), .ZN(new_n582));
  NOR3_X1   g396(.A1(new_n420), .A2(new_n423), .A3(G953), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(G122), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(G116), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n356), .A2(G122), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(KEYINPUT93), .ZN(new_n589));
  XNOR2_X1  g403(.A(G116), .B(G122), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT93), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n211), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n356), .A2(KEYINPUT14), .A3(G122), .ZN(new_n595));
  OAI211_X1 g409(.A(G107), .B(new_n595), .C1(new_n588), .C2(KEYINPUT14), .ZN(new_n596));
  XNOR2_X1  g410(.A(G128), .B(G143), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n597), .B(new_n225), .ZN(new_n598));
  AND3_X1   g412(.A1(new_n594), .A2(new_n596), .A3(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n589), .A2(new_n592), .A3(G107), .ZN(new_n600));
  AOI21_X1  g414(.A(KEYINPUT13), .B1(new_n240), .B2(G143), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n601), .A2(new_n225), .ZN(new_n602));
  OR2_X1    g416(.A1(new_n602), .A2(new_n597), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n597), .ZN(new_n604));
  AOI22_X1  g418(.A1(new_n594), .A2(new_n600), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n584), .B1(new_n599), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n594), .A2(new_n600), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n603), .A2(new_n604), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n594), .A2(new_n596), .A3(new_n598), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n609), .A2(new_n610), .A3(new_n583), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n606), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n327), .ZN(new_n613));
  INV_X1    g427(.A(G478), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n614), .A2(KEYINPUT15), .ZN(new_n615));
  XOR2_X1   g429(.A(new_n613), .B(new_n615), .Z(new_n616));
  NAND2_X1  g430(.A1(new_n582), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(G234), .A2(G237), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n618), .A2(G952), .A3(new_n188), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n618), .A2(G902), .A3(G953), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(KEYINPUT21), .B(G898), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n620), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n617), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n422), .A2(new_n533), .A3(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n217), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G3));
  INV_X1    g442(.A(new_n624), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n614), .A2(G902), .ZN(new_n630));
  AOI21_X1  g444(.A(KEYINPUT33), .B1(new_n612), .B2(KEYINPUT95), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT95), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT33), .ZN(new_n633));
  AOI211_X1 g447(.A(new_n632), .B(new_n633), .C1(new_n606), .C2(new_n611), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n630), .B1(new_n631), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n613), .A2(new_n614), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n638), .A2(new_n582), .ZN(new_n639));
  AND3_X1   g453(.A1(new_n419), .A2(new_n629), .A3(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n421), .ZN(new_n641));
  INV_X1    g455(.A(new_n316), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n276), .B1(new_n290), .B2(new_n291), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT81), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n292), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n642), .B1(new_n646), .B2(new_n190), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n329), .B1(new_n647), .B2(G469), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n641), .B1(new_n648), .B2(new_n328), .ZN(new_n649));
  INV_X1    g463(.A(G472), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n650), .B1(new_n510), .B2(new_n327), .ZN(new_n651));
  OR2_X1    g465(.A1(new_n651), .A2(KEYINPUT94), .ZN(new_n652));
  OAI21_X1  g466(.A(KEYINPUT94), .B1(new_n651), .B2(new_n505), .ZN(new_n653));
  AND2_X1   g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n464), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n640), .A2(new_n649), .A3(new_n654), .A4(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT34), .B(G104), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G6));
  XNOR2_X1  g472(.A(new_n613), .B(new_n615), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n582), .A2(new_n629), .A3(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT96), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n581), .A2(G475), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n550), .A2(new_n561), .A3(new_n553), .ZN(new_n664));
  AND2_X1   g478(.A1(new_n571), .A2(new_n561), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n664), .B1(new_n665), .B2(new_n553), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n577), .B1(new_n666), .B2(new_n578), .ZN(new_n667));
  INV_X1    g481(.A(new_n579), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n663), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n669), .A2(new_n616), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n670), .A2(KEYINPUT96), .A3(new_n629), .ZN(new_n671));
  AND3_X1   g485(.A1(new_n419), .A2(new_n662), .A3(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n672), .A2(new_n649), .A3(new_n654), .A4(new_n655), .ZN(new_n673));
  XOR2_X1   g487(.A(KEYINPUT35), .B(G107), .Z(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G9));
  NAND2_X1  g489(.A1(new_n444), .A2(new_n450), .ZN(new_n676));
  INV_X1    g490(.A(new_n453), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n677), .A2(KEYINPUT36), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n676), .B(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(new_n462), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n460), .A2(new_n680), .ZN(new_n681));
  AND3_X1   g495(.A1(new_n652), .A2(new_n653), .A3(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n422), .A2(new_n625), .A3(new_n682), .ZN(new_n683));
  XOR2_X1   g497(.A(KEYINPUT37), .B(G110), .Z(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G12));
  INV_X1    g499(.A(G900), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n622), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(new_n619), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n670), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(KEYINPUT97), .ZN(new_n690));
  INV_X1    g504(.A(new_n681), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n691), .B1(new_n514), .B2(new_n532), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n422), .A2(new_n690), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G128), .ZN(G30));
  INV_X1    g508(.A(KEYINPUT40), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n688), .B(KEYINPUT39), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n331), .A2(new_n421), .A3(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT99), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n331), .A2(KEYINPUT99), .A3(new_n421), .A4(new_n696), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n695), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n699), .A2(new_n695), .A3(new_n700), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n413), .A2(new_n418), .ZN(new_n704));
  XNOR2_X1  g518(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n413), .A2(new_n418), .A3(new_n705), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n522), .A2(new_n485), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n526), .A2(new_n491), .A3(new_n489), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(new_n327), .ZN(new_n714));
  OAI21_X1  g528(.A(G472), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n514), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n669), .A2(new_n659), .ZN(new_n717));
  NOR3_X1   g531(.A1(new_n681), .A2(new_n717), .A3(new_n333), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n710), .A2(new_n716), .A3(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(new_n719), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n702), .A2(new_n703), .A3(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G143), .ZN(G45));
  NAND3_X1  g536(.A1(new_n669), .A2(new_n637), .A3(new_n688), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n422), .A2(new_n692), .A3(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G146), .ZN(G48));
  OAI211_X1 g540(.A(new_n315), .B(new_n276), .C1(new_n290), .C2(new_n291), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n323), .B1(new_n727), .B2(KEYINPUT82), .ZN(new_n728));
  AOI21_X1  g542(.A(G902), .B1(new_n728), .B2(new_n322), .ZN(new_n729));
  AOI21_X1  g543(.A(KEYINPUT100), .B1(new_n729), .B2(new_n326), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n325), .A2(new_n327), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(G469), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n731), .A2(KEYINPUT100), .A3(G469), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n641), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n735), .A2(new_n533), .A3(new_n640), .ZN(new_n736));
  XNOR2_X1  g550(.A(KEYINPUT41), .B(G113), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n736), .B(new_n737), .ZN(G15));
  NAND3_X1  g552(.A1(new_n735), .A2(new_n533), .A3(new_n672), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G116), .ZN(G18));
  NAND4_X1  g554(.A1(new_n735), .A2(new_n419), .A3(new_n625), .A4(new_n692), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G119), .ZN(G21));
  AOI211_X1 g556(.A(new_n333), .B(new_n717), .C1(new_n413), .C2(new_n418), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n508), .A2(new_n509), .ZN(new_n744));
  INV_X1    g558(.A(new_n489), .ZN(new_n745));
  OAI21_X1  g559(.A(KEYINPUT28), .B1(new_n745), .B2(new_n525), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n485), .B1(new_n746), .B2(new_n518), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n466), .B1(new_n744), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n510), .A2(new_n327), .ZN(new_n749));
  XOR2_X1   g563(.A(KEYINPUT101), .B(G472), .Z(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n655), .A2(new_n748), .A3(new_n751), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n752), .A2(new_n624), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n735), .A2(new_n743), .A3(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G122), .ZN(G24));
  NAND2_X1  g569(.A1(new_n723), .A2(KEYINPUT103), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT103), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n669), .A2(new_n637), .A3(new_n757), .A4(new_n688), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  AOI21_X1  g573(.A(G902), .B1(new_n498), .B2(new_n504), .ZN(new_n760));
  INV_X1    g574(.A(new_n750), .ZN(new_n761));
  OAI211_X1 g575(.A(new_n681), .B(new_n748), .C1(new_n760), .C2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT102), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n751), .A2(KEYINPUT102), .A3(new_n681), .A4(new_n748), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n759), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n735), .A2(new_n766), .A3(new_n419), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G125), .ZN(G27));
  NAND2_X1  g582(.A1(new_n331), .A2(new_n421), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT104), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n704), .A2(new_n333), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n331), .A2(KEYINPUT104), .A3(new_n421), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n771), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n505), .A2(KEYINPUT32), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT105), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n776), .B1(new_n505), .B2(KEYINPUT32), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n511), .A2(KEYINPUT105), .A3(new_n465), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n532), .A2(new_n775), .A3(new_n777), .A4(new_n778), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n779), .A2(new_n655), .A3(new_n756), .A4(new_n758), .ZN(new_n780));
  OAI21_X1  g594(.A(KEYINPUT42), .B1(new_n774), .B2(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n413), .A2(new_n418), .A3(new_n332), .ZN(new_n782));
  AOI211_X1 g596(.A(new_n464), .B(new_n782), .C1(new_n514), .C2(new_n532), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n759), .A2(KEYINPUT42), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n783), .A2(new_n771), .A3(new_n773), .A4(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n781), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(new_n232), .ZN(G33));
  NAND4_X1  g601(.A1(new_n783), .A2(new_n690), .A3(new_n771), .A4(new_n773), .ZN(new_n788));
  XOR2_X1   g602(.A(KEYINPUT106), .B(G134), .Z(new_n789));
  XNOR2_X1  g603(.A(new_n788), .B(new_n789), .ZN(G36));
  NAND2_X1  g604(.A1(new_n582), .A2(new_n637), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(KEYINPUT43), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT43), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n582), .A2(new_n637), .A3(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n792), .A2(new_n681), .A3(new_n794), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n654), .A2(new_n795), .ZN(new_n796));
  OR2_X1    g610(.A1(new_n796), .A2(KEYINPUT44), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(KEYINPUT44), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n797), .A2(new_n772), .A3(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(new_n328), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n304), .A2(KEYINPUT45), .A3(new_n316), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(KEYINPUT107), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT107), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n647), .A2(new_n803), .A3(KEYINPUT45), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(new_n647), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT45), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n326), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n805), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(new_n330), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT46), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n800), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n329), .B1(new_n805), .B2(new_n808), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n813), .A2(KEYINPUT46), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n641), .B1(new_n812), .B2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT108), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n815), .A2(new_n816), .A3(new_n696), .ZN(new_n817));
  OAI21_X1  g631(.A(G469), .B1(new_n647), .B2(KEYINPUT45), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n818), .B1(new_n802), .B2(new_n804), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n811), .B1(new_n819), .B2(new_n329), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n814), .A2(new_n820), .A3(new_n328), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n821), .A2(new_n421), .A3(new_n696), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(KEYINPUT108), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n799), .B1(new_n817), .B2(new_n823), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(new_n227), .ZN(G39));
  NAND4_X1  g639(.A1(new_n514), .A2(new_n532), .A3(new_n464), .A4(new_n724), .ZN(new_n826));
  INV_X1    g640(.A(new_n826), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n328), .B1(new_n813), .B2(KEYINPUT46), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n819), .A2(new_n811), .A3(new_n329), .ZN(new_n829));
  OAI211_X1 g643(.A(KEYINPUT47), .B(new_n421), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(new_n830), .ZN(new_n831));
  AOI21_X1  g645(.A(KEYINPUT47), .B1(new_n821), .B2(new_n421), .ZN(new_n832));
  OAI211_X1 g646(.A(new_n772), .B(new_n827), .C1(new_n831), .C2(new_n832), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n833), .B(G140), .ZN(G42));
  NAND2_X1  g648(.A1(new_n733), .A2(new_n734), .ZN(new_n835));
  XNOR2_X1  g649(.A(new_n835), .B(KEYINPUT49), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n655), .A2(new_n332), .A3(new_n421), .ZN(new_n837));
  NOR4_X1   g651(.A1(new_n710), .A2(new_n716), .A3(new_n791), .A4(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n735), .A2(new_n772), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n792), .A2(new_n620), .A3(new_n794), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n779), .A2(new_n655), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g658(.A(KEYINPUT118), .B(KEYINPUT48), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(new_n715), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n847), .B1(new_n506), .B2(new_n513), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n848), .A2(new_n655), .A3(new_n620), .ZN(new_n849));
  OAI21_X1  g663(.A(KEYINPUT115), .B1(new_n840), .B2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(new_n849), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT115), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n851), .A2(new_n852), .A3(new_n735), .A4(new_n772), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n850), .A2(new_n639), .A3(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT118), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n842), .A2(new_n855), .A3(KEYINPUT48), .A4(new_n843), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n841), .A2(new_n752), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n735), .A2(new_n419), .A3(new_n857), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n858), .A2(G952), .A3(new_n188), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n846), .A2(new_n854), .A3(new_n856), .A4(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n857), .A2(new_n772), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n831), .A2(new_n832), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n835), .A2(new_n641), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n861), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n857), .A2(new_n709), .A3(new_n333), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n835), .A2(new_n421), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT50), .ZN(new_n867));
  OR3_X1    g681(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n867), .B1(new_n865), .B2(new_n866), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n850), .A2(new_n582), .A3(new_n638), .A4(new_n853), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n764), .A2(new_n765), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n842), .A2(new_n872), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n870), .A2(new_n871), .A3(KEYINPUT51), .A4(new_n873), .ZN(new_n874));
  OAI21_X1  g688(.A(KEYINPUT117), .B1(new_n864), .B2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(new_n874), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT117), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n821), .A2(new_n421), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT47), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n880), .A2(new_n830), .A3(new_n863), .ZN(new_n881));
  OAI211_X1 g695(.A(new_n876), .B(new_n877), .C1(new_n881), .C2(new_n861), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n860), .B1(new_n875), .B2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT116), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n870), .A2(new_n871), .A3(new_n873), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n863), .B(KEYINPUT114), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n880), .A2(new_n830), .A3(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(new_n861), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n885), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n884), .B1(new_n889), .B2(KEYINPUT51), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT51), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n861), .B1(new_n862), .B2(new_n886), .ZN(new_n892));
  OAI211_X1 g706(.A(KEYINPUT116), .B(new_n891), .C1(new_n892), .C2(new_n885), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n883), .A2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT54), .ZN(new_n896));
  AND2_X1   g710(.A1(new_n767), .A2(new_n693), .ZN(new_n897));
  INV_X1    g711(.A(new_n688), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n681), .A2(new_n898), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n649), .A2(new_n716), .A3(new_n743), .A4(new_n899), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n725), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n897), .A2(KEYINPUT52), .A3(new_n901), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n767), .A2(new_n693), .A3(new_n725), .A4(new_n900), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT52), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n769), .A2(new_n617), .A3(new_n898), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n907), .A2(new_n692), .A3(new_n772), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n771), .A2(new_n766), .A3(new_n772), .A4(new_n773), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n788), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n786), .A2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT109), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n912), .B1(new_n669), .B2(new_n616), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n670), .A2(KEYINPUT109), .ZN(new_n914));
  AND4_X1   g728(.A1(new_n419), .A2(new_n629), .A3(new_n913), .A4(new_n914), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n915), .A2(new_n649), .A3(new_n655), .A4(new_n654), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n741), .A2(new_n739), .A3(new_n754), .A4(new_n916), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n736), .A2(new_n626), .A3(new_n683), .A4(new_n656), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  AND4_X1   g733(.A1(KEYINPUT53), .A2(new_n906), .A3(new_n911), .A4(new_n919), .ZN(new_n920));
  XOR2_X1   g734(.A(KEYINPUT111), .B(KEYINPUT52), .Z(new_n921));
  NAND2_X1  g735(.A1(new_n767), .A2(new_n693), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n725), .A2(new_n900), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n921), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT112), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n903), .A2(KEYINPUT112), .A3(new_n921), .ZN(new_n927));
  OAI21_X1  g741(.A(KEYINPUT110), .B1(new_n903), .B2(new_n904), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT110), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n897), .A2(new_n901), .A3(new_n929), .A4(KEYINPUT52), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n926), .A2(new_n927), .A3(new_n928), .A4(new_n930), .ZN(new_n931));
  NOR4_X1   g745(.A1(new_n786), .A2(new_n910), .A3(new_n917), .A4(new_n918), .ZN(new_n932));
  AOI21_X1  g746(.A(KEYINPUT53), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n920), .B1(new_n933), .B2(KEYINPUT113), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT113), .ZN(new_n935));
  INV_X1    g749(.A(new_n786), .ZN(new_n936));
  INV_X1    g750(.A(new_n910), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n936), .A2(new_n919), .A3(new_n937), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n930), .A2(new_n928), .ZN(new_n939));
  AND3_X1   g753(.A1(new_n903), .A2(KEYINPUT112), .A3(new_n921), .ZN(new_n940));
  AOI21_X1  g754(.A(KEYINPUT112), .B1(new_n903), .B2(new_n921), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n938), .B1(new_n939), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n935), .B1(new_n943), .B2(KEYINPUT53), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n896), .B1(new_n934), .B2(new_n944), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n931), .A2(KEYINPUT53), .A3(new_n932), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT53), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n902), .A2(new_n905), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n947), .B1(new_n938), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n946), .A2(new_n949), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n950), .A2(KEYINPUT54), .ZN(new_n951));
  NOR3_X1   g765(.A1(new_n895), .A2(new_n945), .A3(new_n951), .ZN(new_n952));
  NOR2_X1   g766(.A1(G952), .A2(G953), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n839), .B1(new_n952), .B2(new_n953), .ZN(G75));
  NOR2_X1   g768(.A1(new_n188), .A2(G952), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n327), .B1(new_n946), .B2(new_n949), .ZN(new_n957));
  AOI21_X1  g771(.A(KEYINPUT56), .B1(new_n957), .B2(G210), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n415), .A2(new_n416), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(new_n348), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(KEYINPUT55), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n956), .B1(new_n958), .B2(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT119), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n957), .A2(new_n963), .A3(G210), .ZN(new_n964));
  XNOR2_X1  g778(.A(KEYINPUT120), .B(KEYINPUT56), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n961), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n957), .A2(G210), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n966), .B1(new_n967), .B2(KEYINPUT119), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n962), .B1(new_n964), .B2(new_n968), .ZN(G51));
  AOI21_X1  g783(.A(new_n896), .B1(new_n946), .B2(new_n949), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n951), .A2(new_n970), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n329), .B(KEYINPUT57), .Z(new_n972));
  OAI21_X1  g786(.A(new_n325), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n957), .A2(new_n819), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n955), .B1(new_n973), .B2(new_n974), .ZN(G54));
  AND3_X1   g789(.A1(new_n957), .A2(KEYINPUT58), .A3(G475), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n956), .B1(new_n976), .B2(new_n666), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n977), .B1(new_n666), .B2(new_n976), .ZN(G60));
  OR2_X1    g792(.A1(new_n631), .A2(new_n634), .ZN(new_n979));
  NAND2_X1  g793(.A1(G478), .A2(G902), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n980), .B(KEYINPUT59), .Z(new_n981));
  INV_X1    g795(.A(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n979), .A2(new_n982), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n956), .B1(new_n971), .B2(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(new_n979), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n982), .B1(new_n945), .B2(new_n951), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n984), .B1(new_n985), .B2(new_n986), .ZN(G63));
  NAND2_X1  g801(.A1(G217), .A2(G902), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n988), .B(KEYINPUT60), .Z(new_n989));
  NAND2_X1  g803(.A1(new_n950), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(new_n461), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n950), .A2(new_n679), .A3(new_n989), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n991), .A2(new_n956), .A3(new_n992), .ZN(new_n993));
  INV_X1    g807(.A(KEYINPUT61), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n991), .A2(KEYINPUT61), .A3(new_n956), .A4(new_n992), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n995), .A2(new_n996), .ZN(G66));
  INV_X1    g811(.A(G224), .ZN(new_n998));
  OAI21_X1  g812(.A(G953), .B1(new_n623), .B2(new_n998), .ZN(new_n999));
  INV_X1    g813(.A(KEYINPUT121), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n919), .A2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g815(.A(KEYINPUT121), .B1(new_n917), .B2(new_n918), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n999), .B1(new_n1003), .B2(G953), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n959), .B1(G898), .B2(new_n188), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1005), .B(KEYINPUT122), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n1004), .B(new_n1006), .ZN(G69));
  NAND2_X1  g821(.A1(new_n827), .A2(new_n772), .ZN(new_n1008));
  NOR2_X1   g822(.A1(new_n862), .A2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n1009), .A2(new_n824), .ZN(new_n1010));
  INV_X1    g824(.A(new_n783), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n699), .A2(new_n700), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n639), .B1(new_n914), .B2(new_n913), .ZN(new_n1013));
  NOR3_X1   g827(.A1(new_n1011), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g828(.A(KEYINPUT62), .ZN(new_n1015));
  AND3_X1   g829(.A1(new_n699), .A2(new_n695), .A3(new_n700), .ZN(new_n1016));
  NOR3_X1   g830(.A1(new_n1016), .A2(new_n701), .A3(new_n719), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n767), .A2(new_n693), .A3(new_n725), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n1015), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g833(.A(new_n1018), .ZN(new_n1020));
  NAND3_X1  g834(.A1(new_n721), .A2(KEYINPUT62), .A3(new_n1020), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n1014), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1010), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n474), .A2(new_n479), .ZN(new_n1024));
  XOR2_X1   g838(.A(new_n1024), .B(KEYINPUT123), .Z(new_n1025));
  OAI21_X1  g839(.A(new_n568), .B1(new_n569), .B2(new_n567), .ZN(new_n1026));
  XNOR2_X1  g840(.A(new_n1025), .B(new_n1026), .ZN(new_n1027));
  AND2_X1   g841(.A1(new_n1027), .A2(new_n188), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n1023), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g843(.A1(new_n936), .A2(new_n788), .A3(new_n1020), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n817), .A2(new_n823), .ZN(new_n1031));
  AND2_X1   g845(.A1(new_n843), .A2(new_n743), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n1030), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g847(.A(G953), .B1(new_n1010), .B2(new_n1033), .ZN(new_n1034));
  NOR2_X1   g848(.A1(new_n188), .A2(G900), .ZN(new_n1035));
  XNOR2_X1  g849(.A(new_n1035), .B(KEYINPUT125), .ZN(new_n1036));
  OR2_X1    g850(.A1(new_n1027), .A2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g851(.A(new_n1029), .B1(new_n1034), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g852(.A(KEYINPUT124), .ZN(new_n1039));
  AOI21_X1  g853(.A(new_n188), .B1(G227), .B2(G900), .ZN(new_n1040));
  AND3_X1   g854(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  AOI21_X1  g855(.A(new_n1040), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1042));
  NOR2_X1   g856(.A1(new_n1041), .A2(new_n1042), .ZN(G72));
  NOR2_X1   g857(.A1(new_n522), .A2(new_n485), .ZN(new_n1044));
  INV_X1    g858(.A(new_n1044), .ZN(new_n1045));
  NAND2_X1  g859(.A1(G472), .A2(G902), .ZN(new_n1046));
  XOR2_X1   g860(.A(new_n1046), .B(KEYINPUT63), .Z(new_n1047));
  AND3_X1   g861(.A1(new_n1045), .A2(new_n711), .A3(new_n1047), .ZN(new_n1048));
  NAND2_X1  g862(.A1(new_n931), .A2(new_n932), .ZN(new_n1049));
  NAND3_X1  g863(.A1(new_n1049), .A2(KEYINPUT113), .A3(new_n947), .ZN(new_n1050));
  INV_X1    g864(.A(new_n920), .ZN(new_n1051));
  NAND2_X1  g865(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NOR2_X1   g866(.A1(new_n933), .A2(KEYINPUT113), .ZN(new_n1053));
  OAI21_X1  g867(.A(new_n1048), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g868(.A(KEYINPUT126), .ZN(new_n1055));
  INV_X1    g869(.A(new_n799), .ZN(new_n1056));
  AOI21_X1  g870(.A(new_n816), .B1(new_n815), .B2(new_n696), .ZN(new_n1057));
  NOR2_X1   g871(.A1(new_n822), .A2(KEYINPUT108), .ZN(new_n1058));
  OAI21_X1  g872(.A(new_n1056), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  NAND4_X1  g873(.A1(new_n1022), .A2(new_n1059), .A3(new_n833), .A4(new_n1003), .ZN(new_n1060));
  NAND2_X1  g874(.A1(new_n1060), .A2(new_n1047), .ZN(new_n1061));
  AOI21_X1  g875(.A(new_n1055), .B1(new_n1061), .B2(new_n712), .ZN(new_n1062));
  AOI211_X1 g876(.A(KEYINPUT126), .B(new_n711), .C1(new_n1060), .C2(new_n1047), .ZN(new_n1063));
  OAI21_X1  g877(.A(new_n1054), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g878(.A(KEYINPUT127), .ZN(new_n1065));
  NAND3_X1  g879(.A1(new_n1010), .A2(new_n1003), .A3(new_n1033), .ZN(new_n1066));
  AOI21_X1  g880(.A(new_n1045), .B1(new_n1066), .B2(new_n1047), .ZN(new_n1067));
  OAI21_X1  g881(.A(new_n1065), .B1(new_n1067), .B2(new_n955), .ZN(new_n1068));
  AND2_X1   g882(.A1(new_n1066), .A2(new_n1047), .ZN(new_n1069));
  OAI211_X1 g883(.A(KEYINPUT127), .B(new_n956), .C1(new_n1069), .C2(new_n1045), .ZN(new_n1070));
  AOI21_X1  g884(.A(new_n1064), .B1(new_n1068), .B2(new_n1070), .ZN(G57));
endmodule


