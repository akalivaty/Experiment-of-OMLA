//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 0 0 0 1 1 0 0 1 0 1 1 0 1 1 0 1 0 1 0 1 0 1 0 0 1 0 0 0 0 0 0 0 0 0 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:58 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT11), .ZN(new_n188));
  INV_X1    g002(.A(G134), .ZN(new_n189));
  OAI21_X1  g003(.A(new_n188), .B1(new_n189), .B2(G137), .ZN(new_n190));
  INV_X1    g004(.A(G137), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(KEYINPUT11), .A3(G134), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n189), .A2(G137), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n190), .A2(new_n192), .A3(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G131), .ZN(new_n195));
  INV_X1    g009(.A(G131), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n190), .A2(new_n192), .A3(new_n196), .A4(new_n193), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n195), .A2(KEYINPUT66), .A3(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G143), .ZN(new_n199));
  OAI21_X1  g013(.A(KEYINPUT64), .B1(new_n199), .B2(G146), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g015(.A(G146), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n201), .A2(new_n202), .A3(G143), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n199), .A2(G146), .ZN(new_n204));
  NAND2_X1  g018(.A1(KEYINPUT0), .A2(G128), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  AND4_X1   g020(.A1(new_n200), .A2(new_n203), .A3(new_n204), .A4(new_n206), .ZN(new_n207));
  OR2_X1    g021(.A1(KEYINPUT0), .A2(G128), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(new_n205), .ZN(new_n209));
  XNOR2_X1  g023(.A(G143), .B(G146), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n207), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT66), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n194), .A2(new_n213), .A3(G131), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n198), .A2(new_n212), .A3(new_n214), .ZN(new_n215));
  XNOR2_X1  g029(.A(G116), .B(G119), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  XNOR2_X1  g031(.A(KEYINPUT2), .B(G113), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  XOR2_X1   g033(.A(KEYINPUT2), .B(G113), .Z(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(new_n216), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n219), .A2(new_n221), .A3(KEYINPUT69), .ZN(new_n222));
  OR3_X1    g036(.A1(new_n220), .A2(KEYINPUT69), .A3(new_n216), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n200), .A2(new_n203), .A3(new_n204), .ZN(new_n225));
  NOR2_X1   g039(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n227), .A2(G128), .A3(new_n228), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n225), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n202), .A2(G143), .ZN(new_n231));
  AND2_X1   g045(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n231), .B1(new_n232), .B2(new_n226), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(KEYINPUT68), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT68), .ZN(new_n235));
  OAI211_X1 g049(.A(new_n231), .B(new_n235), .C1(new_n232), .C2(new_n226), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n234), .A2(new_n236), .A3(G128), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n231), .A2(new_n204), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n230), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(new_n193), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n189), .A2(G137), .ZN(new_n241));
  OAI21_X1  g055(.A(G131), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(new_n197), .ZN(new_n243));
  OAI211_X1 g057(.A(new_n215), .B(new_n224), .C1(new_n239), .C2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT70), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n243), .ZN(new_n247));
  INV_X1    g061(.A(G128), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n248), .B1(new_n233), .B2(KEYINPUT68), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n210), .B1(new_n249), .B2(new_n236), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n247), .B1(new_n250), .B2(new_n230), .ZN(new_n251));
  NAND4_X1  g065(.A1(new_n251), .A2(KEYINPUT70), .A3(new_n224), .A4(new_n215), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n246), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  XNOR2_X1  g068(.A(KEYINPUT26), .B(G101), .ZN(new_n255));
  NOR2_X1   g069(.A1(G237), .A2(G953), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G210), .ZN(new_n257));
  XNOR2_X1  g071(.A(new_n255), .B(new_n257), .ZN(new_n258));
  XNOR2_X1  g072(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n259));
  XNOR2_X1  g073(.A(new_n258), .B(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT65), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n262), .B1(new_n207), .B2(new_n211), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n200), .A2(new_n203), .A3(new_n204), .A4(new_n206), .ZN(new_n264));
  OAI211_X1 g078(.A(new_n264), .B(KEYINPUT65), .C1(new_n210), .C2(new_n209), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n263), .A2(new_n198), .A3(new_n214), .A4(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(KEYINPUT30), .B1(new_n251), .B2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n224), .ZN(new_n269));
  OAI211_X1 g083(.A(new_n215), .B(KEYINPUT30), .C1(new_n239), .C2(new_n243), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n268), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  XNOR2_X1  g085(.A(KEYINPUT72), .B(KEYINPUT31), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n254), .A2(new_n261), .A3(new_n271), .A4(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n270), .ZN(new_n274));
  NOR3_X1   g088(.A1(new_n274), .A2(new_n267), .A3(new_n224), .ZN(new_n275));
  NOR3_X1   g089(.A1(new_n275), .A2(new_n253), .A3(new_n260), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT31), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n273), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n251), .A2(new_n266), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(new_n269), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n246), .A2(new_n280), .A3(new_n252), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(KEYINPUT28), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT28), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n244), .A2(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n261), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n187), .B1(new_n278), .B2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT32), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(KEYINPUT73), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n260), .B1(new_n275), .B2(new_n253), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT29), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n284), .A2(new_n261), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n293), .B1(new_n281), .B2(KEYINPUT28), .ZN(new_n294));
  OAI21_X1  g108(.A(KEYINPUT74), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(G902), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n293), .A2(new_n291), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n251), .A2(new_n215), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(new_n269), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n246), .A2(new_n299), .A3(new_n252), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT75), .ZN(new_n301));
  AND3_X1   g115(.A1(new_n300), .A2(new_n301), .A3(KEYINPUT28), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n301), .B1(new_n300), .B2(KEYINPUT28), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n297), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(new_n294), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT74), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n305), .A2(new_n306), .A3(new_n291), .A4(new_n290), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n295), .A2(new_n296), .A3(new_n304), .A4(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(G472), .ZN(new_n309));
  OR2_X1    g123(.A1(new_n286), .A2(new_n287), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT73), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n286), .A2(new_n311), .A3(new_n287), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n289), .A2(new_n309), .A3(new_n310), .A4(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G140), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G125), .ZN(new_n315));
  INV_X1    g129(.A(G125), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G140), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n315), .A2(new_n317), .A3(KEYINPUT77), .ZN(new_n318));
  OR3_X1    g132(.A1(new_n314), .A2(KEYINPUT77), .A3(G125), .ZN(new_n319));
  AND3_X1   g133(.A1(new_n318), .A2(G146), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(KEYINPUT18), .A2(G131), .ZN(new_n321));
  INV_X1    g135(.A(G237), .ZN(new_n322));
  INV_X1    g136(.A(G953), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n322), .A2(new_n323), .A3(G214), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n324), .A2(new_n199), .ZN(new_n325));
  AOI21_X1  g139(.A(G143), .B1(new_n256), .B2(G214), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n321), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n324), .A2(new_n199), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n256), .A2(G143), .A3(G214), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n328), .A2(KEYINPUT18), .A3(G131), .A4(new_n329), .ZN(new_n330));
  AOI22_X1  g144(.A1(KEYINPUT87), .A2(new_n320), .B1(new_n327), .B2(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n318), .A2(new_n319), .A3(G146), .ZN(new_n332));
  AND2_X1   g146(.A1(new_n315), .A2(new_n317), .ZN(new_n333));
  AOI21_X1  g147(.A(KEYINPUT87), .B1(new_n333), .B2(new_n202), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  AND2_X1   g149(.A1(new_n331), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n328), .A2(new_n329), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(G131), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n328), .A2(new_n196), .A3(new_n329), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n340), .A2(KEYINPUT17), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n318), .A2(new_n319), .A3(KEYINPUT16), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT16), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n315), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(G146), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n342), .A2(new_n202), .A3(new_n344), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n337), .A2(KEYINPUT17), .A3(G131), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n341), .B1(new_n349), .B2(KEYINPUT89), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT89), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n346), .A2(new_n351), .A3(new_n347), .A4(new_n348), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n336), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  XNOR2_X1  g167(.A(G113), .B(G122), .ZN(new_n354));
  INV_X1    g168(.A(G104), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n354), .B(new_n355), .ZN(new_n356));
  AOI22_X1  g170(.A1(new_n345), .A2(G146), .B1(new_n338), .B2(new_n339), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT19), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n358), .B1(new_n318), .B2(new_n319), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n333), .A2(KEYINPUT19), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n202), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  AOI22_X1  g175(.A1(new_n357), .A2(new_n361), .B1(new_n331), .B2(new_n335), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT88), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n356), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n331), .A2(new_n335), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n346), .A2(new_n361), .A3(new_n340), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(KEYINPUT88), .ZN(new_n368));
  AOI22_X1  g182(.A1(new_n353), .A2(new_n356), .B1(new_n364), .B2(new_n368), .ZN(new_n369));
  NOR2_X1   g183(.A1(G475), .A2(G902), .ZN(new_n370));
  XOR2_X1   g184(.A(new_n370), .B(KEYINPUT90), .Z(new_n371));
  OAI21_X1  g185(.A(KEYINPUT20), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n350), .A2(new_n352), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n373), .A2(new_n356), .A3(new_n365), .ZN(new_n374));
  INV_X1    g188(.A(new_n356), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n365), .A2(new_n366), .A3(new_n363), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n368), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT20), .ZN(new_n379));
  INV_X1    g193(.A(new_n371), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n356), .B1(new_n373), .B2(new_n365), .ZN(new_n382));
  AOI211_X1 g196(.A(new_n375), .B(new_n336), .C1(new_n350), .C2(new_n352), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n296), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  AOI22_X1  g198(.A1(new_n372), .A2(new_n381), .B1(G475), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n199), .A2(G128), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n248), .A2(G143), .ZN(new_n387));
  AND2_X1   g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  XNOR2_X1  g202(.A(new_n388), .B(new_n189), .ZN(new_n389));
  INV_X1    g203(.A(G116), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n390), .A2(KEYINPUT14), .A3(G122), .ZN(new_n391));
  XNOR2_X1  g205(.A(G116), .B(G122), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  OAI211_X1 g207(.A(G107), .B(new_n391), .C1(new_n393), .C2(KEYINPUT14), .ZN(new_n394));
  OAI211_X1 g208(.A(new_n389), .B(new_n394), .C1(G107), .C2(new_n393), .ZN(new_n395));
  INV_X1    g209(.A(new_n386), .ZN(new_n396));
  AND2_X1   g210(.A1(new_n396), .A2(KEYINPUT13), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n387), .B1(new_n396), .B2(KEYINPUT13), .ZN(new_n398));
  OAI21_X1  g212(.A(G134), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n388), .A2(new_n189), .ZN(new_n400));
  INV_X1    g214(.A(G107), .ZN(new_n401));
  XNOR2_X1  g215(.A(new_n392), .B(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n399), .A2(new_n400), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n395), .A2(new_n403), .ZN(new_n404));
  XNOR2_X1  g218(.A(KEYINPUT9), .B(G234), .ZN(new_n405));
  INV_X1    g219(.A(G217), .ZN(new_n406));
  NOR3_X1   g220(.A1(new_n405), .A2(new_n406), .A3(G953), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n404), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n395), .A2(new_n403), .A3(new_n407), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(G478), .ZN(new_n412));
  OR2_X1    g226(.A1(new_n412), .A2(KEYINPUT15), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n411), .A2(new_n296), .A3(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n413), .B1(new_n411), .B2(new_n296), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(G234), .A2(G237), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n418), .A2(G952), .A3(new_n323), .ZN(new_n419));
  XNOR2_X1  g233(.A(KEYINPUT21), .B(G898), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n418), .A2(G902), .A3(G953), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n419), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  AND2_X1   g237(.A1(new_n417), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n385), .A2(new_n424), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n425), .B(KEYINPUT91), .ZN(new_n426));
  OAI21_X1  g240(.A(G221), .B1(new_n405), .B2(G902), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  XNOR2_X1  g242(.A(G110), .B(G140), .ZN(new_n429));
  AND2_X1   g243(.A1(new_n323), .A2(G227), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n429), .B(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(G101), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n355), .A2(G107), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n401), .A2(G104), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n433), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT83), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n437), .A2(new_n401), .A3(KEYINPUT3), .A4(G104), .ZN(new_n438));
  NOR3_X1   g252(.A1(new_n355), .A2(KEYINPUT83), .A3(G107), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT3), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n440), .B1(new_n401), .B2(G104), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n438), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n436), .B1(new_n442), .B2(new_n433), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n239), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n231), .A2(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(G128), .ZN(new_n447));
  AND2_X1   g261(.A1(new_n447), .A2(new_n225), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n443), .B1(new_n448), .B2(new_n230), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n445), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n198), .A2(new_n214), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  OAI211_X1 g267(.A(KEYINPUT10), .B(new_n443), .C1(new_n250), .C2(new_n230), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT10), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n449), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n442), .A2(new_n433), .ZN(new_n457));
  OAI211_X1 g271(.A(G101), .B(new_n438), .C1(new_n439), .C2(new_n441), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n457), .A2(KEYINPUT4), .A3(new_n458), .ZN(new_n459));
  OR2_X1    g273(.A1(new_n439), .A2(new_n441), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT4), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n460), .A2(new_n461), .A3(G101), .A4(new_n438), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n459), .A2(new_n212), .A3(new_n462), .ZN(new_n463));
  AND3_X1   g277(.A1(new_n454), .A2(new_n456), .A3(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT84), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n451), .B(new_n465), .ZN(new_n466));
  AOI22_X1  g280(.A1(KEYINPUT12), .A2(new_n453), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT12), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n450), .A2(new_n468), .A3(new_n452), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n432), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n464), .A2(new_n451), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n451), .B(KEYINPUT84), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n454), .A2(new_n456), .A3(new_n463), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NOR3_X1   g288(.A1(new_n471), .A2(new_n474), .A3(new_n431), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n470), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(G469), .B1(new_n476), .B2(G902), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n431), .B1(new_n471), .B2(new_n474), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n453), .A2(KEYINPUT12), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n464), .A2(new_n466), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n479), .A2(new_n480), .A3(new_n469), .A4(new_n432), .ZN(new_n481));
  AOI21_X1  g295(.A(G902), .B1(new_n478), .B2(new_n481), .ZN(new_n482));
  XOR2_X1   g296(.A(KEYINPUT85), .B(G469), .Z(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n428), .B1(new_n477), .B2(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(G214), .B1(G237), .B2(G902), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n239), .A2(new_n316), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n212), .A2(new_n316), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(G224), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n492), .A2(G953), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n491), .B(new_n493), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n459), .A2(new_n223), .A3(new_n222), .A4(new_n462), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n216), .A2(KEYINPUT5), .ZN(new_n496));
  NOR3_X1   g310(.A1(new_n390), .A2(KEYINPUT5), .A3(G119), .ZN(new_n497));
  INV_X1    g311(.A(G113), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI22_X1  g313(.A1(new_n496), .A2(new_n499), .B1(new_n220), .B2(new_n216), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n443), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n495), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(KEYINPUT86), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT86), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n495), .A2(new_n504), .A3(new_n501), .ZN(new_n505));
  XNOR2_X1  g319(.A(G110), .B(G122), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n503), .A2(KEYINPUT6), .A3(new_n505), .A4(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n495), .A2(new_n501), .A3(new_n506), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n506), .B1(new_n502), .B2(KEYINPUT86), .ZN(new_n511));
  AOI21_X1  g325(.A(KEYINPUT6), .B1(new_n511), .B2(new_n505), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n494), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n491), .A2(new_n493), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n506), .B(KEYINPUT8), .ZN(new_n515));
  INV_X1    g329(.A(new_n501), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n443), .A2(new_n500), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT7), .ZN(new_n519));
  NOR3_X1   g333(.A1(new_n250), .A2(G125), .A3(new_n230), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n519), .B1(new_n520), .B2(new_n489), .ZN(new_n521));
  AND4_X1   g335(.A1(new_n514), .A2(new_n509), .A3(new_n518), .A4(new_n521), .ZN(new_n522));
  OR3_X1    g336(.A1(new_n491), .A2(new_n519), .A3(new_n493), .ZN(new_n523));
  AOI21_X1  g337(.A(G902), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n513), .A2(new_n524), .ZN(new_n525));
  OAI21_X1  g339(.A(G210), .B1(G237), .B2(G902), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n513), .A2(new_n524), .A3(new_n526), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n487), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  AND2_X1   g344(.A1(new_n485), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT80), .ZN(new_n532));
  XNOR2_X1  g346(.A(KEYINPUT22), .B(G137), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n323), .A2(G221), .A3(G234), .ZN(new_n534));
  XOR2_X1   g348(.A(new_n533), .B(new_n534), .Z(new_n535));
  XNOR2_X1  g349(.A(new_n535), .B(KEYINPUT79), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n248), .A2(G119), .ZN(new_n538));
  INV_X1    g352(.A(G119), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(G128), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  XNOR2_X1  g355(.A(KEYINPUT24), .B(G110), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT23), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n544), .B1(new_n539), .B2(G128), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n248), .A2(KEYINPUT23), .A3(G119), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n545), .A2(new_n546), .A3(new_n540), .ZN(new_n547));
  OR2_X1    g361(.A1(new_n547), .A2(KEYINPUT76), .ZN(new_n548));
  INV_X1    g362(.A(G110), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n549), .B1(new_n547), .B2(KEYINPUT76), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n543), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(new_n347), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n202), .B1(new_n342), .B2(new_n344), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n551), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT78), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n551), .B(KEYINPUT78), .C1(new_n552), .C2(new_n553), .ZN(new_n557));
  AND2_X1   g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  OR2_X1    g372(.A1(new_n547), .A2(G110), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n541), .A2(new_n542), .ZN(new_n560));
  AOI22_X1  g374(.A1(new_n559), .A2(new_n560), .B1(new_n202), .B2(new_n333), .ZN(new_n561));
  AND2_X1   g375(.A1(new_n561), .A2(new_n346), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n532), .B(new_n537), .C1(new_n558), .C2(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n562), .B1(new_n556), .B2(new_n557), .ZN(new_n564));
  OAI21_X1  g378(.A(KEYINPUT80), .B1(new_n564), .B2(new_n536), .ZN(new_n565));
  INV_X1    g379(.A(new_n535), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n563), .A2(new_n565), .A3(new_n296), .A4(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT25), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AOI211_X1 g384(.A(new_n535), .B(new_n562), .C1(new_n556), .C2(new_n557), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n564), .A2(new_n536), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n571), .B1(new_n572), .B2(new_n532), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n573), .A2(KEYINPUT25), .A3(new_n296), .A4(new_n565), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n406), .B1(G234), .B2(new_n296), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n576), .A2(G902), .ZN(new_n578));
  XOR2_X1   g392(.A(new_n578), .B(KEYINPUT81), .Z(new_n579));
  NAND4_X1  g393(.A1(new_n563), .A2(new_n565), .A3(new_n567), .A4(new_n579), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n580), .B(KEYINPUT82), .ZN(new_n581));
  AND2_X1   g395(.A1(new_n577), .A2(new_n581), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n313), .A2(new_n426), .A3(new_n531), .A4(new_n582), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n583), .B(G101), .ZN(G3));
  INV_X1    g398(.A(G469), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n479), .A2(new_n480), .A3(new_n469), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(new_n431), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n480), .B(new_n432), .C1(new_n451), .C2(new_n464), .ZN(new_n588));
  AOI21_X1  g402(.A(G902), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n484), .B1(new_n585), .B2(new_n589), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n577), .A2(new_n581), .A3(new_n427), .A4(new_n590), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n278), .A2(new_n285), .ZN(new_n592));
  OAI21_X1  g406(.A(G472), .B1(new_n592), .B2(G902), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n286), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  AND3_X1   g409(.A1(new_n513), .A2(new_n524), .A3(new_n526), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n526), .B1(new_n513), .B2(new_n524), .ZN(new_n597));
  OAI211_X1 g411(.A(new_n423), .B(new_n486), .C1(new_n596), .C2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n384), .A2(G475), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n379), .B1(new_n378), .B2(new_n380), .ZN(new_n600));
  AOI211_X1 g414(.A(KEYINPUT20), .B(new_n371), .C1(new_n374), .C2(new_n377), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n599), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n412), .A2(new_n296), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n411), .A2(new_n296), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n604), .B1(new_n605), .B2(G478), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n411), .B(KEYINPUT33), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n606), .B1(new_n608), .B2(G478), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n602), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(KEYINPUT92), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT92), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n602), .A2(new_n609), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n598), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n595), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(KEYINPUT93), .ZN(new_n616));
  XOR2_X1   g430(.A(KEYINPUT34), .B(G104), .Z(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G6));
  AOI21_X1  g432(.A(new_n417), .B1(G475), .B2(new_n384), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n601), .A2(KEYINPUT94), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT94), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n372), .A2(new_n621), .A3(new_n381), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n619), .A2(new_n423), .A3(new_n620), .A4(new_n622), .ZN(new_n623));
  OR2_X1    g437(.A1(new_n623), .A2(KEYINPUT95), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(KEYINPUT95), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n624), .A2(new_n530), .A3(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(new_n595), .ZN(new_n628));
  XOR2_X1   g442(.A(KEYINPUT35), .B(G107), .Z(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G9));
  INV_X1    g444(.A(new_n594), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n564), .B(KEYINPUT96), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n537), .A2(KEYINPUT36), .ZN(new_n633));
  XOR2_X1   g447(.A(new_n632), .B(new_n633), .Z(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n579), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(new_n577), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n426), .A2(new_n531), .A3(new_n631), .A4(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(KEYINPUT37), .B(G110), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(KEYINPUT97), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n637), .B(new_n639), .ZN(G12));
  AND2_X1   g454(.A1(new_n531), .A2(new_n636), .ZN(new_n641));
  AND2_X1   g455(.A1(new_n622), .A2(new_n620), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n419), .B(KEYINPUT99), .ZN(new_n643));
  XNOR2_X1  g457(.A(KEYINPUT98), .B(G900), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n643), .B1(new_n422), .B2(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(KEYINPUT100), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  AND3_X1   g461(.A1(new_n642), .A2(new_n619), .A3(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n641), .A2(new_n313), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(KEYINPUT101), .B(G128), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G30));
  XOR2_X1   g465(.A(KEYINPUT103), .B(KEYINPUT39), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n646), .B(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n485), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g468(.A(new_n654), .B(KEYINPUT40), .Z(new_n655));
  INV_X1    g469(.A(new_n310), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n254), .A2(new_n271), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n261), .ZN(new_n658));
  OAI211_X1 g472(.A(new_n658), .B(new_n296), .C1(new_n261), .C2(new_n300), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n656), .B1(G472), .B2(new_n659), .ZN(new_n660));
  AND2_X1   g474(.A1(new_n289), .A2(new_n312), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n528), .A2(new_n529), .ZN(new_n663));
  XNOR2_X1  g477(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n417), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n602), .A2(new_n666), .ZN(new_n667));
  NOR4_X1   g481(.A1(new_n665), .A2(new_n487), .A3(new_n636), .A4(new_n667), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n655), .A2(new_n662), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G143), .ZN(G45));
  NOR2_X1   g484(.A1(new_n610), .A2(new_n646), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n641), .A2(new_n313), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G146), .ZN(G48));
  NOR2_X1   g487(.A1(new_n482), .A2(new_n585), .ZN(new_n674));
  INV_X1    g488(.A(new_n483), .ZN(new_n675));
  AOI211_X1 g489(.A(G902), .B(new_n675), .C1(new_n478), .C2(new_n481), .ZN(new_n676));
  NOR3_X1   g490(.A1(new_n674), .A2(new_n676), .A3(new_n428), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n313), .A2(new_n614), .A3(new_n582), .A4(new_n677), .ZN(new_n678));
  XOR2_X1   g492(.A(KEYINPUT41), .B(G113), .Z(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(KEYINPUT104), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n678), .B(new_n680), .ZN(G15));
  NAND4_X1  g495(.A1(new_n627), .A2(new_n313), .A3(new_n582), .A4(new_n677), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G116), .ZN(G18));
  INV_X1    g497(.A(KEYINPUT105), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n486), .B1(new_n596), .B2(new_n597), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n478), .A2(new_n481), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(new_n296), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(G469), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n688), .A2(new_n427), .A3(new_n484), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n684), .B1(new_n685), .B2(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n530), .A2(new_n677), .A3(KEYINPUT105), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n692), .A2(new_n313), .A3(new_n426), .A4(new_n636), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G119), .ZN(G21));
  OAI21_X1  g508(.A(new_n284), .B1(new_n302), .B2(new_n303), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n261), .B1(new_n695), .B2(KEYINPUT106), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT106), .ZN(new_n697));
  OAI211_X1 g511(.A(new_n697), .B(new_n284), .C1(new_n302), .C2(new_n303), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n278), .B1(new_n696), .B2(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(new_n187), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n593), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n688), .A2(new_n423), .A3(new_n427), .A4(new_n484), .ZN(new_n703));
  NOR3_X1   g517(.A1(new_n703), .A2(new_n685), .A3(new_n667), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n702), .A2(new_n582), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G122), .ZN(G24));
  INV_X1    g520(.A(new_n636), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n707), .A2(new_n701), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n708), .A2(new_n671), .A3(new_n692), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G125), .ZN(G27));
  NAND3_X1  g524(.A1(new_n309), .A2(new_n310), .A3(new_n288), .ZN(new_n711));
  AND2_X1   g525(.A1(new_n711), .A2(new_n582), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n528), .A2(new_n486), .A3(new_n529), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT108), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n528), .A2(KEYINPUT108), .A3(new_n486), .A4(new_n529), .ZN(new_n716));
  OAI21_X1  g530(.A(KEYINPUT107), .B1(new_n470), .B2(new_n475), .ZN(new_n717));
  OR2_X1    g531(.A1(new_n475), .A2(KEYINPUT107), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n717), .A2(new_n718), .A3(G469), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n585), .A2(new_n296), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n720), .B1(new_n482), .B2(new_n483), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n428), .B1(new_n719), .B2(new_n721), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n715), .A2(new_n671), .A3(new_n716), .A4(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n712), .A2(KEYINPUT42), .A3(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  AND3_X1   g540(.A1(new_n715), .A2(new_n716), .A3(new_n722), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n727), .A2(new_n313), .A3(new_n582), .A4(new_n671), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT42), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT109), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n728), .A2(KEYINPUT109), .A3(new_n729), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n726), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(new_n196), .ZN(G33));
  NAND4_X1  g549(.A1(new_n727), .A2(new_n648), .A3(new_n313), .A4(new_n582), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G134), .ZN(G36));
  INV_X1    g551(.A(new_n606), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n738), .B1(new_n607), .B2(new_n412), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n602), .A2(new_n739), .ZN(new_n740));
  XOR2_X1   g554(.A(new_n740), .B(KEYINPUT43), .Z(new_n741));
  NOR3_X1   g555(.A1(new_n741), .A2(new_n631), .A3(new_n707), .ZN(new_n742));
  OR2_X1    g556(.A1(new_n742), .A2(KEYINPUT44), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n715), .A2(new_n716), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n744), .B1(new_n742), .B2(KEYINPUT44), .ZN(new_n745));
  AND2_X1   g559(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  AND3_X1   g560(.A1(new_n717), .A2(KEYINPUT45), .A3(new_n718), .ZN(new_n747));
  OAI21_X1  g561(.A(G469), .B1(new_n476), .B2(KEYINPUT45), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n749), .A2(new_n720), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n484), .B1(new_n750), .B2(KEYINPUT46), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(KEYINPUT46), .ZN(new_n752));
  OR2_X1    g566(.A1(new_n752), .A2(KEYINPUT110), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(KEYINPUT110), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n751), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n755), .A2(new_n428), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n746), .A2(new_n653), .A3(new_n756), .ZN(new_n757));
  XOR2_X1   g571(.A(KEYINPUT111), .B(G137), .Z(new_n758));
  XNOR2_X1  g572(.A(new_n757), .B(new_n758), .ZN(G39));
  INV_X1    g573(.A(new_n671), .ZN(new_n760));
  NOR4_X1   g574(.A1(new_n313), .A2(new_n744), .A3(new_n760), .A4(new_n582), .ZN(new_n761));
  INV_X1    g575(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n756), .A2(KEYINPUT47), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT47), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n764), .B1(new_n755), .B2(new_n428), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n762), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(new_n314), .ZN(G42));
  NOR2_X1   g581(.A1(new_n741), .A2(new_n643), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n768), .A2(new_n582), .A3(new_n702), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n689), .A2(new_n486), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n769), .A2(new_n665), .A3(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT50), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n771), .B(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(new_n662), .ZN(new_n774));
  INV_X1    g588(.A(new_n419), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n744), .A2(new_n689), .ZN(new_n776));
  AND4_X1   g590(.A1(new_n582), .A2(new_n774), .A3(new_n775), .A4(new_n776), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n602), .A2(new_n609), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n768), .A2(new_n776), .ZN(new_n779));
  AOI22_X1  g593(.A1(new_n777), .A2(new_n778), .B1(new_n708), .B2(new_n779), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n773), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(KEYINPUT51), .ZN(new_n782));
  INV_X1    g596(.A(new_n769), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n783), .A2(new_n744), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n674), .A2(new_n676), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n428), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n763), .A2(new_n765), .A3(new_n786), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n782), .B1(new_n784), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n763), .A2(new_n765), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n786), .B(KEYINPUT118), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n784), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  AOI21_X1  g605(.A(KEYINPUT51), .B1(new_n781), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n779), .A2(new_n712), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(KEYINPUT48), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n769), .A2(new_n692), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n323), .A2(G952), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n611), .A2(new_n613), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n796), .B1(new_n777), .B2(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n794), .A2(new_n795), .A3(new_n798), .ZN(new_n799));
  OR3_X1    g613(.A1(new_n788), .A2(new_n792), .A3(new_n799), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n649), .A2(new_n672), .A3(new_n709), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT52), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n685), .A2(new_n667), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n636), .A2(new_n646), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n662), .A2(new_n803), .A3(new_n722), .A4(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n801), .A2(new_n802), .A3(new_n805), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n805), .A2(new_n649), .A3(new_n672), .A4(new_n709), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(KEYINPUT52), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n313), .A2(new_n582), .A3(new_n677), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n678), .B1(new_n810), .B2(new_n626), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT114), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT113), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n813), .B1(new_n385), .B2(new_n739), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n602), .A2(new_n609), .A3(KEYINPUT113), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n812), .B1(new_n816), .B2(new_n598), .ZN(new_n817));
  INV_X1    g631(.A(new_n598), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n818), .A2(KEYINPUT114), .A3(new_n814), .A4(new_n815), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n595), .A2(new_n817), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(new_n705), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n811), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n602), .A2(new_n417), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n595), .A2(new_n818), .A3(new_n823), .ZN(new_n824));
  AND4_X1   g638(.A1(new_n583), .A2(new_n693), .A3(new_n637), .A4(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT115), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n702), .A2(new_n636), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n826), .B1(new_n827), .B2(new_n723), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n708), .A2(new_n724), .A3(KEYINPUT115), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n666), .A2(new_n646), .ZN(new_n831));
  AND4_X1   g645(.A1(new_n599), .A2(new_n485), .A3(new_n642), .A4(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(new_n744), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n832), .A2(new_n833), .A3(new_n313), .A4(new_n636), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n834), .A2(new_n736), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n822), .A2(new_n825), .A3(new_n830), .A4(new_n835), .ZN(new_n836));
  OAI21_X1  g650(.A(KEYINPUT116), .B1(new_n836), .B2(new_n734), .ZN(new_n837));
  INV_X1    g651(.A(new_n733), .ZN(new_n838));
  AOI21_X1  g652(.A(KEYINPUT109), .B1(new_n728), .B2(new_n729), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n725), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n693), .A2(new_n824), .A3(new_n583), .A4(new_n637), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n841), .A2(new_n811), .A3(new_n821), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n834), .A2(new_n736), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n843), .B1(new_n828), .B2(new_n829), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT116), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n840), .A2(new_n842), .A3(new_n844), .A4(new_n845), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n809), .B1(new_n837), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n649), .A2(new_n709), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(KEYINPUT52), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT53), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n847), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n837), .A2(new_n846), .ZN(new_n853));
  INV_X1    g667(.A(new_n809), .ZN(new_n854));
  AOI21_X1  g668(.A(KEYINPUT53), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g669(.A(KEYINPUT54), .B1(new_n852), .B2(new_n855), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n836), .A2(new_n734), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n850), .B1(new_n848), .B2(KEYINPUT52), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n854), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  XNOR2_X1  g673(.A(KEYINPUT117), .B(KEYINPUT54), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n859), .B(new_n860), .C1(new_n847), .C2(KEYINPUT53), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n856), .A2(new_n861), .ZN(new_n862));
  OAI22_X1  g676(.A1(new_n800), .A2(new_n862), .B1(G952), .B2(G953), .ZN(new_n863));
  XNOR2_X1  g677(.A(new_n785), .B(KEYINPUT49), .ZN(new_n864));
  AND4_X1   g678(.A1(new_n427), .A2(new_n864), .A3(new_n486), .A4(new_n740), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n774), .A2(new_n865), .A3(new_n582), .A4(new_n665), .ZN(new_n866));
  XOR2_X1   g680(.A(new_n866), .B(KEYINPUT112), .Z(new_n867));
  NAND2_X1  g681(.A1(new_n863), .A2(new_n867), .ZN(G75));
  NOR2_X1   g682(.A1(new_n323), .A2(G952), .ZN(new_n869));
  AND4_X1   g683(.A1(new_n806), .A2(new_n857), .A3(new_n808), .A4(new_n858), .ZN(new_n870));
  OAI211_X1 g684(.A(G210), .B(G902), .C1(new_n855), .C2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT56), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n510), .A2(new_n512), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n874), .B(new_n494), .ZN(new_n875));
  XNOR2_X1  g689(.A(KEYINPUT119), .B(KEYINPUT55), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n875), .B(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n869), .B1(new_n873), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n871), .A2(KEYINPUT120), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n859), .B1(new_n847), .B2(KEYINPUT53), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT120), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n880), .A2(new_n881), .A3(G210), .A4(G902), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n877), .A2(KEYINPUT56), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n879), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n878), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(KEYINPUT121), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT121), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n878), .A2(new_n887), .A3(new_n884), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n886), .A2(new_n888), .ZN(G51));
  XNOR2_X1  g703(.A(new_n720), .B(KEYINPUT57), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n853), .A2(new_n854), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(new_n850), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n860), .B1(new_n892), .B2(new_n859), .ZN(new_n893));
  INV_X1    g707(.A(new_n861), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n890), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(new_n686), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n296), .B1(new_n892), .B2(new_n859), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(new_n749), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n869), .B1(new_n896), .B2(new_n898), .ZN(G54));
  AND2_X1   g713(.A1(KEYINPUT58), .A2(G475), .ZN(new_n900));
  AND3_X1   g714(.A1(new_n897), .A2(new_n378), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n378), .B1(new_n897), .B2(new_n900), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n901), .A2(new_n902), .A3(new_n869), .ZN(G60));
  INV_X1    g717(.A(new_n869), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n603), .B(KEYINPUT59), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n905), .B1(new_n856), .B2(new_n861), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n904), .B1(new_n906), .B2(new_n607), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n608), .A2(new_n905), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n908), .B1(new_n893), .B2(new_n894), .ZN(new_n909));
  OR2_X1    g723(.A1(new_n909), .A2(KEYINPUT122), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(KEYINPUT122), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n907), .B1(new_n910), .B2(new_n911), .ZN(G63));
  NAND2_X1  g726(.A1(G217), .A2(G902), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(KEYINPUT60), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n914), .B1(new_n892), .B2(new_n859), .ZN(new_n915));
  AND2_X1   g729(.A1(new_n573), .A2(new_n565), .ZN(new_n916));
  OR2_X1    g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n915), .A2(new_n634), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n917), .A2(new_n904), .A3(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT61), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n917), .A2(KEYINPUT61), .A3(new_n904), .A4(new_n918), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(G66));
  OAI21_X1  g737(.A(G953), .B1(new_n420), .B2(new_n492), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n924), .B1(new_n842), .B2(G953), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n874), .B1(G898), .B2(new_n323), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n925), .B(new_n926), .ZN(G69));
  AOI21_X1  g741(.A(new_n323), .B1(G227), .B2(G900), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n268), .A2(new_n270), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n359), .A2(new_n360), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n930), .B(new_n931), .Z(new_n932));
  AOI21_X1  g746(.A(new_n932), .B1(G900), .B2(G953), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n756), .A2(new_n653), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n712), .A2(new_n803), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n736), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n936), .A2(new_n766), .ZN(new_n937));
  AOI21_X1  g751(.A(KEYINPUT124), .B1(new_n757), .B2(new_n801), .ZN(new_n938));
  AND3_X1   g752(.A1(new_n757), .A2(KEYINPUT124), .A3(new_n801), .ZN(new_n939));
  OAI211_X1 g753(.A(new_n937), .B(new_n840), .C1(new_n938), .C2(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n933), .B1(new_n940), .B2(G953), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n313), .A2(new_n582), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n823), .B1(new_n814), .B2(new_n815), .ZN(new_n943));
  OR4_X1    g757(.A1(new_n942), .A2(new_n654), .A3(new_n744), .A4(new_n943), .ZN(new_n944));
  AND2_X1   g758(.A1(new_n757), .A2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n766), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n801), .A2(new_n669), .ZN(new_n947));
  OR2_X1    g761(.A1(new_n947), .A2(KEYINPUT62), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(KEYINPUT62), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n945), .A2(new_n946), .A3(new_n948), .A4(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n323), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n932), .B(KEYINPUT123), .Z(new_n952));
  NAND2_X1  g766(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT125), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n941), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n954), .B1(new_n941), .B2(new_n953), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n929), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n941), .A2(new_n953), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(KEYINPUT125), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n960), .A2(new_n928), .A3(new_n955), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n958), .A2(new_n961), .ZN(G72));
  NAND2_X1  g776(.A1(G472), .A2(G902), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT63), .Z(new_n964));
  INV_X1    g778(.A(new_n842), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n964), .B1(new_n940), .B2(new_n965), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n657), .A2(new_n261), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n869), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n964), .B1(new_n950), .B2(new_n965), .ZN(new_n969));
  AND2_X1   g783(.A1(new_n969), .A2(KEYINPUT126), .ZN(new_n970));
  OAI211_X1 g784(.A(new_n261), .B(new_n657), .C1(new_n969), .C2(KEYINPUT126), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n968), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n658), .A2(new_n964), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n973), .A2(new_n967), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n974), .B1(new_n852), .B2(new_n855), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT127), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  OR2_X1    g791(.A1(new_n975), .A2(new_n976), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n972), .B1(new_n977), .B2(new_n978), .ZN(G57));
endmodule


