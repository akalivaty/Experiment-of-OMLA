//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 0 0 1 0 1 0 0 0 1 0 1 0 0 1 1 1 1 1 1 0 1 1 0 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 1 0 1 1 1 0 0 0 1 1 1 0 1 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:58 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1252, new_n1253, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NOR3_X1   g0007(.A1(new_n207), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0008(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  INV_X1    g0010(.A(G87), .ZN(new_n211));
  INV_X1    g0011(.A(G250), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(G50), .ZN(new_n214));
  INV_X1    g0014(.A(G226), .ZN(new_n215));
  INV_X1    g0015(.A(G116), .ZN(new_n216));
  INV_X1    g0016(.A(G270), .ZN(new_n217));
  OAI22_X1  g0017(.A1(new_n214), .A2(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  AOI211_X1 g0018(.A(new_n213), .B(new_n218), .C1(G97), .C2(G257), .ZN(new_n219));
  INV_X1    g0019(.A(G238), .ZN(new_n220));
  INV_X1    g0020(.A(G244), .ZN(new_n221));
  XNOR2_X1  g0021(.A(KEYINPUT65), .B(G77), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n202), .B2(new_n220), .C1(new_n221), .C2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT66), .Z(new_n226));
  OAI21_X1  g0026(.A(new_n210), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  OR2_X1    g0027(.A1(new_n227), .A2(KEYINPUT1), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT67), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n210), .A2(G13), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n230), .B(G250), .C1(G257), .C2(G264), .ZN(new_n231));
  INV_X1    g0031(.A(KEYINPUT0), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n206), .A2(new_n214), .ZN(new_n234));
  NAND2_X1  g0034(.A1(G1), .A2(G13), .ZN(new_n235));
  INV_X1    g0035(.A(new_n235), .ZN(new_n236));
  NAND3_X1  g0036(.A1(new_n234), .A2(G20), .A3(new_n236), .ZN(new_n237));
  OAI21_X1  g0037(.A(new_n237), .B1(new_n232), .B2(new_n231), .ZN(new_n238));
  AOI21_X1  g0038(.A(new_n238), .B1(new_n227), .B2(KEYINPUT1), .ZN(new_n239));
  NAND3_X1  g0039(.A1(new_n229), .A2(new_n233), .A3(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT68), .ZN(G361));
  XNOR2_X1  g0041(.A(G238), .B(G244), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G232), .ZN(new_n243));
  XNOR2_X1  g0043(.A(KEYINPUT2), .B(G226), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G250), .B(G257), .Z(new_n246));
  XNOR2_X1  g0046(.A(G264), .B(G270), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G358));
  XOR2_X1   g0049(.A(G68), .B(G77), .Z(new_n250));
  XNOR2_X1  g0050(.A(G50), .B(G58), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(G87), .B(G97), .Z(new_n253));
  XNOR2_X1  g0053(.A(G107), .B(G116), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n252), .B(new_n255), .ZN(G351));
  NAND2_X1  g0056(.A1(KEYINPUT73), .A2(KEYINPUT9), .ZN(new_n257));
  OAI21_X1  g0057(.A(G20), .B1(new_n207), .B2(G50), .ZN(new_n258));
  INV_X1    g0058(.A(G150), .ZN(new_n259));
  NOR2_X1   g0059(.A1(G20), .A2(G33), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  XNOR2_X1  g0061(.A(KEYINPUT8), .B(G58), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT70), .ZN(new_n263));
  INV_X1    g0063(.A(G33), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n263), .B1(new_n264), .B2(G20), .ZN(new_n265));
  INV_X1    g0065(.A(G20), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n266), .A2(KEYINPUT70), .A3(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  OAI221_X1 g0068(.A(new_n258), .B1(new_n259), .B2(new_n261), .C1(new_n262), .C2(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(new_n235), .ZN(new_n271));
  INV_X1    g0071(.A(G13), .ZN(new_n272));
  NOR3_X1   g0072(.A1(new_n272), .A2(new_n266), .A3(G1), .ZN(new_n273));
  AOI22_X1  g0073(.A1(new_n269), .A2(new_n271), .B1(new_n214), .B2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n271), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n275), .B1(G1), .B2(new_n266), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G50), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n274), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT72), .ZN(new_n280));
  XNOR2_X1  g0080(.A(new_n279), .B(new_n280), .ZN(new_n281));
  NOR2_X1   g0081(.A1(KEYINPUT73), .A2(KEYINPUT9), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n257), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n264), .A2(KEYINPUT3), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT3), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  XNOR2_X1  g0087(.A(KEYINPUT69), .B(G1698), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n287), .B1(G222), .B2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G223), .ZN(new_n290));
  INV_X1    g0090(.A(G1698), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n289), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n235), .B1(G33), .B2(G41), .ZN(new_n293));
  XNOR2_X1  g0093(.A(KEYINPUT3), .B(G33), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n292), .B(new_n293), .C1(new_n222), .C2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G1), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n296), .B1(G41), .B2(G45), .ZN(new_n297));
  INV_X1    g0097(.A(G274), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n293), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(new_n297), .ZN(new_n302));
  OAI211_X1 g0102(.A(new_n295), .B(new_n300), .C1(new_n215), .C2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G190), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n305), .B1(G200), .B2(new_n303), .ZN(new_n306));
  XNOR2_X1  g0106(.A(new_n279), .B(KEYINPUT72), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n307), .A2(KEYINPUT73), .A3(KEYINPUT9), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n283), .A2(new_n306), .A3(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(KEYINPUT10), .B1(new_n306), .B2(KEYINPUT74), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n310), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n312), .A2(new_n283), .A3(new_n306), .A4(new_n308), .ZN(new_n313));
  OR2_X1    g0113(.A1(new_n303), .A2(G179), .ZN(new_n314));
  INV_X1    g0114(.A(G169), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n303), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n314), .A2(new_n279), .A3(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n311), .A2(new_n313), .A3(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT13), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n284), .A2(new_n286), .A3(G232), .A4(G1698), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT75), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n294), .A2(KEYINPUT75), .A3(G232), .A4(G1698), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(G33), .A2(G97), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n294), .A2(new_n288), .A3(G226), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(new_n293), .ZN(new_n328));
  INV_X1    g0128(.A(new_n302), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(G238), .ZN(new_n330));
  AND4_X1   g0130(.A1(new_n319), .A2(new_n328), .A3(new_n300), .A4(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n299), .B1(new_n327), .B2(new_n293), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n319), .B1(new_n332), .B2(new_n330), .ZN(new_n333));
  OAI21_X1  g0133(.A(G169), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(KEYINPUT14), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n331), .A2(new_n333), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(G179), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT14), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n338), .B(G169), .C1(new_n331), .C2(new_n333), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n335), .A2(new_n337), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n202), .A2(G20), .ZN(new_n341));
  INV_X1    g0141(.A(G77), .ZN(new_n342));
  OAI221_X1 g0142(.A(new_n341), .B1(new_n214), .B2(new_n261), .C1(new_n268), .C2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(new_n271), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  AOI22_X1  g0145(.A1(new_n345), .A2(KEYINPUT11), .B1(G68), .B2(new_n277), .ZN(new_n346));
  NOR3_X1   g0146(.A1(new_n341), .A2(G1), .A3(new_n272), .ZN(new_n347));
  XNOR2_X1  g0147(.A(new_n347), .B(KEYINPUT12), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n346), .B(new_n349), .C1(KEYINPUT11), .C2(new_n345), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n340), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n350), .B1(new_n336), .B2(G190), .ZN(new_n352));
  INV_X1    g0152(.A(G200), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n352), .B1(new_n353), .B2(new_n336), .ZN(new_n354));
  AND2_X1   g0154(.A1(KEYINPUT69), .A2(G1698), .ZN(new_n355));
  NOR2_X1   g0155(.A1(KEYINPUT69), .A2(G1698), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(G232), .ZN(new_n358));
  OAI221_X1 g0158(.A(new_n294), .B1(new_n220), .B2(new_n291), .C1(new_n357), .C2(new_n358), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n359), .B(new_n293), .C1(G107), .C2(new_n294), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n360), .B(new_n300), .C1(new_n221), .C2(new_n302), .ZN(new_n361));
  OR2_X1    g0161(.A1(new_n361), .A2(G179), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n222), .A2(G20), .ZN(new_n363));
  XNOR2_X1  g0163(.A(KEYINPUT15), .B(G87), .ZN(new_n364));
  OAI221_X1 g0164(.A(new_n363), .B1(new_n261), .B2(new_n262), .C1(new_n268), .C2(new_n364), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n365), .A2(new_n271), .B1(new_n223), .B2(new_n273), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n277), .A2(G77), .ZN(new_n367));
  AND2_X1   g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n361), .A2(new_n315), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n362), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n351), .A2(new_n354), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n361), .A2(G200), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(new_n368), .ZN(new_n374));
  XNOR2_X1  g0174(.A(new_n374), .B(KEYINPUT71), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n361), .A2(new_n304), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT76), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n378), .B1(new_n285), .B2(G33), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(new_n286), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n378), .A2(new_n285), .A3(G33), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n380), .A2(G226), .A3(G1698), .A4(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(KEYINPUT78), .ZN(new_n383));
  NOR3_X1   g0183(.A1(new_n264), .A2(KEYINPUT76), .A3(KEYINPUT3), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n384), .B1(new_n286), .B2(new_n379), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT78), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n385), .A2(new_n386), .A3(G226), .A4(G1698), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n385), .A2(G223), .A3(new_n288), .ZN(new_n388));
  NAND2_X1  g0188(.A1(G33), .A2(G87), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT79), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n383), .A2(new_n387), .A3(new_n388), .A4(new_n391), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n389), .A2(new_n390), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n293), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n329), .A2(G232), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n394), .A2(new_n300), .A3(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(G179), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(KEYINPUT76), .B1(new_n264), .B2(KEYINPUT3), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n264), .A2(KEYINPUT3), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n381), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n401), .A2(new_n357), .ZN(new_n402));
  AOI22_X1  g0202(.A1(G223), .A2(new_n402), .B1(new_n382), .B2(KEYINPUT78), .ZN(new_n403));
  INV_X1    g0203(.A(new_n393), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n403), .A2(new_n404), .A3(new_n387), .A4(new_n391), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n299), .B1(new_n405), .B2(new_n293), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n315), .B1(new_n406), .B2(new_n395), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n203), .B(new_n205), .C1(new_n201), .C2(new_n202), .ZN(new_n408));
  AOI22_X1  g0208(.A1(new_n408), .A2(G20), .B1(G159), .B2(new_n260), .ZN(new_n409));
  AOI21_X1  g0209(.A(G20), .B1(new_n380), .B2(new_n381), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT7), .ZN(new_n411));
  OAI21_X1  g0211(.A(G68), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NOR3_X1   g0212(.A1(new_n385), .A2(KEYINPUT7), .A3(G20), .ZN(new_n413));
  OAI211_X1 g0213(.A(KEYINPUT16), .B(new_n409), .C1(new_n412), .C2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT16), .ZN(new_n415));
  INV_X1    g0215(.A(new_n409), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n411), .B1(new_n294), .B2(G20), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n287), .A2(KEYINPUT7), .A3(new_n266), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n202), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n415), .B1(new_n416), .B2(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n414), .A2(new_n271), .A3(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT77), .ZN(new_n422));
  INV_X1    g0222(.A(new_n273), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(new_n262), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n424), .B1(new_n277), .B2(new_n262), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n421), .A2(new_n422), .A3(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n422), .B1(new_n421), .B2(new_n425), .ZN(new_n428));
  OAI22_X1  g0228(.A1(new_n398), .A2(new_n407), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(KEYINPUT18), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n396), .A2(G200), .ZN(new_n431));
  AND2_X1   g0231(.A1(new_n421), .A2(new_n425), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT80), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n394), .A2(G190), .A3(new_n300), .A4(new_n395), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n431), .A2(new_n432), .A3(new_n433), .A4(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT17), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n421), .A2(new_n425), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n438), .B1(G200), .B2(new_n396), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n439), .A2(new_n433), .A3(KEYINPUT17), .A4(new_n434), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n438), .A2(KEYINPUT77), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(new_n426), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n396), .A2(G169), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n406), .A2(G179), .A3(new_n395), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT18), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n442), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n430), .A2(new_n437), .A3(new_n440), .A4(new_n447), .ZN(new_n448));
  NOR4_X1   g0248(.A1(new_n318), .A2(new_n372), .A3(new_n377), .A4(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT87), .ZN(new_n451));
  OAI21_X1  g0251(.A(G250), .B1(new_n355), .B2(new_n356), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n451), .B1(new_n401), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(G33), .A2(G294), .ZN(new_n454));
  OR2_X1    g0254(.A1(KEYINPUT69), .A2(G1698), .ZN(new_n455));
  NAND2_X1  g0255(.A1(KEYINPUT69), .A2(G1698), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n212), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n457), .A2(new_n380), .A3(KEYINPUT87), .A4(new_n381), .ZN(new_n458));
  AND2_X1   g0258(.A1(G257), .A2(G1698), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n380), .A2(new_n381), .A3(new_n459), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n453), .A2(new_n454), .A3(new_n458), .A4(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(KEYINPUT88), .ZN(new_n462));
  AOI22_X1  g0262(.A1(new_n385), .A2(new_n459), .B1(G33), .B2(G294), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT88), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n463), .A2(new_n464), .A3(new_n453), .A4(new_n458), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n462), .A2(new_n293), .A3(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT5), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT83), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n467), .B1(new_n468), .B2(G41), .ZN(new_n469));
  INV_X1    g0269(.A(G45), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n470), .A2(G1), .ZN(new_n471));
  INV_X1    g0271(.A(G41), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n472), .A2(KEYINPUT83), .A3(KEYINPUT5), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n469), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n301), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(G264), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n466), .A2(new_n477), .ZN(new_n478));
  OR2_X1    g0278(.A1(new_n474), .A2(new_n298), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(new_n304), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT89), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n478), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n466), .A2(KEYINPUT89), .A3(new_n477), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n480), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n482), .B1(new_n486), .B2(G200), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n294), .A2(new_n266), .A3(G87), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT22), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n266), .A2(G107), .ZN(new_n490));
  OR2_X1    g0290(.A1(new_n490), .A2(KEYINPUT23), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(KEYINPUT23), .ZN(new_n492));
  AOI22_X1  g0292(.A1(new_n488), .A2(new_n489), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n385), .A2(KEYINPUT22), .A3(new_n266), .A4(G87), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n266), .A2(G33), .A3(G116), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  OR2_X1    g0296(.A1(new_n496), .A2(KEYINPUT24), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(KEYINPUT24), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n275), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n272), .A2(G1), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n490), .ZN(new_n501));
  AND2_X1   g0301(.A1(new_n501), .A2(KEYINPUT25), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT81), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n264), .A2(G1), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n273), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n504), .A2(new_n503), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n506), .A2(new_n271), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(G107), .ZN(new_n509));
  OAI22_X1  g0309(.A1(new_n508), .A2(new_n509), .B1(KEYINPUT25), .B2(new_n501), .ZN(new_n510));
  NOR3_X1   g0310(.A1(new_n499), .A2(new_n502), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n487), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(G33), .A2(G116), .ZN(new_n513));
  AOI22_X1  g0313(.A1(new_n288), .A2(G238), .B1(G244), .B2(G1698), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n513), .B1(new_n514), .B2(new_n401), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n515), .A2(KEYINPUT84), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT84), .ZN(new_n517));
  OAI22_X1  g0317(.A1(new_n357), .A2(new_n220), .B1(new_n221), .B2(new_n291), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(new_n385), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n517), .B1(new_n519), .B2(new_n513), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n293), .B1(new_n516), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n471), .A2(G274), .ZN(new_n522));
  OR3_X1    g0322(.A1(new_n293), .A2(new_n212), .A3(new_n471), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n521), .A2(G190), .A3(new_n522), .A4(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n508), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(G87), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n265), .A2(G97), .A3(new_n267), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT19), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n266), .B1(new_n325), .B2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(G97), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n211), .A2(new_n530), .A3(new_n509), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n527), .A2(new_n528), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n380), .A2(new_n266), .A3(G68), .A4(new_n381), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n271), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n364), .A2(new_n273), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n526), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n515), .A2(KEYINPUT84), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n519), .A2(new_n517), .A3(new_n513), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n301), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(new_n522), .ZN(new_n542));
  INV_X1    g0342(.A(new_n523), .ZN(new_n543));
  NOR3_X1   g0343(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n524), .B(new_n538), .C1(new_n544), .C2(new_n353), .ZN(new_n545));
  OAI211_X1 g0345(.A(KEYINPUT4), .B(G244), .C1(new_n355), .C2(new_n356), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n546), .B1(new_n212), .B2(new_n291), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n294), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n380), .A2(G244), .A3(new_n288), .A4(new_n381), .ZN(new_n549));
  XOR2_X1   g0349(.A(KEYINPUT82), .B(KEYINPUT4), .Z(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(G33), .A2(G283), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n548), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n293), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n476), .A2(G257), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n554), .A2(new_n397), .A3(new_n555), .A4(new_n479), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n423), .A2(G97), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n525), .A2(G97), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n509), .B1(new_n417), .B2(new_n418), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n261), .A2(new_n342), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT6), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n530), .A2(new_n509), .ZN(new_n563));
  NOR2_X1   g0363(.A1(G97), .A2(G107), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n509), .A2(KEYINPUT6), .A3(G97), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n266), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NOR3_X1   g0367(.A1(new_n560), .A2(new_n561), .A3(new_n567), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n558), .B(new_n559), .C1(new_n568), .C2(new_n275), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n556), .A2(new_n569), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n553), .A2(new_n293), .B1(G257), .B2(new_n476), .ZN(new_n571));
  AOI21_X1  g0371(.A(G169), .B1(new_n571), .B2(new_n479), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n521), .A2(new_n397), .A3(new_n522), .A4(new_n523), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n535), .B(new_n536), .C1(new_n364), .C2(new_n508), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n575), .B(new_n576), .C1(new_n544), .C2(G169), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n571), .A2(new_n479), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(G200), .ZN(new_n579));
  INV_X1    g0379(.A(new_n569), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n579), .B(new_n580), .C1(new_n304), .C2(new_n578), .ZN(new_n581));
  AND4_X1   g0381(.A1(new_n545), .A2(new_n574), .A3(new_n577), .A4(new_n581), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n479), .B1(new_n217), .B2(new_n475), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT85), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n479), .B(KEYINPUT85), .C1(new_n217), .C2(new_n475), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n288), .A2(G257), .B1(G264), .B2(G1698), .ZN(new_n588));
  INV_X1    g0388(.A(G303), .ZN(new_n589));
  OAI22_X1  g0389(.A1(new_n588), .A2(new_n401), .B1(new_n589), .B2(new_n294), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n293), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT86), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n590), .A2(KEYINPUT86), .A3(new_n293), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n587), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n273), .A2(new_n216), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n552), .B(new_n266), .C1(G33), .C2(new_n530), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n597), .B(new_n271), .C1(new_n266), .C2(G116), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT20), .ZN(new_n599));
  AND2_X1   g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n598), .A2(new_n599), .ZN(new_n601));
  OAI221_X1 g0401(.A(new_n596), .B1(new_n508), .B2(new_n216), .C1(new_n600), .C2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n595), .A2(G169), .A3(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT21), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n595), .A2(G200), .ZN(new_n606));
  INV_X1    g0406(.A(new_n602), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n606), .B(new_n607), .C1(new_n304), .C2(new_n595), .ZN(new_n608));
  AND4_X1   g0408(.A1(G179), .A2(new_n587), .A3(new_n593), .A4(new_n594), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n602), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n595), .A2(KEYINPUT21), .A3(G169), .A4(new_n602), .ZN(new_n611));
  AND4_X1   g0411(.A1(new_n605), .A2(new_n608), .A3(new_n610), .A4(new_n611), .ZN(new_n612));
  AND3_X1   g0412(.A1(new_n466), .A2(KEYINPUT89), .A3(new_n477), .ZN(new_n613));
  AOI21_X1  g0413(.A(KEYINPUT89), .B1(new_n466), .B2(new_n477), .ZN(new_n614));
  OAI211_X1 g0414(.A(G179), .B(new_n479), .C1(new_n613), .C2(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(G169), .B1(new_n478), .B2(new_n480), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n511), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n512), .A2(new_n582), .A3(new_n612), .A4(new_n619), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n450), .A2(new_n620), .ZN(G372));
  INV_X1    g0421(.A(new_n317), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n311), .A2(new_n313), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n432), .B1(new_n443), .B2(new_n444), .ZN(new_n624));
  XNOR2_X1  g0424(.A(new_n624), .B(KEYINPUT18), .ZN(new_n625));
  INV_X1    g0425(.A(new_n371), .ZN(new_n626));
  AOI22_X1  g0426(.A1(new_n354), .A2(new_n626), .B1(new_n340), .B2(new_n350), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n437), .A2(new_n440), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n625), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n622), .B1(new_n623), .B2(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n545), .A2(new_n573), .A3(new_n577), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(KEYINPUT26), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n632), .A2(new_n577), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(G200), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT90), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n537), .A2(new_n636), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n526), .A2(new_n535), .A3(KEYINPUT90), .A4(new_n536), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n635), .A2(new_n639), .A3(new_n524), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n577), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT26), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n642), .A2(new_n643), .A3(new_n573), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n574), .A2(new_n581), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n479), .B1(new_n613), .B2(new_n614), .ZN(new_n646));
  AOI22_X1  g0446(.A1(new_n646), .A2(new_n353), .B1(new_n304), .B2(new_n481), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n645), .B(new_n640), .C1(new_n647), .C2(new_n618), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n511), .B1(new_n615), .B2(new_n616), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n605), .A2(new_n610), .A3(new_n611), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n577), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  OAI211_X1 g0451(.A(new_n633), .B(new_n644), .C1(new_n648), .C2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n630), .B1(new_n450), .B2(new_n653), .ZN(G369));
  NOR2_X1   g0454(.A1(new_n272), .A2(G20), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n296), .ZN(new_n656));
  OR2_X1    g0456(.A1(new_n656), .A2(KEYINPUT27), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(KEYINPUT27), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n657), .A2(G213), .A3(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(G343), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n618), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n512), .A2(new_n619), .A3(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n650), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n664), .A2(new_n661), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n649), .A2(new_n661), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n663), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n649), .B1(new_n511), .B2(new_n487), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(new_n665), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n661), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n607), .A2(new_n672), .ZN(new_n673));
  MUX2_X1   g0473(.A(new_n612), .B(new_n650), .S(new_n673), .Z(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(G330), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  AOI22_X1  g0477(.A1(new_n669), .A2(new_n665), .B1(new_n649), .B2(new_n672), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(G399));
  INV_X1    g0479(.A(KEYINPUT91), .ZN(new_n680));
  INV_X1    g0480(.A(new_n230), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n680), .B1(new_n681), .B2(G41), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n230), .A2(KEYINPUT91), .A3(new_n472), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n531), .A2(G116), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n684), .A2(G1), .A3(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n234), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n686), .B1(new_n687), .B2(new_n684), .ZN(new_n688));
  XNOR2_X1  g0488(.A(new_n688), .B(KEYINPUT28), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT30), .ZN(new_n690));
  OAI211_X1 g0490(.A(new_n609), .B(new_n479), .C1(new_n613), .C2(new_n614), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n544), .A2(new_n571), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n690), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT93), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n692), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n486), .A2(KEYINPUT30), .A3(new_n609), .A4(new_n696), .ZN(new_n697));
  OAI211_X1 g0497(.A(KEYINPUT93), .B(new_n690), .C1(new_n691), .C2(new_n692), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n695), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  AND3_X1   g0499(.A1(new_n634), .A2(new_n595), .A3(new_n397), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n646), .A2(new_n700), .A3(new_n578), .ZN(new_n701));
  XNOR2_X1  g0501(.A(new_n701), .B(KEYINPUT94), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n661), .B1(new_n699), .B2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT31), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n693), .A2(new_n697), .A3(new_n701), .ZN(new_n706));
  XOR2_X1   g0506(.A(KEYINPUT92), .B(KEYINPUT31), .Z(new_n707));
  NAND3_X1  g0507(.A1(new_n706), .A2(new_n661), .A3(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n708), .B1(new_n620), .B2(new_n661), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n705), .A2(new_n710), .ZN(new_n711));
  AND2_X1   g0511(.A1(new_n711), .A2(G330), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n631), .A2(new_n643), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT95), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n640), .A2(KEYINPUT26), .A3(new_n577), .A4(new_n573), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n713), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  OR2_X1    g0516(.A1(new_n715), .A2(new_n714), .ZN(new_n717));
  AND3_X1   g0517(.A1(new_n716), .A2(new_n717), .A3(new_n577), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n619), .A2(KEYINPUT96), .A3(new_n664), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT96), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n720), .B1(new_n649), .B2(new_n650), .ZN(new_n721));
  INV_X1    g0521(.A(new_n640), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n722), .B1(new_n487), .B2(new_n511), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n719), .A2(new_n721), .A3(new_n723), .A4(new_n645), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n718), .A2(new_n724), .ZN(new_n725));
  AND4_X1   g0525(.A1(KEYINPUT97), .A2(new_n725), .A3(KEYINPUT29), .A4(new_n672), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n661), .B1(new_n718), .B2(new_n724), .ZN(new_n727));
  AOI21_X1  g0527(.A(KEYINPUT97), .B1(new_n727), .B2(KEYINPUT29), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n652), .A2(new_n672), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT29), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n712), .B1(new_n729), .B2(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n689), .B1(new_n733), .B2(G1), .ZN(G364));
  INV_X1    g0534(.A(new_n684), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n655), .A2(G45), .ZN(new_n736));
  OR2_X1    g0536(.A1(new_n736), .A2(KEYINPUT98), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(KEYINPUT98), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n737), .A2(G1), .A3(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n735), .A2(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n740), .B1(new_n674), .B2(G330), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n741), .B1(G330), .B2(new_n674), .ZN(new_n742));
  NAND2_X1  g0542(.A1(G20), .A2(G179), .ZN(new_n743));
  XOR2_X1   g0543(.A(new_n743), .B(KEYINPUT99), .Z(new_n744));
  NAND3_X1  g0544(.A1(new_n744), .A2(G190), .A3(new_n353), .ZN(new_n745));
  INV_X1    g0545(.A(G322), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(G179), .A2(G200), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n748), .A2(G20), .A3(new_n304), .ZN(new_n749));
  INV_X1    g0549(.A(G329), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n353), .A2(G179), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n751), .A2(G20), .A3(G190), .ZN(new_n752));
  OAI221_X1 g0552(.A(new_n287), .B1(new_n749), .B2(new_n750), .C1(new_n752), .C2(new_n589), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n744), .A2(G190), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(new_n353), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n753), .B1(new_n755), .B2(G326), .ZN(new_n756));
  INV_X1    g0556(.A(G283), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n751), .A2(G20), .A3(new_n304), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n756), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  AND3_X1   g0559(.A1(new_n744), .A2(new_n304), .A3(G200), .ZN(new_n760));
  XNOR2_X1  g0560(.A(KEYINPUT33), .B(G317), .ZN(new_n761));
  AOI211_X1 g0561(.A(new_n747), .B(new_n759), .C1(new_n760), .C2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(G294), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n266), .B1(new_n748), .B2(G190), .ZN(new_n764));
  OR2_X1    g0564(.A1(new_n764), .A2(KEYINPUT102), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(KEYINPUT102), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(G311), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n744), .A2(new_n304), .A3(new_n353), .ZN(new_n769));
  INV_X1    g0569(.A(KEYINPUT101), .ZN(new_n770));
  AND2_X1   g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n769), .A2(new_n770), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  OAI221_X1 g0573(.A(new_n762), .B1(new_n763), .B2(new_n767), .C1(new_n768), .C2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n760), .ZN(new_n775));
  OAI22_X1  g0575(.A1(new_n775), .A2(new_n202), .B1(new_n530), .B2(new_n767), .ZN(new_n776));
  INV_X1    g0576(.A(new_n752), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G87), .ZN(new_n778));
  INV_X1    g0578(.A(G159), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n749), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n780), .B(KEYINPUT32), .ZN(new_n781));
  INV_X1    g0581(.A(new_n755), .ZN(new_n782));
  OAI211_X1 g0582(.A(new_n778), .B(new_n781), .C1(new_n782), .C2(new_n214), .ZN(new_n783));
  XOR2_X1   g0583(.A(new_n745), .B(KEYINPUT100), .Z(new_n784));
  AOI211_X1 g0584(.A(new_n776), .B(new_n783), .C1(G58), .C2(new_n784), .ZN(new_n785));
  OAI221_X1 g0585(.A(new_n785), .B1(new_n509), .B2(new_n758), .C1(new_n223), .C2(new_n773), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n774), .B1(new_n786), .B2(new_n287), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n235), .B1(G20), .B2(new_n315), .ZN(new_n788));
  NOR2_X1   g0588(.A1(G13), .A2(G33), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(G20), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(new_n788), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n385), .A2(new_n681), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n234), .A2(new_n470), .ZN(new_n794));
  OAI211_X1 g0594(.A(new_n793), .B(new_n794), .C1(new_n252), .C2(new_n470), .ZN(new_n795));
  INV_X1    g0595(.A(G355), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n294), .A2(new_n230), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n795), .B1(G116), .B2(new_n230), .C1(new_n796), .C2(new_n797), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n787), .A2(new_n788), .B1(new_n792), .B2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n791), .ZN(new_n800));
  OAI211_X1 g0600(.A(new_n799), .B(new_n740), .C1(new_n674), .C2(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n742), .A2(new_n801), .ZN(G396));
  NOR2_X1   g0602(.A1(new_n368), .A2(new_n672), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n371), .B1(new_n377), .B2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n371), .A2(new_n661), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n730), .A2(new_n807), .ZN(new_n808));
  AND2_X1   g0608(.A1(new_n804), .A2(new_n806), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n652), .A2(new_n809), .A3(new_n672), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n712), .B(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n740), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n758), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(G68), .ZN(new_n816));
  OAI221_X1 g0616(.A(new_n816), .B1(new_n214), .B2(new_n752), .C1(new_n767), .C2(new_n201), .ZN(new_n817));
  INV_X1    g0617(.A(G132), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n784), .A2(G143), .B1(G150), .B2(new_n760), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n819), .B1(new_n779), .B2(new_n773), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n820), .B1(G137), .B2(new_n755), .ZN(new_n821));
  XOR2_X1   g0621(.A(new_n821), .B(KEYINPUT104), .Z(new_n822));
  INV_X1    g0622(.A(KEYINPUT34), .ZN(new_n823));
  OAI221_X1 g0623(.A(new_n385), .B1(new_n818), .B2(new_n749), .C1(new_n822), .C2(new_n823), .ZN(new_n824));
  AOI211_X1 g0624(.A(new_n817), .B(new_n824), .C1(new_n823), .C2(new_n822), .ZN(new_n825));
  INV_X1    g0625(.A(new_n767), .ZN(new_n826));
  AOI22_X1  g0626(.A1(G303), .A2(new_n755), .B1(new_n826), .B2(G97), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(new_n763), .B2(new_n745), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n773), .A2(new_n216), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n294), .B1(new_n777), .B2(G107), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT103), .ZN(new_n831));
  INV_X1    g0631(.A(new_n749), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n830), .A2(new_n831), .B1(G311), .B2(new_n832), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n833), .B1(new_n831), .B2(new_n830), .C1(new_n211), .C2(new_n758), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n775), .A2(new_n757), .ZN(new_n835));
  NOR4_X1   g0635(.A1(new_n828), .A2(new_n829), .A3(new_n834), .A4(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n788), .B1(new_n825), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n807), .A2(new_n789), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n788), .A2(new_n789), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(new_n342), .ZN(new_n840));
  NAND4_X1  g0640(.A1(new_n837), .A2(new_n740), .A3(new_n838), .A4(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n814), .A2(new_n841), .ZN(G384));
  NAND2_X1  g0642(.A1(new_n350), .A2(new_n661), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n351), .A2(new_n354), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(KEYINPUT105), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT105), .ZN(new_n846));
  NAND4_X1  g0646(.A1(new_n351), .A2(new_n846), .A3(new_n354), .A4(new_n843), .ZN(new_n847));
  OAI21_X1  g0647(.A(KEYINPUT106), .B1(new_n351), .B2(new_n672), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT106), .ZN(new_n849));
  NAND4_X1  g0649(.A1(new_n340), .A2(new_n849), .A3(new_n350), .A4(new_n661), .ZN(new_n850));
  AOI22_X1  g0650(.A1(new_n845), .A2(new_n847), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  NAND4_X1  g0651(.A1(new_n669), .A2(new_n582), .A3(new_n612), .A4(new_n672), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(new_n707), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(new_n703), .ZN(new_n854));
  OAI211_X1 g0654(.A(KEYINPUT31), .B(new_n661), .C1(new_n699), .C2(new_n702), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n807), .B(new_n851), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT40), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT38), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n445), .A2(new_n438), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n439), .A2(new_n434), .ZN(new_n860));
  INV_X1    g0660(.A(new_n659), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n861), .B1(new_n427), .B2(new_n428), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n859), .A2(new_n860), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(KEYINPUT37), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n442), .B1(new_n445), .B2(new_n861), .ZN(new_n865));
  AOI21_X1  g0665(.A(KEYINPUT37), .B1(new_n439), .B2(new_n434), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AND2_X1   g0667(.A1(new_n864), .A2(new_n867), .ZN(new_n868));
  AND2_X1   g0668(.A1(new_n437), .A2(new_n440), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n862), .B1(new_n625), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n858), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n409), .B1(new_n412), .B2(new_n413), .ZN(new_n872));
  AND2_X1   g0672(.A1(new_n872), .A2(new_n415), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n414), .A2(new_n271), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n425), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n861), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n448), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n445), .A2(new_n875), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n879), .A2(new_n860), .A3(new_n876), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(KEYINPUT37), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(new_n867), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n878), .A2(new_n882), .A3(KEYINPUT38), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n857), .B1(new_n871), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n845), .A2(new_n847), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n848), .A2(new_n850), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n807), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  AND3_X1   g0687(.A1(new_n442), .A2(new_n445), .A3(new_n446), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n446), .B1(new_n442), .B2(new_n445), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n876), .B1(new_n890), .B2(new_n869), .ZN(new_n891));
  AOI22_X1  g0691(.A1(new_n880), .A2(KEYINPUT37), .B1(new_n866), .B2(new_n865), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n858), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(new_n883), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT94), .ZN(new_n895));
  XNOR2_X1  g0695(.A(new_n701), .B(new_n895), .ZN(new_n896));
  NAND4_X1  g0696(.A1(new_n896), .A2(new_n697), .A3(new_n695), .A4(new_n698), .ZN(new_n897));
  AOI22_X1  g0697(.A1(new_n897), .A2(new_n661), .B1(new_n852), .B2(new_n707), .ZN(new_n898));
  INV_X1    g0698(.A(new_n855), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n887), .B(new_n894), .C1(new_n898), .C2(new_n899), .ZN(new_n900));
  AOI22_X1  g0700(.A1(new_n856), .A2(new_n884), .B1(new_n900), .B2(new_n857), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n854), .A2(new_n855), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(new_n449), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n901), .B(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(G330), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n725), .A2(KEYINPUT29), .A3(new_n672), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT97), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n727), .A2(KEYINPUT97), .A3(KEYINPUT29), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n908), .A2(new_n449), .A3(new_n732), .A4(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n630), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT39), .ZN(new_n912));
  NOR3_X1   g0712(.A1(new_n891), .A2(new_n858), .A3(new_n892), .ZN(new_n913));
  INV_X1    g0713(.A(new_n862), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n624), .B(new_n446), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n914), .B1(new_n915), .B2(new_n628), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n864), .A2(new_n867), .ZN(new_n917));
  AOI21_X1  g0717(.A(KEYINPUT38), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n912), .B1(new_n913), .B2(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n351), .A2(new_n661), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n893), .A2(KEYINPUT39), .A3(new_n883), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n810), .A2(new_n806), .ZN(new_n923));
  INV_X1    g0723(.A(new_n851), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n923), .A2(new_n894), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n915), .A2(new_n659), .ZN(new_n926));
  AND3_X1   g0726(.A1(new_n922), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n911), .B(new_n927), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n905), .B(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(new_n296), .B2(new_n655), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n565), .A2(new_n566), .ZN(new_n931));
  OAI211_X1 g0731(.A(G20), .B(new_n236), .C1(new_n931), .C2(KEYINPUT35), .ZN(new_n932));
  AOI211_X1 g0732(.A(new_n216), .B(new_n932), .C1(KEYINPUT35), .C2(new_n931), .ZN(new_n933));
  XOR2_X1   g0733(.A(new_n933), .B(KEYINPUT36), .Z(new_n934));
  OAI21_X1  g0734(.A(new_n222), .B1(new_n201), .B2(new_n202), .ZN(new_n935));
  OAI22_X1  g0735(.A1(new_n687), .A2(new_n935), .B1(G50), .B2(new_n202), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n936), .A2(G1), .A3(new_n272), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n930), .A2(new_n934), .A3(new_n937), .ZN(G367));
  NAND2_X1  g0738(.A1(new_n777), .A2(G116), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT46), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n832), .A2(G317), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n940), .B(new_n941), .C1(new_n530), .C2(new_n758), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n401), .B1(new_n782), .B2(new_n768), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n944), .B1(new_n763), .B2(new_n775), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n945), .B1(G303), .B2(new_n784), .ZN(new_n946));
  OAI221_X1 g0746(.A(new_n946), .B1(new_n509), .B2(new_n767), .C1(new_n757), .C2(new_n773), .ZN(new_n947));
  INV_X1    g0747(.A(G143), .ZN(new_n948));
  OAI22_X1  g0748(.A1(new_n782), .A2(new_n948), .B1(new_n202), .B2(new_n767), .ZN(new_n949));
  AND2_X1   g0749(.A1(new_n832), .A2(G137), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n745), .A2(new_n259), .ZN(new_n951));
  OAI221_X1 g0751(.A(new_n294), .B1(new_n752), .B2(new_n201), .C1(new_n223), .C2(new_n758), .ZN(new_n952));
  NOR4_X1   g0752(.A1(new_n949), .A2(new_n950), .A3(new_n951), .A4(new_n952), .ZN(new_n953));
  OAI221_X1 g0753(.A(new_n953), .B1(new_n214), .B2(new_n773), .C1(new_n779), .C2(new_n775), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n947), .A2(new_n954), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(KEYINPUT47), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n813), .B1(new_n956), .B2(new_n788), .ZN(new_n957));
  INV_X1    g0757(.A(new_n793), .ZN(new_n958));
  OAI221_X1 g0758(.A(new_n792), .B1(new_n230), .B2(new_n364), .C1(new_n958), .C2(new_n248), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n637), .A2(new_n638), .A3(new_n661), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n642), .A2(new_n960), .ZN(new_n961));
  OR2_X1    g0761(.A1(new_n577), .A2(new_n960), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n961), .A2(new_n791), .A3(new_n962), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n957), .A2(new_n959), .A3(new_n963), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n908), .A2(new_n732), .A3(new_n909), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n711), .A2(G330), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT108), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n671), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n668), .A2(KEYINPUT108), .A3(new_n670), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n969), .A2(new_n675), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(KEYINPUT109), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT109), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n969), .A2(new_n973), .A3(new_n675), .A4(new_n970), .ZN(new_n974));
  AND3_X1   g0774(.A1(new_n972), .A2(new_n677), .A3(new_n974), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n574), .B(new_n581), .C1(new_n580), .C2(new_n672), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n573), .A2(new_n661), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OR3_X1    g0778(.A1(new_n678), .A2(KEYINPUT44), .A3(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(KEYINPUT44), .B1(new_n678), .B2(new_n978), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  AND3_X1   g0781(.A1(new_n678), .A2(KEYINPUT45), .A3(new_n978), .ZN(new_n982));
  AOI21_X1  g0782(.A(KEYINPUT45), .B1(new_n678), .B2(new_n978), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n981), .A2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n967), .B1(new_n975), .B2(new_n986), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n684), .B(KEYINPUT41), .Z(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(KEYINPUT110), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n972), .A2(new_n677), .A3(new_n974), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n733), .B1(new_n991), .B2(new_n985), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT110), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n992), .A2(new_n993), .A3(new_n988), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n739), .B1(new_n990), .B2(new_n994), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n670), .A2(new_n976), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT42), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n574), .B1(new_n619), .B2(new_n976), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n998), .B(KEYINPUT107), .Z(new_n999));
  NAND2_X1  g0799(.A1(new_n999), .A2(new_n672), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n961), .A2(new_n962), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n997), .A2(new_n1000), .B1(KEYINPUT43), .B2(new_n1001), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n1001), .A2(KEYINPUT43), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1002), .B(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n978), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n677), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1004), .B(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n964), .B1(new_n995), .B2(new_n1008), .ZN(G387));
  NAND2_X1  g0809(.A1(new_n975), .A2(new_n739), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n755), .A2(G159), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT111), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n767), .A2(new_n364), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n745), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1013), .B1(G50), .B2(new_n1014), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n758), .A2(new_n530), .B1(new_n259), .B2(new_n749), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n262), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1016), .B1(new_n760), .B2(new_n1017), .ZN(new_n1018));
  AND3_X1   g0818(.A1(new_n1012), .A2(new_n1015), .A3(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n777), .A2(new_n222), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n773), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1021), .A2(G68), .ZN(new_n1022));
  NAND4_X1  g0822(.A1(new_n1019), .A2(new_n385), .A3(new_n1020), .A4(new_n1022), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n784), .A2(G317), .B1(G311), .B2(new_n760), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n1024), .B1(new_n589), .B2(new_n773), .C1(new_n746), .C2(new_n782), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT48), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n1026), .B1(new_n757), .B2(new_n767), .C1(new_n763), .C2(new_n752), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT49), .ZN(new_n1028));
  OR2_X1    g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n385), .B1(G326), .B2(new_n832), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n758), .A2(new_n216), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1023), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n793), .B1(new_n245), .B2(new_n470), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n685), .B2(new_n797), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n202), .A2(new_n342), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1017), .A2(new_n214), .ZN(new_n1038));
  AOI211_X1 g0838(.A(G116), .B(new_n531), .C1(new_n1038), .C2(KEYINPUT50), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1039), .B(new_n470), .C1(KEYINPUT50), .C2(new_n1038), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1036), .B1(new_n1037), .B2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1041), .B1(G107), .B2(new_n230), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n1034), .A2(new_n788), .B1(new_n792), .B2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n663), .A2(new_n667), .A3(new_n791), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n735), .B1(new_n975), .B2(new_n733), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n991), .A2(new_n967), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n1010), .B1(new_n1045), .B2(new_n813), .C1(new_n1046), .C2(new_n1047), .ZN(G393));
  OAI21_X1  g0848(.A(new_n676), .B1(new_n981), .B2(new_n984), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n983), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n678), .A2(KEYINPUT45), .A3(new_n978), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND4_X1  g0852(.A1(new_n1052), .A2(new_n677), .A3(new_n980), .A4(new_n979), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1049), .A2(new_n1053), .A3(new_n739), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(G317), .A2(new_n755), .B1(new_n1014), .B2(G311), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT52), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n758), .A2(new_n509), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n777), .A2(G283), .B1(new_n832), .B2(G322), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n287), .B1(new_n1058), .B2(KEYINPUT113), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n1057), .B(new_n1059), .C1(KEYINPUT113), .C2(new_n1058), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n1060), .B1(new_n216), .B2(new_n767), .C1(new_n763), .C2(new_n773), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n1056), .B(new_n1061), .C1(G303), .C2(new_n760), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(G150), .A2(new_n755), .B1(new_n1014), .B2(G159), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT51), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n758), .A2(new_n211), .B1(new_n948), .B2(new_n749), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n401), .B(new_n1065), .C1(G68), .C2(new_n777), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1066), .ZN(new_n1067));
  OR2_X1    g0867(.A1(new_n1067), .A2(KEYINPUT112), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n826), .A2(G77), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1067), .A2(KEYINPUT112), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n760), .A2(G50), .ZN(new_n1071));
  NAND4_X1  g0871(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .A4(new_n1071), .ZN(new_n1072));
  AOI211_X1 g0872(.A(new_n1064), .B(new_n1072), .C1(new_n1017), .C2(new_n1021), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n788), .B1(new_n1062), .B2(new_n1073), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n792), .B1(new_n530), .B2(new_n230), .C1(new_n958), .C2(new_n255), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1074), .A2(new_n740), .A3(new_n1075), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT114), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1077), .B1(new_n800), .B2(new_n978), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1049), .A2(new_n1053), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n991), .B2(new_n967), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n735), .ZN(new_n1081));
  NOR3_X1   g0881(.A1(new_n991), .A2(new_n967), .A3(new_n985), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n1054), .B(new_n1078), .C1(new_n1081), .C2(new_n1082), .ZN(G390));
  OAI22_X1  g0883(.A1(new_n773), .A2(new_n530), .B1(new_n509), .B2(new_n775), .ZN(new_n1084));
  XOR2_X1   g0884(.A(new_n1084), .B(KEYINPUT115), .Z(new_n1085));
  NAND2_X1  g0885(.A1(new_n832), .A2(G294), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n778), .A2(new_n816), .A3(new_n287), .A4(new_n1086), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n1069), .B1(new_n216), .B2(new_n745), .C1(new_n782), .C2(new_n757), .ZN(new_n1088));
  NOR3_X1   g0888(.A1(new_n1085), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n826), .A2(G159), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(KEYINPUT54), .B(G143), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n773), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n760), .A2(G137), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n752), .A2(new_n259), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1094), .B(KEYINPUT53), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n815), .A2(G50), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n287), .B1(new_n832), .B2(G125), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n1093), .A2(new_n1095), .A3(new_n1096), .A4(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(G128), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n782), .A2(new_n1099), .B1(new_n818), .B2(new_n745), .ZN(new_n1100));
  NOR3_X1   g0900(.A1(new_n1092), .A2(new_n1098), .A3(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1089), .B1(new_n1090), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n1103), .A2(new_n788), .B1(new_n262), .B2(new_n839), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n921), .ZN(new_n1105));
  AOI21_X1  g0905(.A(KEYINPUT39), .B1(new_n871), .B2(new_n883), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n740), .B(new_n1104), .C1(new_n1107), .C2(new_n790), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n851), .B1(new_n810), .B2(new_n806), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n1109), .A2(new_n920), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n920), .B1(new_n871), .B2(new_n883), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n805), .B1(new_n727), .B2(new_n804), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1111), .B1(new_n1112), .B2(new_n851), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n809), .A2(G330), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(KEYINPUT31), .B1(new_n897), .B2(new_n661), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n924), .B(new_n1115), .C1(new_n1116), .C2(new_n709), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  AND3_X1   g0918(.A1(new_n1110), .A2(new_n1113), .A3(new_n1118), .ZN(new_n1119));
  AOI211_X1 g0919(.A(new_n851), .B(new_n1114), .C1(new_n854), .C2(new_n855), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1120), .B1(new_n1110), .B2(new_n1113), .ZN(new_n1121));
  OR2_X1    g0921(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n739), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1108), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n902), .A2(new_n449), .A3(G330), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n910), .A2(new_n630), .A3(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n924), .B1(new_n711), .B2(new_n1115), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n923), .B1(new_n1120), .B2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1114), .B1(new_n854), .B2(new_n855), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n1117), .B(new_n1112), .C1(new_n1131), .C2(new_n924), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1128), .B(new_n1133), .C1(new_n1119), .C2(new_n1121), .ZN(new_n1134));
  AND2_X1   g0934(.A1(new_n1134), .A2(new_n735), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1128), .A2(new_n1133), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1123), .A2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1125), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(G378));
  INV_X1    g0939(.A(KEYINPUT118), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(KEYINPUT117), .B(KEYINPUT56), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT55), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n623), .A2(new_n1143), .A3(new_n317), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n318), .A2(KEYINPUT55), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n307), .A2(new_n659), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  AND3_X1   g0947(.A1(new_n1144), .A2(new_n1145), .A3(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1147), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1142), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(new_n1146), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1144), .A2(new_n1145), .A3(new_n1147), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1152), .A2(new_n1141), .A3(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1150), .A2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n922), .A2(new_n925), .A3(new_n926), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1156), .B1(new_n901), .B2(G330), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n900), .A2(new_n857), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n902), .A2(new_n887), .A3(new_n884), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1158), .A2(G330), .A3(new_n1159), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1160), .A2(new_n927), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1155), .B1(new_n1157), .B2(new_n1161), .ZN(new_n1162));
  AND2_X1   g0962(.A1(new_n1150), .A2(new_n1154), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1160), .A2(new_n927), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n1156), .A2(G330), .A3(new_n1158), .A4(new_n1159), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1163), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n1162), .A2(new_n1166), .B1(new_n1134), .B2(new_n1128), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1140), .B1(new_n1167), .B2(KEYINPUT57), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n684), .B1(new_n1167), .B2(KEYINPUT57), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT57), .ZN(new_n1170));
  AND3_X1   g0970(.A1(new_n1163), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1163), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1127), .B1(new_n1122), .B2(new_n1133), .ZN(new_n1174));
  OAI211_X1 g0974(.A(KEYINPUT118), .B(new_n1170), .C1(new_n1173), .C2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1168), .A2(new_n1169), .A3(new_n1175), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n739), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n839), .A2(new_n214), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(G125), .A2(new_n755), .B1(new_n826), .B2(G150), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(new_n1179), .B(KEYINPUT116), .ZN(new_n1180));
  OAI22_X1  g0980(.A1(new_n745), .A2(new_n1099), .B1(new_n752), .B2(new_n1091), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1181), .B1(new_n1021), .B2(G137), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1180), .B(new_n1182), .C1(new_n818), .C2(new_n775), .ZN(new_n1183));
  XOR2_X1   g0983(.A(new_n1183), .B(KEYINPUT59), .Z(new_n1184));
  AOI21_X1  g0984(.A(G41), .B1(new_n832), .B2(G124), .ZN(new_n1185));
  AOI21_X1  g0985(.A(G33), .B1(new_n815), .B2(G159), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n782), .A2(new_n216), .B1(new_n775), .B2(new_n530), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n401), .B1(new_n767), .B2(new_n202), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n815), .A2(G58), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n832), .A2(G283), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1020), .A2(new_n1190), .A3(new_n472), .A4(new_n1191), .ZN(new_n1192));
  NOR3_X1   g0992(.A1(new_n1188), .A2(new_n1189), .A3(new_n1192), .ZN(new_n1193));
  OAI221_X1 g0993(.A(new_n1193), .B1(new_n509), .B2(new_n745), .C1(new_n364), .C2(new_n773), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(new_n1194), .B(KEYINPUT58), .ZN(new_n1195));
  AOI21_X1  g0995(.A(G41), .B1(new_n385), .B2(G33), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1187), .B(new_n1195), .C1(G50), .C2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n813), .B1(new_n1197), .B2(new_n788), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1178), .B(new_n1198), .C1(new_n1155), .C2(new_n790), .ZN(new_n1199));
  AND2_X1   g0999(.A1(new_n1177), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1176), .A2(new_n1200), .ZN(G375));
  NAND2_X1  g1001(.A1(new_n851), .A2(new_n789), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n385), .B1(new_n1099), .B2(new_n749), .ZN(new_n1203));
  OAI221_X1 g1003(.A(new_n1190), .B1(new_n779), .B2(new_n752), .C1(new_n775), .C2(new_n1091), .ZN(new_n1204));
  AOI211_X1 g1004(.A(new_n1203), .B(new_n1204), .C1(G132), .C2(new_n755), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n784), .A2(G137), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1021), .A2(G150), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(G50), .B2(new_n826), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n287), .B1(new_n749), .B2(new_n589), .C1(new_n758), .C2(new_n342), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n1210), .B(new_n1013), .C1(G97), .C2(new_n777), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(G294), .A2(new_n755), .B1(new_n1014), .B2(G283), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1211), .B(new_n1212), .C1(new_n509), .C2(new_n773), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(G116), .B2(new_n760), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n788), .B1(new_n1209), .B2(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n813), .B1(new_n202), .B2(new_n839), .ZN(new_n1216));
  XOR2_X1   g1016(.A(new_n1216), .B(KEYINPUT121), .Z(new_n1217));
  NAND3_X1  g1017(.A1(new_n1202), .A2(new_n1215), .A3(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT120), .ZN(new_n1219));
  XOR2_X1   g1019(.A(new_n739), .B(KEYINPUT119), .Z(new_n1220));
  AOI21_X1  g1020(.A(new_n1219), .B1(new_n1133), .B2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1220), .ZN(new_n1222));
  AOI211_X1 g1022(.A(KEYINPUT120), .B(new_n1222), .C1(new_n1130), .C2(new_n1132), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1218), .B1(new_n1221), .B2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1224), .A2(KEYINPUT122), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1132), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n902), .A2(new_n924), .A3(new_n1115), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n709), .B1(new_n704), .B2(new_n703), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n851), .B1(new_n1228), .B2(new_n1114), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n1227), .A2(new_n1229), .B1(new_n806), .B2(new_n810), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1220), .B1(new_n1226), .B2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(KEYINPUT120), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1133), .A2(new_n1219), .A3(new_n1220), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT122), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1234), .A2(new_n1235), .A3(new_n1218), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1225), .A2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1136), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n988), .B1(new_n1133), .B2(new_n1128), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1237), .B1(new_n1238), .B2(new_n1239), .ZN(G381));
  NOR2_X1   g1040(.A1(G375), .A2(G378), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(G381), .A2(G384), .ZN(new_n1242));
  AND3_X1   g1042(.A1(new_n992), .A2(new_n993), .A3(new_n988), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n993), .B1(new_n992), .B2(new_n988), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1124), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(new_n1004), .B(new_n1006), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(G390), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1247), .A2(new_n964), .A3(new_n1248), .ZN(new_n1249));
  NOR3_X1   g1049(.A1(new_n1249), .A2(G396), .A3(G393), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1241), .A2(new_n1242), .A3(new_n1250), .ZN(G407));
  INV_X1    g1051(.A(G213), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1252), .B1(new_n1241), .B2(new_n660), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(G407), .ZN(G409));
  XNOR2_X1  g1054(.A(G393), .B(G396), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1248), .B1(new_n1247), .B2(new_n964), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n964), .ZN(new_n1258));
  AOI211_X1 g1058(.A(new_n1258), .B(G390), .C1(new_n1245), .C2(new_n1246), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1256), .B1(new_n1257), .B2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT61), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(G387), .A2(G390), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1262), .A2(new_n1255), .A3(new_n1249), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1260), .A2(new_n1261), .A3(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT123), .ZN(new_n1265));
  XNOR2_X1  g1065(.A(new_n1264), .B(new_n1265), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1252), .A2(G343), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1176), .A2(G378), .A3(new_n1200), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1134), .A2(new_n1128), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1220), .B1(new_n1269), .B2(new_n988), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1199), .B1(new_n1270), .B2(new_n1173), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(new_n1138), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1267), .B1(new_n1268), .B2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1267), .A2(G2897), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1127), .A2(new_n1130), .A3(KEYINPUT60), .A4(new_n1132), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1136), .A2(new_n735), .A3(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1133), .ZN(new_n1278));
  AOI21_X1  g1078(.A(KEYINPUT60), .B1(new_n1278), .B2(new_n1127), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1277), .A2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(G384), .B1(new_n1237), .B2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(G384), .ZN(new_n1283));
  AOI211_X1 g1083(.A(new_n1283), .B(new_n1280), .C1(new_n1225), .C2(new_n1236), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1275), .B1(new_n1282), .B2(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1235), .B1(new_n1234), .B2(new_n1218), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1218), .ZN(new_n1287));
  AOI211_X1 g1087(.A(KEYINPUT122), .B(new_n1287), .C1(new_n1232), .C2(new_n1233), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1281), .B1(new_n1286), .B2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(new_n1283), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1237), .A2(G384), .A3(new_n1281), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1290), .A2(new_n1291), .A3(new_n1274), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1285), .A2(new_n1292), .ZN(new_n1293));
  OR2_X1    g1093(.A1(new_n1273), .A2(new_n1293), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1282), .A2(new_n1284), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1273), .A2(KEYINPUT63), .A3(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1273), .A2(new_n1295), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT63), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1266), .A2(new_n1294), .A3(new_n1296), .A4(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT62), .ZN(new_n1301));
  OR2_X1    g1101(.A1(new_n1301), .A2(KEYINPUT124), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(KEYINPUT124), .ZN(new_n1303));
  AND4_X1   g1103(.A1(new_n1273), .A2(new_n1295), .A3(new_n1302), .A4(new_n1303), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1261), .B1(new_n1273), .B2(new_n1293), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1302), .B1(new_n1273), .B2(new_n1295), .ZN(new_n1306));
  NOR3_X1   g1106(.A1(new_n1304), .A2(new_n1305), .A3(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1260), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1263), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1300), .B1(new_n1307), .B2(new_n1310), .ZN(G405));
  INV_X1    g1111(.A(KEYINPUT125), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1268), .A2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1315), .A2(G375), .A3(new_n1138), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1316), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1315), .B1(new_n1138), .B2(G375), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1314), .B1(new_n1317), .B2(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT126), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1320), .B1(new_n1308), .B2(new_n1309), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(G375), .A2(new_n1138), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1322), .A2(new_n1295), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1323), .A2(new_n1313), .A3(new_n1316), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1319), .A2(new_n1321), .A3(new_n1324), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1260), .A2(KEYINPUT126), .A3(new_n1263), .ZN(new_n1326));
  XNOR2_X1  g1126(.A(new_n1326), .B(KEYINPUT127), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1325), .A2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT127), .ZN(new_n1329));
  XNOR2_X1  g1129(.A(new_n1326), .B(new_n1329), .ZN(new_n1330));
  NAND4_X1  g1130(.A1(new_n1330), .A2(new_n1321), .A3(new_n1324), .A4(new_n1319), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1328), .A2(new_n1331), .ZN(G402));
endmodule


