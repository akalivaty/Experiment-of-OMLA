//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 0 0 1 1 1 1 1 0 1 0 1 1 1 0 1 1 0 1 0 0 0 1 1 0 1 0 1 1 0 0 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 0 1 1 0 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:11 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n784, new_n785,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n984, new_n985,
    new_n986, new_n987, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026;
  XNOR2_X1  g000(.A(KEYINPUT72), .B(G902), .ZN(new_n187));
  INV_X1    g001(.A(G234), .ZN(new_n188));
  OAI21_X1  g002(.A(G217), .B1(new_n187), .B2(new_n188), .ZN(new_n189));
  XOR2_X1   g003(.A(new_n189), .B(KEYINPUT74), .Z(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT77), .B(KEYINPUT78), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT22), .B(G137), .ZN(new_n193));
  INV_X1    g007(.A(G953), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n194), .A2(G221), .A3(G234), .ZN(new_n195));
  OR2_X1    g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n193), .A2(new_n195), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n192), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n196), .A2(new_n192), .A3(new_n197), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT23), .ZN(new_n202));
  INV_X1    g016(.A(G119), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n202), .B1(new_n203), .B2(G128), .ZN(new_n204));
  INV_X1    g018(.A(G128), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n205), .A2(KEYINPUT23), .A3(G119), .ZN(new_n206));
  OAI211_X1 g020(.A(new_n204), .B(new_n206), .C1(G119), .C2(new_n205), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G110), .ZN(new_n208));
  XOR2_X1   g022(.A(KEYINPUT24), .B(G110), .Z(new_n209));
  XNOR2_X1  g023(.A(G119), .B(G128), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G140), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G125), .ZN(new_n214));
  INV_X1    g028(.A(G125), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G140), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n214), .A2(new_n216), .A3(KEYINPUT75), .ZN(new_n217));
  OR3_X1    g031(.A1(new_n215), .A2(KEYINPUT75), .A3(G140), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n217), .A2(new_n218), .A3(KEYINPUT16), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT16), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n214), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G146), .ZN(new_n223));
  INV_X1    g037(.A(G146), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n219), .A2(new_n224), .A3(new_n221), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n212), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g040(.A(KEYINPUT76), .B(G110), .ZN(new_n227));
  OAI22_X1  g041(.A1(new_n207), .A2(new_n227), .B1(new_n210), .B2(new_n209), .ZN(new_n228));
  XNOR2_X1  g042(.A(G125), .B(G140), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(new_n224), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n224), .B1(new_n219), .B2(new_n221), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n201), .B1(new_n226), .B2(new_n233), .ZN(new_n234));
  AND2_X1   g048(.A1(new_n208), .A2(new_n211), .ZN(new_n235));
  AND3_X1   g049(.A1(new_n219), .A2(new_n224), .A3(new_n221), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n235), .B1(new_n236), .B2(new_n232), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n223), .A2(new_n230), .A3(new_n228), .ZN(new_n238));
  AND3_X1   g052(.A1(new_n196), .A2(new_n192), .A3(new_n197), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n239), .A2(new_n198), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n237), .A2(new_n238), .A3(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n187), .B1(new_n234), .B2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT25), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n191), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n187), .ZN(new_n245));
  AND3_X1   g059(.A1(new_n237), .A2(new_n238), .A3(new_n240), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n240), .B1(new_n237), .B2(new_n238), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n245), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(KEYINPUT25), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n244), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n234), .A2(new_n241), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n190), .A2(G902), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  AND2_X1   g067(.A1(new_n250), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(G143), .ZN(new_n255));
  OAI21_X1  g069(.A(KEYINPUT64), .B1(new_n255), .B2(G146), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT64), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n257), .A2(new_n224), .A3(G143), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n255), .A2(G146), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n256), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n255), .A2(G146), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT1), .ZN(new_n262));
  OAI21_X1  g076(.A(G128), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n260), .A2(new_n263), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n205), .A2(KEYINPUT1), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n256), .A2(new_n258), .A3(new_n259), .A4(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(G104), .ZN(new_n268));
  OAI21_X1  g082(.A(KEYINPUT3), .B1(new_n268), .B2(G107), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT3), .ZN(new_n270));
  INV_X1    g084(.A(G107), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n270), .A2(new_n271), .A3(G104), .ZN(new_n272));
  INV_X1    g086(.A(G101), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n268), .A2(G107), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n269), .A2(new_n272), .A3(new_n273), .A4(new_n274), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n268), .A2(G107), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n271), .A2(G104), .ZN(new_n277));
  OAI21_X1  g091(.A(G101), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  AND2_X1   g092(.A1(new_n275), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n267), .A2(new_n279), .ZN(new_n280));
  XNOR2_X1  g094(.A(KEYINPUT80), .B(KEYINPUT10), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n269), .A2(new_n272), .A3(new_n274), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT79), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n284), .A2(new_n285), .A3(G101), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n286), .A2(KEYINPUT4), .A3(new_n275), .ZN(new_n287));
  NAND2_X1  g101(.A1(KEYINPUT0), .A2(G128), .ZN(new_n288));
  OR2_X1    g102(.A1(KEYINPUT0), .A2(G128), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n224), .A2(G143), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n288), .B(new_n289), .C1(new_n261), .C2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(new_n288), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n256), .A2(new_n258), .A3(new_n292), .A4(new_n259), .ZN(new_n293));
  AND2_X1   g107(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT4), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n284), .A2(new_n285), .A3(new_n295), .A4(G101), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n287), .A2(new_n294), .A3(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G134), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(G137), .ZN(new_n299));
  INV_X1    g113(.A(G137), .ZN(new_n300));
  AOI21_X1  g114(.A(KEYINPUT65), .B1(new_n300), .B2(G134), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT11), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n299), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  AOI211_X1 g117(.A(KEYINPUT65), .B(KEYINPUT11), .C1(new_n300), .C2(G134), .ZN(new_n304));
  NOR3_X1   g118(.A1(new_n303), .A2(G131), .A3(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G131), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n300), .A2(G134), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT65), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n308), .B1(new_n298), .B2(G137), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n307), .B1(new_n309), .B2(KEYINPUT11), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n301), .A2(new_n302), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n306), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n305), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT10), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n262), .B1(G143), .B2(new_n224), .ZN(new_n315));
  OAI22_X1  g129(.A1(new_n315), .A2(new_n205), .B1(new_n261), .B2(new_n290), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n314), .B1(new_n316), .B2(new_n266), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(new_n279), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n283), .A2(new_n297), .A3(new_n313), .A4(new_n318), .ZN(new_n319));
  XNOR2_X1  g133(.A(G110), .B(G140), .ZN(new_n320));
  AND2_X1   g134(.A1(new_n194), .A2(G227), .ZN(new_n321));
  XNOR2_X1  g135(.A(new_n320), .B(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n319), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(new_n313), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n275), .A2(new_n278), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n327), .B1(new_n266), .B2(new_n264), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n318), .B1(new_n328), .B2(new_n281), .ZN(new_n329));
  AND3_X1   g143(.A1(new_n287), .A2(new_n294), .A3(new_n296), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n326), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT12), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n310), .A2(new_n306), .A3(new_n311), .ZN(new_n333));
  OAI21_X1  g147(.A(G131), .B1(new_n303), .B2(new_n304), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n327), .A2(new_n266), .A3(new_n316), .ZN(new_n335));
  AOI221_X4 g149(.A(new_n332), .B1(new_n333), .B2(new_n334), .C1(new_n280), .C2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n280), .A2(new_n335), .ZN(new_n337));
  AOI21_X1  g151(.A(KEYINPUT12), .B1(new_n337), .B2(new_n326), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n319), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  AOI22_X1  g153(.A1(new_n325), .A2(new_n331), .B1(new_n339), .B2(new_n322), .ZN(new_n340));
  OAI21_X1  g154(.A(G469), .B1(new_n340), .B2(G902), .ZN(new_n341));
  INV_X1    g155(.A(G469), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n336), .A2(new_n338), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n343), .A2(new_n324), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n323), .B1(new_n331), .B2(new_n319), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n342), .B(new_n245), .C1(new_n344), .C2(new_n345), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n346), .A2(KEYINPUT81), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT81), .ZN(new_n348));
  INV_X1    g162(.A(new_n319), .ZN(new_n349));
  AOI22_X1  g163(.A1(new_n280), .A2(new_n282), .B1(new_n279), .B2(new_n317), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n313), .B1(new_n350), .B2(new_n297), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n322), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  OAI211_X1 g166(.A(new_n319), .B(new_n323), .C1(new_n336), .C2(new_n338), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n187), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n348), .B1(new_n354), .B2(new_n342), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n341), .B1(new_n347), .B2(new_n355), .ZN(new_n356));
  XNOR2_X1  g170(.A(KEYINPUT9), .B(G234), .ZN(new_n357));
  OAI21_X1  g171(.A(G221), .B1(new_n357), .B2(G902), .ZN(new_n358));
  OAI21_X1  g172(.A(G214), .B1(G237), .B2(G902), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  OAI21_X1  g174(.A(G210), .B1(G237), .B2(G902), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n203), .A2(G116), .ZN(new_n363));
  INV_X1    g177(.A(G116), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(G119), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  XNOR2_X1  g180(.A(KEYINPUT2), .B(G113), .ZN(new_n367));
  OAI21_X1  g181(.A(KEYINPUT66), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(G113), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(KEYINPUT2), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT2), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(G113), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  XNOR2_X1  g187(.A(G116), .B(G119), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT66), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n373), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n368), .A2(new_n376), .ZN(new_n377));
  AND2_X1   g191(.A1(KEYINPUT82), .A2(KEYINPUT5), .ZN(new_n378));
  NOR2_X1   g192(.A1(KEYINPUT82), .A2(KEYINPUT5), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n364), .A2(G119), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n369), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  OAI211_X1 g196(.A(new_n363), .B(new_n365), .C1(new_n378), .C2(new_n379), .ZN(new_n383));
  AOI21_X1  g197(.A(KEYINPUT83), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  OR2_X1    g198(.A1(KEYINPUT82), .A2(KEYINPUT5), .ZN(new_n385));
  NAND2_X1  g199(.A1(KEYINPUT82), .A2(KEYINPUT5), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n381), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  AND4_X1   g201(.A1(KEYINPUT83), .A2(new_n383), .A3(new_n387), .A4(G113), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n377), .B(new_n279), .C1(new_n384), .C2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n366), .A2(new_n367), .ZN(new_n390));
  NOR3_X1   g204(.A1(new_n366), .A2(new_n367), .A3(KEYINPUT66), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n375), .B1(new_n373), .B2(new_n374), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n390), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n393), .A2(new_n287), .A3(new_n296), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n389), .A2(new_n394), .ZN(new_n395));
  XNOR2_X1  g209(.A(G110), .B(G122), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n389), .A2(new_n394), .A3(new_n396), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n398), .A2(KEYINPUT6), .A3(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT6), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n395), .A2(new_n401), .A3(new_n397), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n291), .A2(new_n293), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(G125), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n316), .A2(new_n215), .A3(new_n266), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(G224), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n407), .A2(G953), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n406), .B(new_n408), .ZN(new_n409));
  AND3_X1   g223(.A1(new_n400), .A2(new_n402), .A3(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(G902), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n396), .B(KEYINPUT8), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n377), .B1(new_n384), .B2(new_n388), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT5), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n382), .B1(new_n415), .B2(new_n366), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n416), .A2(new_n377), .A3(new_n279), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT84), .ZN(new_n418));
  AOI22_X1  g232(.A1(new_n414), .A2(new_n327), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  OR2_X1    g233(.A1(new_n417), .A2(new_n418), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n413), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n408), .ZN(new_n422));
  AND2_X1   g236(.A1(new_n422), .A2(KEYINPUT86), .ZN(new_n423));
  OAI21_X1  g237(.A(KEYINPUT7), .B1(new_n422), .B2(KEYINPUT86), .ZN(new_n424));
  OR3_X1    g238(.A1(new_n406), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n404), .A2(KEYINPUT85), .A3(new_n405), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n422), .A2(KEYINPUT7), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n426), .B(new_n427), .C1(KEYINPUT85), .C2(new_n405), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n425), .A2(new_n399), .A3(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n411), .B1(new_n421), .B2(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n362), .B1(new_n410), .B2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n421), .ZN(new_n432));
  AND3_X1   g246(.A1(new_n425), .A2(new_n399), .A3(new_n428), .ZN(new_n433));
  AOI21_X1  g247(.A(G902), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n400), .A2(new_n402), .A3(new_n409), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n434), .A2(new_n361), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n360), .B1(new_n431), .B2(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n356), .A2(new_n358), .A3(new_n437), .ZN(new_n438));
  XNOR2_X1  g252(.A(G113), .B(G122), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n439), .B(new_n268), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n217), .A2(new_n218), .A3(KEYINPUT19), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(KEYINPUT90), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT90), .ZN(new_n444));
  INV_X1    g258(.A(new_n229), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n444), .B1(new_n445), .B2(KEYINPUT19), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n443), .B1(new_n442), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(new_n224), .ZN(new_n448));
  INV_X1    g262(.A(G237), .ZN(new_n449));
  AND4_X1   g263(.A1(G143), .A2(new_n449), .A3(new_n194), .A4(G214), .ZN(new_n450));
  NOR2_X1   g264(.A1(G237), .A2(G953), .ZN(new_n451));
  AOI21_X1  g265(.A(G143), .B1(new_n451), .B2(G214), .ZN(new_n452));
  OAI21_X1  g266(.A(G131), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n449), .A2(new_n194), .A3(G214), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(new_n255), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n451), .A2(G143), .A3(G214), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n455), .A2(new_n306), .A3(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n232), .B1(new_n453), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n448), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n217), .A2(new_n218), .A3(G146), .ZN(new_n460));
  AOI21_X1  g274(.A(KEYINPUT88), .B1(new_n229), .B2(new_n224), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AND2_X1   g276(.A1(KEYINPUT87), .A2(KEYINPUT18), .ZN(new_n463));
  OAI211_X1 g277(.A(G131), .B(new_n463), .C1(new_n450), .C2(new_n452), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(G131), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n455), .A2(new_n456), .A3(new_n465), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n217), .A2(new_n218), .A3(KEYINPUT88), .A4(G146), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n462), .A2(new_n464), .A3(new_n466), .A4(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT89), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n306), .B1(new_n455), .B2(new_n456), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n450), .A2(new_n452), .ZN(new_n472));
  AOI22_X1  g286(.A1(new_n471), .A2(new_n463), .B1(new_n472), .B2(new_n465), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n473), .A2(KEYINPUT89), .A3(new_n462), .A4(new_n467), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n470), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n440), .B1(new_n459), .B2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT17), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n453), .A2(new_n477), .A3(new_n457), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n471), .A2(KEYINPUT17), .ZN(new_n479));
  AND2_X1   g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n236), .A2(new_n232), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n440), .B(KEYINPUT91), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n475), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(KEYINPUT92), .ZN(new_n485));
  AOI22_X1  g299(.A1(new_n470), .A2(new_n474), .B1(new_n480), .B2(new_n481), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT92), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n486), .A2(new_n487), .A3(new_n483), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n476), .B1(new_n485), .B2(new_n488), .ZN(new_n489));
  NOR2_X1   g303(.A1(G475), .A2(G902), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(KEYINPUT20), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n459), .A2(new_n475), .ZN(new_n493));
  INV_X1    g307(.A(new_n440), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AND4_X1   g309(.A1(new_n487), .A2(new_n475), .A3(new_n482), .A4(new_n483), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n487), .B1(new_n486), .B2(new_n483), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT20), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n498), .A2(new_n499), .A3(new_n490), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n492), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(G478), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n502), .A2(KEYINPUT15), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(G122), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(G116), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n364), .A2(G122), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(KEYINPUT93), .ZN(new_n509));
  XNOR2_X1  g323(.A(G116), .B(G122), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT93), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(new_n271), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n364), .A2(KEYINPUT14), .A3(G122), .ZN(new_n515));
  OAI211_X1 g329(.A(G107), .B(new_n515), .C1(new_n508), .C2(KEYINPUT14), .ZN(new_n516));
  OR3_X1    g330(.A1(new_n205), .A2(KEYINPUT94), .A3(G143), .ZN(new_n517));
  OAI21_X1  g331(.A(KEYINPUT94), .B1(new_n205), .B2(G143), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n205), .A2(G143), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n519), .A2(new_n298), .A3(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n298), .B1(new_n519), .B2(new_n520), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n514), .B(new_n516), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n513), .A2(new_n271), .ZN(new_n525));
  AOI21_X1  g339(.A(G107), .B1(new_n509), .B2(new_n512), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n521), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT13), .ZN(new_n528));
  AOI22_X1  g342(.A1(new_n519), .A2(new_n528), .B1(new_n205), .B2(G143), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n517), .A2(KEYINPUT13), .A3(new_n518), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n298), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n524), .B1(new_n527), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(G217), .ZN(new_n533));
  NOR3_X1   g347(.A1(new_n357), .A2(new_n533), .A3(G953), .ZN(new_n534));
  XOR2_X1   g348(.A(new_n532), .B(new_n534), .Z(new_n535));
  AOI21_X1  g349(.A(new_n504), .B1(new_n535), .B2(new_n245), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n532), .B(new_n534), .ZN(new_n537));
  NOR3_X1   g351(.A1(new_n537), .A2(new_n187), .A3(new_n503), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(G234), .A2(G237), .ZN(new_n540));
  AND3_X1   g354(.A1(new_n187), .A2(G953), .A3(new_n540), .ZN(new_n541));
  XNOR2_X1  g355(.A(KEYINPUT21), .B(G898), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  XNOR2_X1  g357(.A(KEYINPUT95), .B(G952), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n544), .A2(G953), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(new_n540), .ZN(new_n546));
  AND2_X1   g360(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n486), .A2(new_n440), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n549), .B1(new_n485), .B2(new_n488), .ZN(new_n550));
  OAI21_X1  g364(.A(G475), .B1(new_n550), .B2(G902), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n501), .A2(new_n539), .A3(new_n548), .A4(new_n551), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n438), .A2(new_n552), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n294), .B1(new_n305), .B2(new_n312), .ZN(new_n554));
  AOI22_X1  g368(.A1(new_n368), .A2(new_n376), .B1(new_n366), .B2(new_n367), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n316), .A2(new_n266), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n298), .A2(G137), .ZN(new_n557));
  OAI21_X1  g371(.A(G131), .B1(new_n557), .B2(new_n307), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n556), .A2(new_n333), .A3(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n554), .A2(new_n555), .A3(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  AND3_X1   g375(.A1(new_n556), .A2(new_n333), .A3(new_n558), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n403), .B1(new_n334), .B2(new_n333), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n393), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(KEYINPUT69), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n554), .A2(new_n559), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT69), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n566), .A2(new_n567), .A3(new_n393), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n561), .B1(new_n565), .B2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT28), .ZN(new_n570));
  OAI21_X1  g384(.A(KEYINPUT70), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n567), .B1(new_n566), .B2(new_n393), .ZN(new_n572));
  AOI211_X1 g386(.A(KEYINPUT69), .B(new_n555), .C1(new_n554), .C2(new_n559), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n560), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT70), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n574), .A2(new_n575), .A3(KEYINPUT28), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n451), .A2(G210), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n577), .B(KEYINPUT27), .ZN(new_n578));
  XNOR2_X1  g392(.A(KEYINPUT26), .B(G101), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n578), .B(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n581), .B1(new_n560), .B2(new_n570), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n571), .A2(new_n576), .A3(new_n582), .ZN(new_n583));
  NOR3_X1   g397(.A1(new_n562), .A2(new_n563), .A3(KEYINPUT30), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT30), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n585), .B1(new_n554), .B2(new_n559), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n393), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(new_n560), .ZN(new_n588));
  AOI21_X1  g402(.A(KEYINPUT29), .B1(new_n588), .B2(new_n581), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n583), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(KEYINPUT71), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT71), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n583), .A2(new_n592), .A3(new_n589), .ZN(new_n593));
  AND2_X1   g407(.A1(new_n564), .A2(new_n560), .ZN(new_n594));
  OR2_X1    g408(.A1(new_n594), .A2(new_n570), .ZN(new_n595));
  AND2_X1   g409(.A1(new_n582), .A2(KEYINPUT29), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n187), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n591), .A2(new_n593), .A3(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n598), .A2(KEYINPUT73), .A3(G472), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n560), .A2(new_n570), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n571), .A2(new_n576), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(new_n581), .ZN(new_n602));
  XNOR2_X1  g416(.A(KEYINPUT67), .B(KEYINPUT31), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n587), .A2(new_n560), .A3(new_n580), .A4(new_n603), .ZN(new_n604));
  OAI21_X1  g418(.A(KEYINPUT30), .B1(new_n562), .B2(new_n563), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n554), .A2(new_n585), .A3(new_n559), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n555), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NOR3_X1   g421(.A1(new_n607), .A2(new_n561), .A3(new_n581), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT31), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n604), .B(KEYINPUT68), .C1(new_n608), .C2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT68), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n608), .A2(new_n611), .A3(new_n603), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n602), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT32), .ZN(new_n615));
  NOR2_X1   g429(.A1(G472), .A2(G902), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  AOI22_X1  g431(.A1(new_n601), .A2(new_n581), .B1(new_n610), .B2(new_n612), .ZN(new_n618));
  INV_X1    g432(.A(new_n616), .ZN(new_n619));
  OAI21_X1  g433(.A(KEYINPUT32), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n599), .A2(new_n621), .ZN(new_n622));
  AOI21_X1  g436(.A(KEYINPUT73), .B1(new_n598), .B2(G472), .ZN(new_n623));
  OAI211_X1 g437(.A(new_n254), .B(new_n553), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(KEYINPUT96), .B(G101), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(G3));
  INV_X1    g440(.A(KEYINPUT33), .ZN(new_n627));
  INV_X1    g441(.A(new_n532), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n627), .B1(new_n628), .B2(new_n534), .ZN(new_n629));
  XOR2_X1   g443(.A(new_n534), .B(KEYINPUT97), .Z(new_n630));
  AOI21_X1  g444(.A(KEYINPUT98), .B1(new_n532), .B2(new_n630), .ZN(new_n631));
  AND3_X1   g445(.A1(new_n532), .A2(KEYINPUT98), .A3(new_n630), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n629), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(KEYINPUT99), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n535), .A2(new_n627), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT99), .ZN(new_n636));
  OAI211_X1 g450(.A(new_n629), .B(new_n636), .C1(new_n631), .C2(new_n632), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n187), .A2(new_n502), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n634), .A2(new_n635), .A3(new_n637), .A4(new_n638), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n502), .B1(new_n537), .B2(new_n187), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NOR3_X1   g455(.A1(new_n489), .A2(KEYINPUT20), .A3(new_n491), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n499), .B1(new_n498), .B2(new_n490), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n551), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n437), .A2(new_n548), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT100), .ZN(new_n647));
  NOR3_X1   g461(.A1(new_n645), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  AOI22_X1  g462(.A1(new_n501), .A2(new_n551), .B1(new_n639), .B2(new_n640), .ZN(new_n649));
  NOR3_X1   g463(.A1(new_n410), .A2(new_n362), .A3(new_n430), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n361), .B1(new_n434), .B2(new_n435), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n359), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n652), .A2(new_n547), .ZN(new_n653));
  AOI21_X1  g467(.A(KEYINPUT100), .B1(new_n649), .B2(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n648), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n187), .B1(new_n602), .B2(new_n613), .ZN(new_n656));
  INV_X1    g470(.A(G472), .ZN(new_n657));
  OAI22_X1  g471(.A1(new_n656), .A2(new_n657), .B1(new_n619), .B2(new_n618), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n356), .A2(new_n254), .A3(new_n358), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n655), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT34), .B(G104), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G6));
  NOR3_X1   g477(.A1(new_n658), .A2(new_n659), .A3(new_n646), .ZN(new_n664));
  INV_X1    g478(.A(new_n539), .ZN(new_n665));
  INV_X1    g479(.A(new_n644), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n664), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT35), .B(G107), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G9));
  OAI22_X1  g483(.A1(new_n226), .A2(new_n233), .B1(new_n240), .B2(KEYINPUT36), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT36), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n237), .A2(new_n238), .A3(new_n201), .A4(new_n671), .ZN(new_n672));
  AND3_X1   g486(.A1(new_n670), .A2(new_n672), .A3(new_n252), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  OAI211_X1 g488(.A(new_n243), .B(new_n245), .C1(new_n246), .C2(new_n247), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n190), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n243), .B1(new_n251), .B2(new_n245), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n674), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(KEYINPUT101), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT101), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n250), .A2(new_n680), .A3(new_n674), .ZN(new_n681));
  AND3_X1   g495(.A1(new_n679), .A2(new_n681), .A3(KEYINPUT102), .ZN(new_n682));
  AOI21_X1  g496(.A(KEYINPUT102), .B1(new_n679), .B2(new_n681), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n684), .A2(new_n438), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n657), .B1(new_n614), .B2(new_n245), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n618), .A2(new_n619), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n686), .A2(new_n552), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  XOR2_X1   g503(.A(KEYINPUT37), .B(G110), .Z(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G12));
  INV_X1    g505(.A(KEYINPUT73), .ZN(new_n692));
  AND3_X1   g506(.A1(new_n583), .A2(new_n592), .A3(new_n589), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n592), .B1(new_n583), .B2(new_n589), .ZN(new_n694));
  INV_X1    g508(.A(new_n597), .ZN(new_n695));
  NOR3_X1   g509(.A1(new_n693), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n692), .B1(new_n696), .B2(new_n657), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n697), .A2(new_n621), .A3(new_n599), .ZN(new_n698));
  INV_X1    g512(.A(G900), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n541), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(new_n546), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n665), .A2(new_n501), .A3(new_n551), .A4(new_n701), .ZN(new_n702));
  NOR3_X1   g516(.A1(new_n684), .A2(new_n438), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n698), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G128), .ZN(G30));
  NOR2_X1   g519(.A1(new_n650), .A2(new_n651), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(KEYINPUT38), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n539), .B1(new_n501), .B2(new_n551), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n679), .A2(new_n681), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n710), .A2(new_n360), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n708), .A2(new_n709), .A3(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(new_n358), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n346), .A2(KEYINPUT81), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n354), .A2(new_n348), .A3(new_n342), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n713), .B1(new_n716), .B2(new_n341), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n701), .B(KEYINPUT39), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n712), .B1(KEYINPUT40), .B2(new_n719), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n720), .B1(KEYINPUT40), .B2(new_n719), .ZN(new_n721));
  INV_X1    g535(.A(new_n588), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n722), .A2(new_n581), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  AOI21_X1  g538(.A(G902), .B1(new_n594), .B2(new_n581), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n657), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n726), .B1(new_n617), .B2(new_n620), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n721), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(KEYINPUT103), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G143), .ZN(G45));
  NAND3_X1  g544(.A1(new_n641), .A2(new_n644), .A3(new_n701), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n698), .A2(new_n685), .A3(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G146), .ZN(G48));
  NAND2_X1  g548(.A1(new_n352), .A2(new_n353), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n342), .B1(new_n735), .B2(new_n245), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  OAI211_X1 g551(.A(new_n358), .B(new_n737), .C1(new_n347), .C2(new_n355), .ZN(new_n738));
  INV_X1    g552(.A(new_n254), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n698), .A2(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(new_n655), .ZN(new_n743));
  XNOR2_X1  g557(.A(KEYINPUT41), .B(G113), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n743), .B(new_n744), .ZN(G15));
  NAND2_X1  g559(.A1(new_n666), .A2(new_n665), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n746), .A2(new_n646), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n742), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G116), .ZN(G18));
  NOR2_X1   g563(.A1(new_n738), .A2(new_n652), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT102), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n680), .B1(new_n250), .B2(new_n674), .ZN(new_n752));
  AOI211_X1 g566(.A(KEYINPUT101), .B(new_n673), .C1(new_n244), .C2(new_n249), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n751), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n679), .A2(new_n681), .A3(KEYINPUT102), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(new_n552), .ZN(new_n757));
  AND3_X1   g571(.A1(new_n750), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n758), .B1(new_n622), .B2(new_n623), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(KEYINPUT104), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT104), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n698), .A2(new_n761), .A3(new_n758), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G119), .ZN(G21));
  NOR2_X1   g578(.A1(new_n604), .A2(KEYINPUT68), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n611), .B1(new_n608), .B2(new_n603), .ZN(new_n766));
  OAI21_X1  g580(.A(KEYINPUT31), .B1(new_n588), .B2(new_n581), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n765), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n580), .B1(new_n595), .B2(new_n600), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n616), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  XOR2_X1   g584(.A(KEYINPUT105), .B(G472), .Z(new_n771));
  OAI211_X1 g585(.A(new_n770), .B(new_n254), .C1(new_n656), .C2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n644), .A2(new_n548), .A3(new_n665), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n437), .A2(new_n716), .A3(new_n358), .A4(new_n737), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n773), .A2(new_n776), .A3(KEYINPUT106), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT106), .ZN(new_n778));
  AOI211_X1 g592(.A(new_n713), .B(new_n736), .C1(new_n714), .C2(new_n715), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n779), .A2(new_n709), .A3(new_n437), .A4(new_n548), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n778), .B1(new_n780), .B2(new_n772), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n777), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G122), .ZN(G24));
  OAI211_X1 g597(.A(new_n710), .B(new_n770), .C1(new_n656), .C2(new_n771), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n784), .A2(new_n731), .A3(new_n775), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(new_n215), .ZN(G27));
  INV_X1    g600(.A(KEYINPUT108), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n787), .A2(KEYINPUT42), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n254), .B1(new_n622), .B2(new_n623), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT107), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n706), .A2(new_n790), .A3(new_n359), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n431), .A2(new_n436), .A3(new_n359), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(KEYINPUT107), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n717), .A2(new_n791), .A3(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n795), .A2(new_n649), .A3(new_n701), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n788), .B1(new_n789), .B2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(new_n701), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n794), .A2(new_n645), .A3(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(new_n788), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n799), .A2(new_n698), .A3(new_n254), .A4(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n797), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(G131), .ZN(G33));
  AND2_X1   g617(.A1(new_n599), .A2(new_n621), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n739), .B1(new_n804), .B2(new_n697), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n702), .A2(KEYINPUT109), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n702), .A2(KEYINPUT109), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n806), .A2(new_n807), .A3(new_n794), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n805), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(G134), .ZN(G36));
  OR2_X1    g624(.A1(new_n340), .A2(KEYINPUT45), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n340), .A2(KEYINPUT45), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n811), .A2(G469), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(G469), .A2(G902), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT46), .ZN(new_n816));
  AOI22_X1  g630(.A1(new_n815), .A2(new_n816), .B1(new_n715), .B2(new_n714), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n817), .B1(new_n816), .B2(new_n815), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n818), .A2(new_n358), .A3(new_n718), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n791), .A2(new_n793), .ZN(new_n820));
  INV_X1    g634(.A(new_n820), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n666), .A2(new_n641), .ZN(new_n823));
  NAND2_X1  g637(.A1(KEYINPUT110), .A2(KEYINPUT43), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  XOR2_X1   g639(.A(KEYINPUT110), .B(KEYINPUT43), .Z(new_n826));
  OAI21_X1  g640(.A(new_n825), .B1(new_n823), .B2(new_n826), .ZN(new_n827));
  AND2_X1   g641(.A1(new_n658), .A2(new_n710), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT44), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n827), .A2(KEYINPUT44), .A3(new_n828), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n822), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  XOR2_X1   g647(.A(KEYINPUT111), .B(G137), .Z(new_n834));
  XNOR2_X1  g648(.A(new_n833), .B(new_n834), .ZN(G39));
  NAND2_X1  g649(.A1(new_n818), .A2(new_n358), .ZN(new_n836));
  XOR2_X1   g650(.A(new_n836), .B(KEYINPUT47), .Z(new_n837));
  NOR2_X1   g651(.A1(new_n622), .A2(new_n623), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n821), .A2(new_n254), .A3(new_n731), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n837), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n840), .B(KEYINPUT112), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n841), .B(G140), .ZN(G42));
  NAND2_X1  g656(.A1(new_n716), .A2(new_n737), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n843), .A2(new_n358), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n837), .A2(new_n844), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n827), .A2(new_n540), .A3(new_n545), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(new_n773), .ZN(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(new_n820), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n845), .B1(KEYINPUT118), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n850), .B1(KEYINPUT118), .B2(new_n849), .ZN(new_n851));
  NOR4_X1   g665(.A1(new_n847), .A2(new_n359), .A3(new_n708), .A4(new_n738), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n852), .B(KEYINPUT50), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n846), .A2(new_n779), .A3(new_n820), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n854), .A2(new_n784), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n739), .A2(new_n546), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n727), .A2(new_n779), .A3(new_n820), .A4(new_n856), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n857), .A2(new_n644), .A3(new_n641), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n851), .A2(new_n853), .A3(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT51), .ZN(new_n861));
  OR2_X1    g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n860), .A2(new_n861), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n545), .B1(new_n857), .B2(new_n645), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n854), .A2(new_n789), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n865), .B(KEYINPUT48), .ZN(new_n866));
  AOI211_X1 g680(.A(new_n864), .B(new_n866), .C1(new_n750), .C2(new_n848), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n862), .A2(new_n863), .A3(new_n867), .ZN(new_n868));
  OAI211_X1 g682(.A(new_n698), .B(new_n740), .C1(new_n655), .C2(new_n747), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n746), .A2(new_n645), .ZN(new_n870));
  AOI22_X1  g684(.A1(new_n664), .A2(new_n870), .B1(new_n685), .B2(new_n688), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n869), .A2(new_n624), .A3(new_n782), .A4(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(new_n762), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n761), .B1(new_n698), .B2(new_n758), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n785), .B1(new_n698), .B2(new_n703), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n678), .A2(new_n798), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n709), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n879), .A2(new_n438), .ZN(new_n880));
  INV_X1    g694(.A(new_n726), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n615), .B1(new_n614), .B2(new_n616), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n618), .A2(KEYINPUT32), .A3(new_n619), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n881), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n880), .A2(new_n884), .A3(KEYINPUT114), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT114), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n717), .A2(new_n709), .A3(new_n437), .A4(new_n878), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n886), .B1(new_n727), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n877), .A2(new_n889), .A3(new_n733), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT52), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n877), .A2(new_n889), .A3(new_n733), .A4(KEYINPUT52), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n501), .A2(new_n539), .A3(new_n551), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n895), .B1(new_n755), .B2(new_n754), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n820), .A2(new_n896), .A3(new_n717), .A4(new_n701), .ZN(new_n897));
  OAI21_X1  g711(.A(KEYINPUT113), .B1(new_n838), .B2(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT113), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n794), .A2(new_n798), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n698), .A2(new_n899), .A3(new_n900), .A4(new_n896), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n784), .A2(new_n731), .ZN(new_n903));
  AOI22_X1  g717(.A1(new_n805), .A2(new_n808), .B1(new_n903), .B2(new_n795), .ZN(new_n904));
  AND2_X1   g718(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n876), .A2(new_n894), .A3(new_n802), .A4(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT53), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT115), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n894), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n892), .A2(KEYINPUT115), .A3(new_n893), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n802), .A2(new_n902), .A3(new_n904), .ZN(new_n913));
  AND3_X1   g727(.A1(new_n871), .A2(new_n782), .A3(new_n624), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n914), .A2(new_n763), .A3(new_n869), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n912), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n908), .B1(new_n917), .B2(new_n907), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT54), .ZN(new_n919));
  OR2_X1    g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AND3_X1   g734(.A1(new_n892), .A2(KEYINPUT115), .A3(new_n893), .ZN(new_n921));
  AOI21_X1  g735(.A(KEYINPUT115), .B1(new_n892), .B2(new_n893), .ZN(new_n922));
  OAI211_X1 g736(.A(new_n916), .B(KEYINPUT53), .C1(new_n921), .C2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT117), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n912), .A2(KEYINPUT117), .A3(KEYINPUT53), .A4(new_n916), .ZN(new_n926));
  AND3_X1   g740(.A1(new_n906), .A2(KEYINPUT116), .A3(new_n907), .ZN(new_n927));
  AOI21_X1  g741(.A(KEYINPUT116), .B1(new_n906), .B2(new_n907), .ZN(new_n928));
  OAI211_X1 g742(.A(new_n925), .B(new_n926), .C1(new_n927), .C2(new_n928), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n920), .B1(KEYINPUT54), .B2(new_n929), .ZN(new_n930));
  OAI22_X1  g744(.A1(new_n868), .A2(new_n930), .B1(G952), .B2(G953), .ZN(new_n931));
  NOR4_X1   g745(.A1(new_n708), .A2(new_n739), .A3(new_n713), .A4(new_n360), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n823), .B1(KEYINPUT49), .B2(new_n843), .ZN(new_n933));
  OAI211_X1 g747(.A(new_n932), .B(new_n933), .C1(KEYINPUT49), .C2(new_n843), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n931), .B1(new_n884), .B2(new_n934), .ZN(G75));
  NAND3_X1  g749(.A1(new_n929), .A2(new_n187), .A3(new_n362), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n400), .A2(new_n402), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(new_n409), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n938), .B(KEYINPUT55), .Z(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(KEYINPUT121), .ZN(new_n940));
  OR2_X1    g754(.A1(new_n939), .A2(KEYINPUT121), .ZN(new_n941));
  XOR2_X1   g755(.A(KEYINPUT120), .B(KEYINPUT56), .Z(new_n942));
  AND4_X1   g756(.A1(new_n936), .A2(new_n940), .A3(new_n941), .A4(new_n942), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n194), .A2(G952), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(KEYINPUT122), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(KEYINPUT56), .B1(new_n936), .B2(KEYINPUT119), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n947), .B1(KEYINPUT119), .B2(new_n936), .ZN(new_n948));
  AOI211_X1 g762(.A(new_n943), .B(new_n946), .C1(new_n948), .C2(new_n939), .ZN(G51));
  XNOR2_X1  g763(.A(new_n929), .B(KEYINPUT54), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n814), .B(KEYINPUT57), .Z(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(new_n735), .ZN(new_n953));
  INV_X1    g767(.A(new_n813), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n929), .A2(new_n187), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n944), .B1(new_n953), .B2(new_n955), .ZN(G54));
  NAND4_X1  g770(.A1(new_n929), .A2(KEYINPUT58), .A3(G475), .A4(new_n187), .ZN(new_n957));
  AND2_X1   g771(.A1(new_n957), .A2(new_n489), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n957), .A2(new_n489), .ZN(new_n959));
  NOR3_X1   g773(.A1(new_n958), .A2(new_n959), .A3(new_n944), .ZN(G60));
  AND3_X1   g774(.A1(new_n634), .A2(new_n635), .A3(new_n637), .ZN(new_n961));
  NAND2_X1  g775(.A1(G478), .A2(G902), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n962), .B(KEYINPUT59), .ZN(new_n963));
  AND3_X1   g777(.A1(new_n950), .A2(new_n961), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n961), .B1(new_n930), .B2(new_n963), .ZN(new_n965));
  NOR3_X1   g779(.A1(new_n964), .A2(new_n965), .A3(new_n946), .ZN(G63));
  AND2_X1   g780(.A1(new_n670), .A2(new_n672), .ZN(new_n967));
  NAND2_X1  g781(.A1(G217), .A2(G902), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n968), .B(KEYINPUT60), .Z(new_n969));
  AND3_X1   g783(.A1(new_n929), .A2(KEYINPUT123), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(KEYINPUT123), .B1(new_n929), .B2(new_n969), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n967), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n929), .A2(new_n969), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT123), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(new_n251), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n929), .A2(KEYINPUT123), .A3(new_n969), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n975), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n972), .A2(new_n978), .A3(new_n945), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT61), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n972), .A2(new_n978), .A3(KEYINPUT61), .A4(new_n945), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n981), .A2(new_n982), .ZN(G66));
  OAI21_X1  g797(.A(G953), .B1(new_n542), .B2(new_n407), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n984), .B1(new_n876), .B2(G953), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n937), .B1(G898), .B2(new_n194), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n986), .B(KEYINPUT124), .Z(new_n987));
  XNOR2_X1  g801(.A(new_n985), .B(new_n987), .ZN(G69));
  NAND2_X1  g802(.A1(new_n605), .A2(new_n606), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n989), .B(new_n447), .Z(new_n990));
  INV_X1    g804(.A(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(new_n729), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n877), .A2(new_n733), .ZN(new_n993));
  OR3_X1    g807(.A1(new_n992), .A2(KEYINPUT62), .A3(new_n993), .ZN(new_n994));
  OAI21_X1  g808(.A(KEYINPUT62), .B1(new_n992), .B2(new_n993), .ZN(new_n995));
  AND2_X1   g809(.A1(new_n841), .A2(new_n833), .ZN(new_n996));
  INV_X1    g810(.A(new_n870), .ZN(new_n997));
  NOR4_X1   g811(.A1(new_n789), .A2(new_n821), .A3(new_n719), .A4(new_n997), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n998), .B(KEYINPUT125), .ZN(new_n999));
  NAND4_X1  g813(.A1(new_n994), .A2(new_n995), .A3(new_n996), .A4(new_n999), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n991), .B1(new_n1000), .B2(new_n194), .ZN(new_n1001));
  INV_X1    g815(.A(new_n808), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n709), .A2(new_n437), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n1002), .B1(new_n819), .B2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n993), .B1(new_n1004), .B2(new_n805), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n996), .A2(new_n802), .A3(new_n1005), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n1006), .A2(G953), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n990), .B1(G900), .B2(G953), .ZN(new_n1008));
  INV_X1    g822(.A(new_n1008), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n194), .B1(G227), .B2(G900), .ZN(new_n1011));
  OR3_X1    g825(.A1(new_n1001), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n1011), .B1(new_n1001), .B2(new_n1010), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1012), .A2(new_n1013), .ZN(G72));
  XNOR2_X1  g828(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1015));
  NOR2_X1   g829(.A1(new_n657), .A2(new_n411), .ZN(new_n1016));
  XNOR2_X1  g830(.A(new_n1015), .B(new_n1016), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n1017), .B1(new_n1000), .B2(new_n915), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1018), .A2(new_n723), .ZN(new_n1019));
  NOR2_X1   g833(.A1(new_n588), .A2(new_n580), .ZN(new_n1020));
  INV_X1    g834(.A(new_n1020), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n724), .A2(new_n1021), .A3(new_n1017), .ZN(new_n1022));
  XNOR2_X1  g836(.A(new_n1022), .B(KEYINPUT127), .ZN(new_n1023));
  OR2_X1    g837(.A1(new_n918), .A2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g838(.A(new_n1017), .B1(new_n1006), .B2(new_n915), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n944), .B1(new_n1025), .B2(new_n1020), .ZN(new_n1026));
  AND3_X1   g840(.A1(new_n1019), .A2(new_n1024), .A3(new_n1026), .ZN(G57));
endmodule


