//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 0 0 0 1 0 0 1 1 0 0 0 1 0 1 1 0 1 1 0 1 0 1 0 0 1 0 1 1 0 0 1 0 1 0 1 1 1 1 1 1 1 0 1 0 1 1 0 1 0 0 1 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n728, new_n729,
    new_n731, new_n732, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n818, new_n819, new_n821,
    new_n822, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n881,
    new_n882, new_n884, new_n885, new_n886, new_n887, new_n888, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n902, new_n903, new_n904, new_n906,
    new_n907, new_n908, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n929, new_n930,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n939,
    new_n940;
  XNOR2_X1  g000(.A(G113gat), .B(G120gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT69), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G127gat), .B(G134gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(KEYINPUT70), .B(KEYINPUT1), .ZN(new_n206));
  INV_X1    g005(.A(G120gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n207), .A2(KEYINPUT69), .A3(G113gat), .ZN(new_n208));
  NAND4_X1  g007(.A1(new_n204), .A2(new_n205), .A3(new_n206), .A4(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(new_n205), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n210), .B1(KEYINPUT1), .B2(new_n202), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G148gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(G141gat), .ZN(new_n214));
  INV_X1    g013(.A(G141gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(G148gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n214), .A2(new_n216), .A3(KEYINPUT72), .ZN(new_n217));
  XNOR2_X1  g016(.A(G155gat), .B(G162gat), .ZN(new_n218));
  INV_X1    g017(.A(G155gat), .ZN(new_n219));
  INV_X1    g018(.A(G162gat), .ZN(new_n220));
  OAI21_X1  g019(.A(KEYINPUT2), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT72), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n222), .A2(new_n215), .A3(G148gat), .ZN(new_n223));
  NAND4_X1  g022(.A1(new_n217), .A2(new_n218), .A3(new_n221), .A4(new_n223), .ZN(new_n224));
  AND2_X1   g023(.A1(G155gat), .A2(G162gat), .ZN(new_n225));
  NOR2_X1   g024(.A1(G155gat), .A2(G162gat), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(G141gat), .B(G148gat), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n227), .B1(new_n228), .B2(KEYINPUT2), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n224), .A2(new_n229), .ZN(new_n230));
  OR3_X1    g029(.A1(new_n212), .A2(KEYINPUT4), .A3(new_n230), .ZN(new_n231));
  OAI21_X1  g030(.A(KEYINPUT4), .B1(new_n212), .B2(new_n230), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT74), .ZN(new_n234));
  AND3_X1   g033(.A1(new_n224), .A2(KEYINPUT73), .A3(new_n229), .ZN(new_n235));
  AOI21_X1  g034(.A(KEYINPUT73), .B1(new_n224), .B2(new_n229), .ZN(new_n236));
  OAI211_X1 g035(.A(new_n234), .B(KEYINPUT3), .C1(new_n235), .C2(new_n236), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n230), .A2(KEYINPUT3), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n237), .A2(new_n212), .A3(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT73), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n230), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n224), .A2(KEYINPUT73), .A3(new_n229), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n234), .B1(new_n244), .B2(KEYINPUT3), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n233), .B1(new_n240), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(G225gat), .A2(G233gat), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  OR2_X1    g048(.A1(new_n212), .A2(new_n230), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n235), .A2(new_n236), .ZN(new_n251));
  INV_X1    g050(.A(new_n212), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n250), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  OR2_X1    g052(.A1(new_n253), .A2(new_n248), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n249), .A2(KEYINPUT39), .A3(new_n254), .ZN(new_n255));
  XNOR2_X1  g054(.A(KEYINPUT79), .B(KEYINPUT39), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n246), .A2(new_n248), .A3(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(G1gat), .B(G29gat), .ZN(new_n258));
  INV_X1    g057(.A(G85gat), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n258), .B(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(KEYINPUT0), .B(G57gat), .ZN(new_n261));
  XOR2_X1   g060(.A(new_n260), .B(new_n261), .Z(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  AND3_X1   g062(.A1(new_n257), .A2(KEYINPUT80), .A3(new_n263), .ZN(new_n264));
  AOI21_X1  g063(.A(KEYINPUT80), .B1(new_n257), .B2(new_n263), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n255), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT81), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT40), .ZN(new_n268));
  AND3_X1   g067(.A1(new_n266), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n267), .B1(new_n266), .B2(new_n268), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(G197gat), .B(G204gat), .ZN(new_n272));
  INV_X1    g071(.A(G211gat), .ZN(new_n273));
  INV_X1    g072(.A(G218gat), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n272), .B1(KEYINPUT22), .B2(new_n275), .ZN(new_n276));
  XOR2_X1   g075(.A(G211gat), .B(G218gat), .Z(new_n277));
  XOR2_X1   g076(.A(new_n276), .B(new_n277), .Z(new_n278));
  NAND2_X1  g077(.A1(G226gat), .A2(G233gat), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(G169gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(KEYINPUT23), .ZN(new_n282));
  INV_X1    g081(.A(G176gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(KEYINPUT65), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT65), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(G176gat), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n282), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  NOR2_X1   g086(.A1(G169gat), .A2(G176gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(G169gat), .A2(G176gat), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n288), .B1(KEYINPUT23), .B2(new_n289), .ZN(new_n290));
  OAI21_X1  g089(.A(KEYINPUT66), .B1(new_n287), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(G183gat), .A2(G190gat), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT24), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NOR2_X1   g093(.A1(G183gat), .A2(G190gat), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n292), .A2(new_n293), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT64), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n292), .A2(KEYINPUT64), .A3(new_n293), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n296), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n289), .A2(KEYINPUT23), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n281), .A2(new_n283), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT66), .ZN(new_n305));
  XNOR2_X1  g104(.A(KEYINPUT65), .B(G176gat), .ZN(new_n306));
  OAI211_X1 g105(.A(new_n304), .B(new_n305), .C1(new_n306), .C2(new_n282), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n291), .A2(new_n301), .A3(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT25), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT67), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n308), .A2(KEYINPUT67), .A3(new_n309), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n296), .A2(new_n297), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n281), .A2(new_n283), .A3(KEYINPUT23), .ZN(new_n315));
  NAND4_X1  g114(.A1(new_n314), .A2(KEYINPUT25), .A3(new_n304), .A4(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n312), .A2(new_n313), .A3(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(KEYINPUT27), .B(G183gat), .ZN(new_n318));
  INV_X1    g117(.A(G190gat), .ZN(new_n319));
  AOI21_X1  g118(.A(KEYINPUT68), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  XOR2_X1   g119(.A(new_n320), .B(KEYINPUT28), .Z(new_n321));
  OR2_X1    g120(.A1(new_n303), .A2(KEYINPUT26), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n303), .A2(KEYINPUT26), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n322), .A2(new_n289), .A3(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n321), .A2(new_n324), .A3(new_n292), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n317), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT29), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n280), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n279), .B1(new_n317), .B2(new_n325), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n278), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n329), .ZN(new_n331));
  INV_X1    g130(.A(new_n278), .ZN(new_n332));
  AOI21_X1  g131(.A(KEYINPUT29), .B1(new_n317), .B2(new_n325), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n331), .B(new_n332), .C1(new_n280), .C2(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(G8gat), .B(G36gat), .ZN(new_n335));
  XNOR2_X1  g134(.A(G64gat), .B(G92gat), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n335), .B(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n330), .A2(new_n334), .A3(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT30), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n326), .A2(new_n327), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(new_n279), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n332), .B1(new_n343), .B2(new_n331), .ZN(new_n344));
  NOR3_X1   g143(.A1(new_n328), .A2(new_n278), .A3(new_n329), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n337), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND4_X1  g145(.A1(new_n330), .A2(new_n334), .A3(KEYINPUT30), .A4(new_n338), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n341), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT82), .ZN(new_n349));
  OAI211_X1 g148(.A(new_n247), .B(new_n233), .C1(new_n240), .C2(new_n245), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT5), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n351), .B1(new_n253), .B2(new_n248), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n350), .A2(new_n352), .A3(KEYINPUT75), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT3), .ZN(new_n354));
  OAI21_X1  g153(.A(KEYINPUT74), .B1(new_n251), .B2(new_n354), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n355), .A2(new_n237), .A3(new_n212), .A4(new_n239), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n356), .A2(new_n351), .A3(new_n247), .A4(new_n233), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n353), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(KEYINPUT75), .B1(new_n350), .B2(new_n352), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n349), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n350), .A2(new_n352), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT75), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND4_X1  g162(.A1(new_n363), .A2(KEYINPUT82), .A3(new_n357), .A4(new_n353), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n360), .A2(new_n262), .A3(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n255), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n257), .A2(new_n263), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT80), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n257), .A2(KEYINPUT80), .A3(new_n263), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n366), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(KEYINPUT40), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n271), .A2(new_n348), .A3(new_n365), .A4(new_n372), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n354), .B1(new_n278), .B2(KEYINPUT29), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(new_n244), .ZN(new_n375));
  INV_X1    g174(.A(G228gat), .ZN(new_n376));
  INV_X1    g175(.A(G233gat), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n278), .B1(new_n238), .B2(KEYINPUT29), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n375), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  XNOR2_X1  g180(.A(KEYINPUT76), .B(G22gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n374), .A2(new_n230), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n378), .B1(new_n383), .B2(new_n379), .ZN(new_n384));
  OR3_X1    g183(.A1(new_n381), .A2(new_n382), .A3(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT77), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n382), .B1(new_n381), .B2(new_n384), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  XNOR2_X1  g187(.A(G78gat), .B(G106gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(KEYINPUT31), .B(G50gat), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n389), .B(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n384), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(new_n380), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n394), .A2(KEYINPUT77), .A3(new_n382), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n388), .A2(new_n392), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n394), .A2(G22gat), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n397), .A2(new_n385), .A3(new_n391), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT37), .ZN(new_n400));
  AND3_X1   g199(.A1(new_n330), .A2(new_n334), .A3(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n400), .B1(new_n330), .B2(new_n334), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT38), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n403), .A2(new_n404), .A3(new_n337), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT83), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n403), .A2(KEYINPUT83), .A3(new_n404), .A4(new_n337), .ZN(new_n409));
  OAI211_X1 g208(.A(KEYINPUT6), .B(new_n262), .C1(new_n358), .C2(new_n359), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n358), .A2(new_n359), .ZN(new_n412));
  AOI21_X1  g211(.A(KEYINPUT6), .B1(new_n412), .B2(new_n263), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n411), .B1(new_n365), .B2(new_n413), .ZN(new_n414));
  OAI21_X1  g213(.A(KEYINPUT37), .B1(new_n344), .B2(new_n345), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n330), .A2(new_n334), .A3(new_n400), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n415), .A2(new_n337), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(KEYINPUT38), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n409), .A2(new_n414), .A3(new_n418), .A4(new_n339), .ZN(new_n419));
  OAI211_X1 g218(.A(new_n373), .B(new_n399), .C1(new_n408), .C2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT78), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT36), .ZN(new_n422));
  XOR2_X1   g221(.A(G71gat), .B(G99gat), .Z(new_n423));
  XNOR2_X1  g222(.A(G15gat), .B(G43gat), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n423), .B(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(G227gat), .A2(G233gat), .ZN(new_n426));
  AND3_X1   g225(.A1(new_n308), .A2(KEYINPUT67), .A3(new_n309), .ZN(new_n427));
  AOI21_X1  g226(.A(KEYINPUT67), .B1(new_n308), .B2(new_n309), .ZN(new_n428));
  INV_X1    g227(.A(new_n316), .ZN(new_n429));
  NOR3_X1   g228(.A1(new_n427), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n325), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n212), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n317), .A2(new_n252), .A3(new_n325), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n426), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n425), .B1(new_n434), .B2(KEYINPUT33), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n432), .A2(new_n426), .A3(new_n433), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT34), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(KEYINPUT71), .ZN(new_n438));
  AND2_X1   g237(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n435), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n436), .A2(new_n438), .ZN(new_n441));
  INV_X1    g240(.A(new_n426), .ZN(new_n442));
  AND3_X1   g241(.A1(new_n317), .A2(new_n252), .A3(new_n325), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n252), .B1(new_n317), .B2(new_n325), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n442), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT33), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n441), .B1(new_n447), .B2(new_n425), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n437), .A2(KEYINPUT71), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT32), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n449), .B1(new_n434), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n449), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n445), .A2(KEYINPUT32), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NOR3_X1   g253(.A1(new_n440), .A2(new_n448), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n435), .A2(new_n439), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n447), .A2(new_n441), .A3(new_n425), .ZN(new_n457));
  AOI22_X1  g256(.A1(new_n456), .A2(new_n457), .B1(new_n451), .B2(new_n453), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n422), .B1(new_n455), .B2(new_n458), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n454), .B1(new_n440), .B2(new_n448), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n456), .A2(new_n457), .A3(new_n451), .A4(new_n453), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n460), .A2(KEYINPUT36), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  AND3_X1   g262(.A1(new_n341), .A2(new_n346), .A3(new_n347), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n262), .B1(new_n358), .B2(new_n359), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT6), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n363), .A2(new_n263), .A3(new_n357), .A4(new_n353), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(new_n410), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n399), .B1(new_n464), .B2(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n421), .B1(new_n463), .B2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n399), .ZN(new_n472));
  INV_X1    g271(.A(new_n469), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n472), .B1(new_n473), .B2(new_n348), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n474), .A2(KEYINPUT78), .A3(new_n462), .A4(new_n459), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n420), .A2(new_n471), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n477), .A2(new_n469), .A3(new_n464), .A4(new_n399), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(KEYINPUT35), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT85), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT84), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n482), .B1(new_n455), .B2(new_n458), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n460), .A2(KEYINPUT84), .A3(new_n461), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n414), .A2(KEYINPUT35), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n485), .A2(new_n464), .A3(new_n399), .A4(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n478), .A2(KEYINPUT85), .A3(KEYINPUT35), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n481), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n476), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT86), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n476), .A2(new_n489), .A3(KEYINPUT86), .ZN(new_n493));
  XNOR2_X1  g292(.A(G15gat), .B(G22gat), .ZN(new_n494));
  INV_X1    g293(.A(G1gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(KEYINPUT16), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n497), .B1(G1gat), .B2(new_n494), .ZN(new_n498));
  OR2_X1    g297(.A1(new_n498), .A2(G8gat), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(G8gat), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  OR2_X1    g300(.A1(G29gat), .A2(G36gat), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n502), .B(KEYINPUT14), .ZN(new_n503));
  XNOR2_X1  g302(.A(KEYINPUT88), .B(G29gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(G36gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  XOR2_X1   g305(.A(G43gat), .B(G50gat), .Z(new_n507));
  INV_X1    g306(.A(KEYINPUT15), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n505), .A2(KEYINPUT89), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n507), .A2(new_n508), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT89), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n504), .A2(new_n513), .A3(G36gat), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n511), .A2(new_n503), .A3(new_n512), .A4(new_n514), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n510), .B1(new_n515), .B2(new_n509), .ZN(new_n516));
  AND2_X1   g315(.A1(new_n501), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n516), .B(KEYINPUT17), .ZN(new_n518));
  AND2_X1   g317(.A1(new_n499), .A2(new_n500), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(G229gat), .A2(G233gat), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n521), .B(KEYINPUT90), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n520), .A2(KEYINPUT18), .A3(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n517), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT17), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n516), .B(new_n525), .ZN(new_n526));
  OAI211_X1 g325(.A(new_n522), .B(new_n524), .C1(new_n526), .C2(new_n501), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT18), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  XOR2_X1   g328(.A(new_n522), .B(KEYINPUT13), .Z(new_n530));
  NOR2_X1   g329(.A1(new_n501), .A2(new_n516), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n530), .B1(new_n517), .B2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT91), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  OAI211_X1 g333(.A(KEYINPUT91), .B(new_n530), .C1(new_n517), .C2(new_n531), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n523), .A2(new_n529), .A3(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(G113gat), .B(G141gat), .ZN(new_n538));
  INV_X1    g337(.A(G197gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n538), .B(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(KEYINPUT11), .B(G169gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n540), .B(new_n541), .ZN(new_n542));
  XOR2_X1   g341(.A(KEYINPUT87), .B(KEYINPUT12), .Z(new_n543));
  XNOR2_X1  g342(.A(new_n542), .B(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n537), .A2(new_n545), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n523), .A2(new_n529), .A3(new_n536), .A4(new_n544), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT92), .ZN(new_n548));
  AND2_X1   g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n547), .A2(new_n548), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n546), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n492), .A2(new_n493), .A3(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(G64gat), .ZN(new_n553));
  AND2_X1   g352(.A1(new_n553), .A2(G57gat), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n553), .A2(G57gat), .ZN(new_n555));
  AND2_X1   g354(.A1(G71gat), .A2(G78gat), .ZN(new_n556));
  OAI22_X1  g355(.A1(new_n554), .A2(new_n555), .B1(KEYINPUT9), .B2(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(G71gat), .B(G78gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n557), .B(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n501), .B1(KEYINPUT21), .B2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT94), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n560), .B(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n562), .B(new_n563), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n559), .A2(KEYINPUT21), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  OR2_X1    g365(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n564), .A2(new_n566), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  XOR2_X1   g368(.A(G127gat), .B(G155gat), .Z(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(KEYINPUT93), .ZN(new_n571));
  XOR2_X1   g370(.A(G183gat), .B(G211gat), .Z(new_n572));
  NAND2_X1  g371(.A1(G231gat), .A2(G233gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  XOR2_X1   g373(.A(new_n571), .B(new_n574), .Z(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n569), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n567), .A2(new_n568), .A3(new_n575), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(G99gat), .A2(G106gat), .ZN(new_n580));
  INV_X1    g379(.A(G92gat), .ZN(new_n581));
  AOI22_X1  g380(.A1(KEYINPUT8), .A2(new_n580), .B1(new_n259), .B2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT7), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n583), .B1(new_n259), .B2(new_n581), .ZN(new_n584));
  NAND3_X1  g383(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n582), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  XOR2_X1   g385(.A(G99gat), .B(G106gat), .Z(new_n587));
  OR2_X1    g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n586), .A2(new_n587), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n588), .A2(KEYINPUT96), .A3(new_n589), .ZN(new_n590));
  OR3_X1    g389(.A1(new_n586), .A2(KEYINPUT96), .A3(new_n587), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(new_n516), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT41), .ZN(new_n594));
  NAND2_X1  g393(.A1(G232gat), .A2(G233gat), .ZN(new_n595));
  OAI221_X1 g394(.A(new_n593), .B1(new_n594), .B2(new_n595), .C1(new_n526), .C2(new_n592), .ZN(new_n596));
  XOR2_X1   g395(.A(G190gat), .B(G218gat), .Z(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n596), .B(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n595), .A2(new_n594), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(new_n220), .ZN(new_n601));
  XNOR2_X1  g400(.A(KEYINPUT95), .B(G134gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  OR3_X1    g402(.A1(new_n599), .A2(KEYINPUT97), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n599), .A2(new_n603), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n596), .A2(new_n598), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(KEYINPUT97), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n604), .A2(new_n605), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n579), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n559), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n611), .A2(new_n590), .A3(new_n591), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n559), .A2(new_n588), .A3(new_n589), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(G230gat), .A2(G233gat), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  OR2_X1    g416(.A1(new_n617), .A2(KEYINPUT98), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(KEYINPUT98), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT10), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n612), .A2(new_n620), .A3(new_n613), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n592), .A2(KEYINPUT10), .A3(new_n559), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n616), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n618), .A2(new_n619), .A3(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(G120gat), .B(G148gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(G176gat), .B(G204gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  OR2_X1    g427(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n625), .A2(new_n628), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n610), .A2(new_n632), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n552), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(new_n473), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g435(.A1(new_n634), .A2(new_n348), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(G8gat), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(KEYINPUT42), .ZN(new_n639));
  XNOR2_X1  g438(.A(KEYINPUT99), .B(KEYINPUT16), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(G8gat), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n637), .A2(new_n641), .ZN(new_n642));
  MUX2_X1   g441(.A(new_n639), .B(KEYINPUT42), .S(new_n642), .Z(G1325gat));
  INV_X1    g442(.A(KEYINPUT100), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n463), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(KEYINPUT100), .B1(new_n459), .B2(new_n462), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  AND3_X1   g447(.A1(new_n634), .A2(G15gat), .A3(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(G15gat), .B1(new_n634), .B2(new_n485), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n649), .A2(new_n650), .ZN(G1326gat));
  NAND2_X1  g450(.A1(new_n634), .A2(new_n472), .ZN(new_n652));
  XNOR2_X1  g451(.A(KEYINPUT43), .B(G22gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(G1327gat));
  INV_X1    g453(.A(KEYINPUT44), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n608), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n492), .A2(new_n493), .A3(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n488), .ZN(new_n658));
  AOI21_X1  g457(.A(KEYINPUT85), .B1(new_n478), .B2(KEYINPUT35), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  OAI21_X1  g459(.A(KEYINPUT81), .B1(new_n371), .B2(KEYINPUT40), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n266), .A2(new_n267), .A3(new_n268), .ZN(new_n662));
  AND4_X1   g461(.A1(new_n365), .A2(new_n661), .A3(new_n372), .A4(new_n662), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n472), .B1(new_n663), .B2(new_n348), .ZN(new_n664));
  AND2_X1   g463(.A1(new_n414), .A2(new_n418), .ZN(new_n665));
  NAND4_X1  g464(.A1(new_n665), .A2(new_n339), .A3(new_n407), .A4(new_n409), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n470), .B1(new_n664), .B2(new_n666), .ZN(new_n667));
  AOI22_X1  g466(.A1(new_n660), .A2(new_n487), .B1(new_n667), .B2(new_n647), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n655), .B1(new_n668), .B2(new_n608), .ZN(new_n669));
  AND2_X1   g468(.A1(new_n657), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n551), .ZN(new_n671));
  NOR3_X1   g470(.A1(new_n579), .A2(new_n671), .A3(new_n631), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n504), .B1(new_n673), .B2(new_n469), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n579), .A2(new_n631), .ZN(new_n675));
  NAND4_X1  g474(.A1(new_n492), .A2(new_n493), .A3(new_n551), .A4(new_n675), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n676), .A2(new_n469), .A3(new_n608), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT45), .ZN(new_n678));
  INV_X1    g477(.A(new_n504), .ZN(new_n679));
  AND3_X1   g478(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n678), .B1(new_n677), .B2(new_n679), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n674), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(KEYINPUT101), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT101), .ZN(new_n684));
  OAI211_X1 g483(.A(new_n674), .B(new_n684), .C1(new_n681), .C2(new_n680), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n683), .A2(new_n685), .ZN(G1328gat));
  NOR2_X1   g485(.A1(new_n676), .A2(new_n608), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n464), .A2(G36gat), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  OR2_X1    g488(.A1(new_n689), .A2(KEYINPUT46), .ZN(new_n690));
  OAI21_X1  g489(.A(G36gat), .B1(new_n673), .B2(new_n464), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n689), .A2(KEYINPUT46), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n690), .A2(new_n691), .A3(new_n692), .ZN(G1329gat));
  OAI21_X1  g492(.A(G43gat), .B1(new_n673), .B2(new_n647), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT47), .ZN(new_n695));
  INV_X1    g494(.A(G43gat), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n687), .A2(new_n696), .A3(new_n485), .ZN(new_n697));
  AND3_X1   g496(.A1(new_n694), .A2(new_n695), .A3(new_n697), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n695), .B1(new_n694), .B2(new_n697), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n698), .A2(new_n699), .ZN(G1330gat));
  OAI21_X1  g499(.A(G50gat), .B1(new_n673), .B2(new_n399), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n687), .A2(KEYINPUT102), .ZN(new_n702));
  INV_X1    g501(.A(G50gat), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT102), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n704), .B1(new_n676), .B2(new_n608), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n702), .A2(new_n703), .A3(new_n472), .A4(new_n705), .ZN(new_n706));
  OR2_X1    g505(.A1(KEYINPUT103), .A2(KEYINPUT48), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n701), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(KEYINPUT103), .A2(KEYINPUT48), .ZN(new_n709));
  XOR2_X1   g508(.A(new_n709), .B(KEYINPUT104), .Z(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n701), .A2(new_n706), .A3(new_n710), .A4(new_n707), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(G1331gat));
  NOR2_X1   g513(.A1(new_n668), .A2(new_n551), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n609), .A2(new_n632), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(new_n473), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(G57gat), .ZN(G1332gat));
  INV_X1    g519(.A(KEYINPUT49), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n348), .B1(new_n721), .B2(new_n553), .ZN(new_n722));
  XOR2_X1   g521(.A(new_n722), .B(KEYINPUT105), .Z(new_n723));
  NAND2_X1  g522(.A1(new_n718), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n721), .A2(new_n553), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n724), .B(new_n725), .ZN(G1333gat));
  OAI21_X1  g525(.A(G71gat), .B1(new_n717), .B2(new_n647), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n718), .A2(new_n485), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n727), .B1(new_n728), .B2(G71gat), .ZN(new_n729));
  XOR2_X1   g528(.A(new_n729), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g529(.A1(new_n717), .A2(new_n399), .ZN(new_n731));
  XOR2_X1   g530(.A(KEYINPUT106), .B(G78gat), .Z(new_n732));
  XNOR2_X1  g531(.A(new_n731), .B(new_n732), .ZN(G1335gat));
  NOR2_X1   g532(.A1(new_n579), .A2(new_n551), .ZN(new_n734));
  AND3_X1   g533(.A1(new_n657), .A2(new_n669), .A3(new_n734), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n735), .A2(KEYINPUT107), .A3(new_n473), .A4(new_n631), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT107), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n657), .A2(new_n669), .A3(new_n631), .A4(new_n734), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n737), .B1(new_n738), .B2(new_n469), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n736), .A2(G85gat), .A3(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT108), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n668), .A2(new_n608), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n742), .A2(KEYINPUT51), .A3(new_n734), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  AOI21_X1  g543(.A(KEYINPUT51), .B1(new_n742), .B2(new_n734), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n741), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n742), .A2(new_n734), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT51), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n749), .A2(KEYINPUT108), .A3(new_n743), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n469), .A2(new_n632), .A3(G85gat), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n746), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n740), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(KEYINPUT109), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT109), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n740), .A2(new_n752), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n754), .A2(new_n756), .ZN(G1336gat));
  INV_X1    g556(.A(KEYINPUT52), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n464), .A2(new_n632), .A3(G92gat), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n759), .B1(new_n744), .B2(new_n745), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n758), .B1(new_n760), .B2(KEYINPUT110), .ZN(new_n761));
  OAI21_X1  g560(.A(G92gat), .B1(new_n738), .B2(new_n464), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n761), .B(new_n763), .ZN(G1337gat));
  OAI21_X1  g563(.A(G99gat), .B1(new_n738), .B2(new_n647), .ZN(new_n765));
  INV_X1    g564(.A(G99gat), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n746), .A2(new_n750), .A3(new_n766), .A4(new_n485), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n765), .B1(new_n767), .B2(new_n632), .ZN(G1338gat));
  NAND3_X1  g567(.A1(new_n735), .A2(new_n472), .A3(new_n631), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(G106gat), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT53), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n744), .A2(new_n745), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n399), .A2(new_n632), .A3(G106gat), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n770), .B(new_n771), .C1(new_n772), .C2(new_n774), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n774), .A2(KEYINPUT111), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n772), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n774), .A2(KEYINPUT111), .ZN(new_n778));
  AOI22_X1  g577(.A1(new_n777), .A2(new_n778), .B1(G106gat), .B2(new_n769), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n775), .B1(new_n779), .B2(new_n771), .ZN(G1339gat));
  INV_X1    g579(.A(KEYINPUT112), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n621), .A2(new_n616), .A3(new_n622), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n624), .A2(new_n781), .A3(KEYINPUT54), .A4(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(KEYINPUT54), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT54), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n781), .A2(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n784), .B1(new_n623), .B2(new_n786), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n783), .A2(new_n787), .A3(new_n628), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT55), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n783), .A2(new_n787), .A3(KEYINPUT55), .A4(new_n628), .ZN(new_n791));
  AND3_X1   g590(.A1(new_n790), .A2(new_n629), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n551), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n547), .B(new_n548), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n520), .A2(new_n522), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n517), .A2(new_n531), .A3(new_n530), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n542), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n794), .A2(new_n631), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n793), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(new_n608), .ZN(new_n800));
  AND3_X1   g599(.A1(new_n604), .A2(new_n605), .A3(new_n607), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n794), .A2(new_n797), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n801), .A2(new_n802), .A3(new_n792), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n579), .B1(new_n800), .B2(new_n803), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n609), .A2(new_n551), .A3(new_n631), .ZN(new_n805));
  OR2_X1    g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n806), .A2(new_n473), .ZN(new_n807));
  INV_X1    g606(.A(new_n485), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n808), .A2(new_n348), .A3(new_n472), .ZN(new_n809));
  AND2_X1   g608(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(G113gat), .B1(new_n811), .B2(new_n671), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n807), .A2(new_n399), .A3(new_n477), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n813), .A2(new_n348), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(new_n551), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n812), .B1(new_n815), .B2(G113gat), .ZN(new_n816));
  XNOR2_X1  g615(.A(new_n816), .B(KEYINPUT113), .ZN(G1340gat));
  OAI21_X1  g616(.A(G120gat), .B1(new_n811), .B2(new_n632), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n814), .A2(new_n207), .A3(new_n631), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(G1341gat));
  AOI21_X1  g619(.A(G127gat), .B1(new_n814), .B2(new_n579), .ZN(new_n821));
  AND3_X1   g620(.A1(new_n810), .A2(G127gat), .A3(new_n579), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n821), .A2(new_n822), .ZN(G1342gat));
  NOR4_X1   g622(.A1(new_n813), .A2(G134gat), .A3(new_n348), .A4(new_n608), .ZN(new_n824));
  XNOR2_X1  g623(.A(KEYINPUT114), .B(KEYINPUT56), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  OR2_X1    g625(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(G134gat), .B1(new_n811), .B2(new_n608), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n824), .A2(new_n826), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(G1343gat));
  INV_X1    g629(.A(new_n579), .ZN(new_n831));
  OR2_X1    g630(.A1(new_n790), .A2(KEYINPUT115), .ZN(new_n832));
  NOR2_X1   g631(.A1(KEYINPUT115), .A2(KEYINPUT55), .ZN(new_n833));
  OR2_X1    g632(.A1(new_n788), .A2(new_n833), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n551), .A2(new_n832), .A3(new_n629), .A4(new_n834), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n835), .A2(KEYINPUT116), .A3(new_n798), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(KEYINPUT116), .B1(new_n835), .B2(new_n798), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n837), .A2(new_n838), .A3(new_n801), .ZN(new_n839));
  INV_X1    g638(.A(new_n803), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n831), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(new_n805), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n843), .A2(KEYINPUT117), .A3(KEYINPUT57), .A4(new_n472), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n835), .A2(new_n798), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT116), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n847), .A2(new_n608), .A3(new_n836), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n579), .B1(new_n848), .B2(new_n803), .ZN(new_n849));
  OAI211_X1 g648(.A(KEYINPUT57), .B(new_n472), .C1(new_n849), .C2(new_n805), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n472), .B1(new_n804), .B2(new_n805), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT57), .ZN(new_n852));
  AOI21_X1  g651(.A(KEYINPUT117), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n648), .A2(new_n469), .A3(new_n348), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n844), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  OAI21_X1  g655(.A(G141gat), .B1(new_n856), .B2(new_n671), .ZN(new_n857));
  NAND2_X1  g656(.A1(KEYINPUT118), .A2(KEYINPUT58), .ZN(new_n858));
  NOR4_X1   g657(.A1(new_n851), .A2(new_n469), .A3(new_n348), .A4(new_n648), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n859), .A2(new_n215), .A3(new_n551), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n857), .A2(new_n858), .A3(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(KEYINPUT118), .A2(KEYINPUT58), .ZN(new_n862));
  XNOR2_X1  g661(.A(new_n862), .B(KEYINPUT119), .ZN(new_n863));
  INV_X1    g662(.A(new_n863), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n861), .B(new_n864), .ZN(G1344gat));
  NAND4_X1  g664(.A1(new_n844), .A2(new_n854), .A3(new_n631), .A4(new_n855), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT59), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n866), .A2(new_n867), .A3(G148gat), .ZN(new_n868));
  OAI211_X1 g667(.A(new_n852), .B(new_n472), .C1(new_n849), .C2(new_n805), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n851), .A2(KEYINPUT57), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n869), .A2(new_n631), .A3(new_n855), .A4(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(G148gat), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(KEYINPUT59), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n868), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n859), .A2(new_n213), .A3(new_n631), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT120), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n874), .A2(KEYINPUT120), .A3(new_n875), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(G1345gat));
  AOI21_X1  g679(.A(G155gat), .B1(new_n859), .B2(new_n579), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n856), .A2(new_n831), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n881), .B1(new_n882), .B2(G155gat), .ZN(G1346gat));
  NOR2_X1   g682(.A1(new_n856), .A2(new_n608), .ZN(new_n884));
  OR2_X1    g683(.A1(new_n884), .A2(KEYINPUT121), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(KEYINPUT121), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n885), .A2(G162gat), .A3(new_n886), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n859), .A2(new_n220), .A3(new_n801), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(G1347gat));
  NAND2_X1  g688(.A1(new_n469), .A2(new_n348), .ZN(new_n890));
  AOI211_X1 g689(.A(new_n472), .B(new_n890), .C1(new_n461), .C2(new_n460), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n806), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n892), .A2(new_n281), .A3(new_n551), .ZN(new_n893));
  XOR2_X1   g692(.A(new_n893), .B(KEYINPUT122), .Z(new_n894));
  NOR2_X1   g693(.A1(new_n808), .A2(new_n890), .ZN(new_n895));
  OR2_X1    g694(.A1(new_n895), .A2(KEYINPUT123), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n472), .B1(new_n895), .B2(KEYINPUT123), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n806), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(G169gat), .B1(new_n898), .B2(new_n671), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n894), .A2(new_n899), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n900), .B(KEYINPUT124), .ZN(G1348gat));
  AOI21_X1  g700(.A(G176gat), .B1(new_n892), .B2(new_n631), .ZN(new_n902));
  INV_X1    g701(.A(new_n898), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n631), .A2(new_n306), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n902), .B1(new_n903), .B2(new_n904), .ZN(G1349gat));
  NAND3_X1  g704(.A1(new_n892), .A2(new_n318), .A3(new_n579), .ZN(new_n906));
  OAI21_X1  g705(.A(G183gat), .B1(new_n898), .B2(new_n831), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g707(.A(new_n908), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g708(.A(G190gat), .B1(new_n898), .B2(new_n608), .ZN(new_n910));
  OR2_X1    g709(.A1(new_n910), .A2(KEYINPUT125), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(KEYINPUT125), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n911), .A2(KEYINPUT61), .A3(new_n912), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n892), .A2(new_n319), .A3(new_n801), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT61), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n910), .A2(KEYINPUT125), .A3(new_n915), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n913), .A2(new_n914), .A3(new_n916), .ZN(G1351gat));
  AND2_X1   g716(.A1(new_n869), .A2(new_n870), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n648), .A2(new_n890), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OR3_X1    g719(.A1(new_n920), .A2(KEYINPUT126), .A3(new_n671), .ZN(new_n921));
  OAI21_X1  g720(.A(KEYINPUT126), .B1(new_n920), .B2(new_n671), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n921), .A2(G197gat), .A3(new_n922), .ZN(new_n923));
  NOR3_X1   g722(.A1(new_n851), .A2(new_n648), .A3(new_n890), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n924), .A2(new_n539), .A3(new_n551), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n923), .A2(new_n925), .ZN(G1352gat));
  INV_X1    g725(.A(G204gat), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n924), .A2(new_n927), .A3(new_n631), .ZN(new_n928));
  XOR2_X1   g727(.A(new_n928), .B(KEYINPUT62), .Z(new_n929));
  AND3_X1   g728(.A1(new_n918), .A2(new_n631), .A3(new_n919), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n929), .B1(new_n927), .B2(new_n930), .ZN(G1353gat));
  NAND3_X1  g730(.A1(new_n924), .A2(new_n273), .A3(new_n579), .ZN(new_n932));
  NAND4_X1  g731(.A1(new_n869), .A2(new_n579), .A3(new_n870), .A4(new_n919), .ZN(new_n933));
  AND3_X1   g732(.A1(new_n933), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n934));
  AOI21_X1  g733(.A(KEYINPUT63), .B1(new_n933), .B2(G211gat), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n932), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT127), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n936), .B(new_n937), .ZN(G1354gat));
  OAI21_X1  g737(.A(G218gat), .B1(new_n920), .B2(new_n608), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n924), .A2(new_n274), .A3(new_n801), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(G1355gat));
endmodule


