//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 0 1 1 0 1 1 1 0 1 1 0 0 0 0 1 0 0 0 1 0 1 0 1 1 1 0 1 1 1 1 1 1 1 0 1 1 1 0 1 1 1 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:31 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n560, new_n562, new_n563, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n585, new_n586, new_n587, new_n588, new_n589,
    new_n590, new_n591, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n629, new_n630,
    new_n633, new_n634, new_n635, new_n636, new_n638, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1253, new_n1254, new_n1255;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT64), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  AOI22_X1  g030(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n453), .ZN(G319));
  XNOR2_X1  g031(.A(KEYINPUT3), .B(G2104), .ZN(new_n457));
  AOI22_X1  g032(.A1(new_n457), .A2(G137), .B1(G101), .B2(G2104), .ZN(new_n458));
  OAI21_X1  g033(.A(KEYINPUT66), .B1(new_n458), .B2(G2105), .ZN(new_n459));
  INV_X1    g034(.A(KEYINPUT65), .ZN(new_n460));
  AOI22_X1  g035(.A1(new_n457), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  OAI21_X1  g037(.A(new_n460), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(G101), .A2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G137), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n464), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT66), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n471), .A2(new_n472), .A3(new_n462), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n466), .A2(new_n468), .A3(G125), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n476), .A2(KEYINPUT65), .A3(G2105), .ZN(new_n477));
  NAND4_X1  g052(.A1(new_n459), .A2(new_n463), .A3(new_n473), .A4(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  OAI21_X1  g054(.A(KEYINPUT67), .B1(new_n469), .B2(G2105), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT67), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n457), .A2(new_n481), .A3(new_n462), .ZN(new_n482));
  AND2_X1   g057(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n457), .A2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  AOI22_X1  g060(.A1(new_n483), .A2(G136), .B1(G124), .B2(new_n485), .ZN(new_n486));
  OR2_X1    g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n488));
  XNOR2_X1  g063(.A(new_n488), .B(KEYINPUT68), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT69), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n486), .A2(KEYINPUT69), .A3(new_n489), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(G162));
  NAND3_X1  g069(.A1(new_n466), .A2(new_n468), .A3(G126), .ZN(new_n495));
  NAND2_X1  g070(.A1(G114), .A2(G2104), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G2105), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n465), .A2(G2105), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(G102), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n466), .A2(new_n468), .A3(G138), .A4(new_n462), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n457), .A2(KEYINPUT4), .A3(G138), .A4(new_n462), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n498), .A2(new_n500), .A3(new_n503), .A4(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(G164));
  NAND2_X1  g081(.A1(G75), .A2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(KEYINPUT5), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT70), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT5), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n510), .B1(new_n511), .B2(G543), .ZN(new_n512));
  NOR3_X1   g087(.A1(new_n508), .A2(KEYINPUT70), .A3(KEYINPUT5), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n509), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G62), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n507), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  XNOR2_X1  g091(.A(KEYINPUT6), .B(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G543), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n516), .A2(G651), .B1(G50), .B2(new_n519), .ZN(new_n520));
  OAI211_X1 g095(.A(new_n517), .B(new_n509), .C1(new_n512), .C2(new_n513), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(KEYINPUT71), .ZN(new_n522));
  OAI21_X1  g097(.A(KEYINPUT70), .B1(new_n508), .B2(KEYINPUT5), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n510), .A2(new_n511), .A3(G543), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n523), .A2(new_n524), .B1(KEYINPUT5), .B2(new_n508), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT71), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n525), .A2(new_n526), .A3(new_n517), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n522), .A2(G88), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n520), .A2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(G166));
  NAND3_X1  g105(.A1(new_n522), .A2(G89), .A3(new_n527), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n519), .A2(G51), .ZN(new_n532));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT7), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n525), .A2(G63), .A3(G651), .ZN(new_n535));
  NAND4_X1  g110(.A1(new_n531), .A2(new_n532), .A3(new_n534), .A4(new_n535), .ZN(G286));
  INV_X1    g111(.A(G286), .ZN(G168));
  INV_X1    g112(.A(G64), .ZN(new_n538));
  INV_X1    g113(.A(G77), .ZN(new_n539));
  OAI22_X1  g114(.A1(new_n514), .A2(new_n538), .B1(new_n539), .B2(new_n508), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(KEYINPUT72), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT72), .ZN(new_n542));
  OAI221_X1 g117(.A(new_n542), .B1(new_n539), .B2(new_n508), .C1(new_n514), .C2(new_n538), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n541), .A2(G651), .A3(new_n543), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n522), .A2(G90), .A3(new_n527), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT73), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n519), .A2(G52), .ZN(new_n547));
  AND3_X1   g122(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n546), .B1(new_n545), .B2(new_n547), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n544), .B1(new_n548), .B2(new_n549), .ZN(G301));
  INV_X1    g125(.A(G301), .ZN(G171));
  NAND2_X1  g126(.A1(G68), .A2(G543), .ZN(new_n552));
  INV_X1    g127(.A(G56), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n514), .B2(new_n553), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n554), .A2(G651), .B1(G43), .B2(new_n519), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n522), .A2(G81), .A3(new_n527), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(G153));
  AND3_X1   g134(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G36), .ZN(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n560), .A2(new_n563), .ZN(G188));
  INV_X1    g139(.A(KEYINPUT74), .ZN(new_n565));
  AOI21_X1  g140(.A(KEYINPUT75), .B1(new_n565), .B2(KEYINPUT9), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n566), .B1(KEYINPUT75), .B2(KEYINPUT9), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n519), .A2(G53), .A3(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(G53), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n566), .B1(new_n518), .B2(new_n569), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n525), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n571));
  INV_X1    g146(.A(G651), .ZN(new_n572));
  OAI211_X1 g147(.A(new_n568), .B(new_n570), .C1(new_n571), .C2(new_n572), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n522), .A2(G91), .A3(new_n527), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(new_n575));
  OAI21_X1  g150(.A(KEYINPUT76), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(G78), .A2(G543), .ZN(new_n577));
  INV_X1    g152(.A(G65), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n514), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n519), .A2(G53), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n579), .A2(G651), .B1(new_n580), .B2(new_n566), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT76), .ZN(new_n582));
  NAND4_X1  g157(.A1(new_n581), .A2(new_n582), .A3(new_n574), .A4(new_n568), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n576), .A2(new_n583), .ZN(G299));
  INV_X1    g159(.A(KEYINPUT77), .ZN(new_n585));
  AND3_X1   g160(.A1(new_n522), .A2(G88), .A3(new_n527), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n519), .A2(G50), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n525), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n588), .B2(new_n572), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n585), .B1(new_n586), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n520), .A2(KEYINPUT77), .A3(new_n528), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(G303));
  NAND3_X1  g167(.A1(new_n522), .A2(G87), .A3(new_n527), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n517), .A2(G49), .A3(G543), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT78), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n594), .B(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(G651), .B1(new_n525), .B2(G74), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n593), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(KEYINPUT79), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT79), .ZN(new_n600));
  NAND4_X1  g175(.A1(new_n593), .A2(new_n596), .A3(new_n600), .A4(new_n597), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n599), .A2(new_n601), .ZN(G288));
  NAND3_X1  g177(.A1(new_n522), .A2(G86), .A3(new_n527), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n519), .A2(G48), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n525), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n606), .B2(new_n572), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(G305));
  NAND3_X1  g184(.A1(new_n522), .A2(G85), .A3(new_n527), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n525), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n611));
  XNOR2_X1  g186(.A(KEYINPUT80), .B(G47), .ZN(new_n612));
  OAI221_X1 g187(.A(new_n610), .B1(new_n572), .B2(new_n611), .C1(new_n518), .C2(new_n612), .ZN(G290));
  NAND3_X1  g188(.A1(new_n522), .A2(G92), .A3(new_n527), .ZN(new_n614));
  XOR2_X1   g189(.A(KEYINPUT81), .B(KEYINPUT10), .Z(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(G79), .A2(G543), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT82), .ZN(new_n619));
  INV_X1    g194(.A(G66), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n514), .B2(new_n620), .ZN(new_n621));
  AOI22_X1  g196(.A1(new_n621), .A2(G651), .B1(G54), .B2(new_n519), .ZN(new_n622));
  NAND4_X1  g197(.A1(new_n522), .A2(new_n527), .A3(G92), .A4(new_n615), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n617), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  INV_X1    g199(.A(G868), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(G171), .B2(new_n625), .ZN(G284));
  OAI21_X1  g202(.A(new_n626), .B1(G171), .B2(new_n625), .ZN(G321));
  NOR2_X1   g203(.A1(G286), .A2(new_n625), .ZN(new_n629));
  INV_X1    g204(.A(G299), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n629), .B1(new_n630), .B2(new_n625), .ZN(G297));
  AOI21_X1  g206(.A(new_n629), .B1(new_n630), .B2(new_n625), .ZN(G280));
  OR2_X1    g207(.A1(new_n624), .A2(G559), .ZN(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(new_n634));
  INV_X1    g209(.A(new_n624), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n634), .B1(G860), .B2(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(KEYINPUT83), .Z(G148));
  NAND2_X1  g212(.A1(new_n557), .A2(new_n625), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n638), .B1(new_n634), .B2(new_n625), .ZN(G323));
  XNOR2_X1  g214(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g215(.A1(new_n483), .A2(G135), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n485), .A2(G123), .ZN(new_n642));
  OR2_X1    g217(.A1(G99), .A2(G2105), .ZN(new_n643));
  OAI211_X1 g218(.A(new_n643), .B(G2104), .C1(G111), .C2(new_n462), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n641), .A2(new_n642), .A3(new_n644), .ZN(new_n645));
  INV_X1    g220(.A(KEYINPUT85), .ZN(new_n646));
  AOI22_X1  g221(.A1(new_n645), .A2(G2096), .B1(new_n646), .B2(G2100), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n457), .A2(new_n499), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT12), .ZN(new_n649));
  XOR2_X1   g224(.A(KEYINPUT84), .B(KEYINPUT13), .Z(new_n650));
  NOR2_X1   g225(.A1(new_n646), .A2(G2100), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n649), .B(new_n652), .ZN(new_n653));
  OAI211_X1 g228(.A(new_n647), .B(new_n653), .C1(G2096), .C2(new_n645), .ZN(G156));
  XNOR2_X1  g229(.A(KEYINPUT15), .B(G2430), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2435), .ZN(new_n656));
  XOR2_X1   g231(.A(G2427), .B(G2438), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n658), .A2(KEYINPUT14), .ZN(new_n659));
  XOR2_X1   g234(.A(G2451), .B(G2454), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(KEYINPUT86), .B(KEYINPUT16), .Z(new_n662));
  XNOR2_X1  g237(.A(G1341), .B(G1348), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n661), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2443), .B(G2446), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n665), .B(new_n666), .Z(new_n667));
  AND2_X1   g242(.A1(new_n667), .A2(G14), .ZN(G401));
  XOR2_X1   g243(.A(G2084), .B(G2090), .Z(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2067), .B(G2678), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT87), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G2072), .B(G2078), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n670), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n675), .B(KEYINPUT88), .Z(new_n676));
  XOR2_X1   g251(.A(new_n674), .B(KEYINPUT17), .Z(new_n677));
  OAI21_X1  g252(.A(new_n676), .B1(new_n677), .B2(new_n672), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n677), .A2(new_n672), .A3(new_n669), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n673), .A2(new_n674), .A3(new_n669), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n680), .B(KEYINPUT18), .Z(new_n681));
  NAND3_X1  g256(.A1(new_n678), .A2(new_n679), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(G2096), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(G2100), .Z(G227));
  XOR2_X1   g259(.A(G1956), .B(G2474), .Z(new_n685));
  XOR2_X1   g260(.A(G1961), .B(G1966), .Z(new_n686));
  NOR2_X1   g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1971), .B(G1976), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT19), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n685), .A2(new_n686), .ZN(new_n692));
  OR2_X1    g267(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(KEYINPUT20), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n691), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n688), .A2(new_n690), .A3(new_n692), .ZN(new_n696));
  OAI211_X1 g271(.A(new_n695), .B(new_n696), .C1(new_n694), .C2(new_n693), .ZN(new_n697));
  XOR2_X1   g272(.A(G1991), .B(G1996), .Z(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT89), .B(KEYINPUT90), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n697), .B(new_n700), .ZN(new_n701));
  XOR2_X1   g276(.A(G1981), .B(G1986), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT91), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n701), .B(new_n705), .ZN(G229));
  INV_X1    g281(.A(KEYINPUT28), .ZN(new_n707));
  AND2_X1   g282(.A1(KEYINPUT92), .A2(G29), .ZN(new_n708));
  NOR2_X1   g283(.A1(KEYINPUT92), .A2(G29), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(G26), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n707), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(new_n710), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n713), .A2(KEYINPUT28), .A3(G26), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n483), .A2(G140), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n485), .A2(G128), .ZN(new_n716));
  OR2_X1    g291(.A1(G104), .A2(G2105), .ZN(new_n717));
  OAI211_X1 g292(.A(new_n717), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n715), .A2(new_n716), .A3(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT96), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND4_X1  g296(.A1(new_n715), .A2(KEYINPUT96), .A3(new_n716), .A4(new_n718), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(G29), .ZN(new_n725));
  OAI211_X1 g300(.A(new_n712), .B(new_n714), .C1(new_n724), .C2(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(G2067), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n713), .B1(new_n492), .B2(new_n493), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n710), .A2(G35), .ZN(new_n729));
  OR3_X1    g304(.A1(new_n728), .A2(KEYINPUT29), .A3(new_n729), .ZN(new_n730));
  OAI21_X1  g305(.A(KEYINPUT29), .B1(new_n728), .B2(new_n729), .ZN(new_n731));
  AOI21_X1  g306(.A(G2090), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n558), .A2(G16), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G16), .B2(G19), .ZN(new_n734));
  INV_X1    g309(.A(G1341), .ZN(new_n735));
  AND2_X1   g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT30), .B(G28), .ZN(new_n737));
  AND2_X1   g312(.A1(new_n737), .A2(new_n725), .ZN(new_n738));
  NOR4_X1   g313(.A1(new_n727), .A2(new_n732), .A3(new_n736), .A4(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(G171), .A2(G16), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(G5), .B2(G16), .ZN(new_n741));
  INV_X1    g316(.A(G1961), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  XOR2_X1   g318(.A(KEYINPUT27), .B(G1996), .Z(new_n744));
  INV_X1    g319(.A(new_n744), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n480), .A2(G141), .A3(new_n482), .ZN(new_n746));
  NAND3_X1  g321(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT26), .Z(new_n748));
  AND2_X1   g323(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  AND3_X1   g324(.A1(new_n457), .A2(G129), .A3(G2105), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT99), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n499), .A2(G105), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n749), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n753), .A2(G29), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n725), .A2(G32), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT100), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n743), .B1(new_n745), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n483), .A2(G139), .ZN(new_n760));
  AOI22_X1  g335(.A1(new_n457), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n761));
  OR2_X1    g336(.A1(new_n761), .A2(new_n462), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n499), .A2(G103), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT25), .Z(new_n764));
  NAND3_X1  g339(.A1(new_n760), .A2(new_n762), .A3(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n766), .A2(G29), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G29), .B2(G33), .ZN(new_n768));
  INV_X1    g343(.A(G2072), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(G2084), .ZN(new_n771));
  XOR2_X1   g346(.A(KEYINPUT97), .B(KEYINPUT24), .Z(new_n772));
  INV_X1    g347(.A(G34), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n710), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT98), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(new_n773), .B2(new_n772), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(new_n725), .B2(new_n478), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n770), .B1(new_n771), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n713), .A2(G27), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G164), .B2(new_n713), .ZN(new_n780));
  INV_X1    g355(.A(G2078), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(G168), .A2(G16), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G16), .B2(G21), .ZN(new_n784));
  INV_X1    g359(.A(G1966), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  AND2_X1   g361(.A1(new_n786), .A2(KEYINPUT102), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n786), .A2(KEYINPUT102), .ZN(new_n788));
  OAI211_X1 g363(.A(new_n778), .B(new_n782), .C1(new_n787), .C2(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(new_n789), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n784), .A2(new_n785), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(KEYINPUT101), .Z(new_n792));
  NAND4_X1  g367(.A1(new_n739), .A2(new_n759), .A3(new_n790), .A4(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(G16), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n794), .A2(KEYINPUT23), .A3(G20), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT23), .ZN(new_n796));
  INV_X1    g371(.A(G20), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n796), .B1(new_n797), .B2(G16), .ZN(new_n798));
  OAI211_X1 g373(.A(new_n795), .B(new_n798), .C1(new_n630), .C2(new_n794), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(G1956), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n768), .A2(new_n769), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(new_n758), .B2(new_n745), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n730), .A2(G2090), .A3(new_n731), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n734), .A2(new_n735), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n794), .A2(G4), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(new_n635), .B2(new_n794), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n807), .A2(G1348), .ZN(new_n808));
  AND2_X1   g383(.A1(new_n807), .A2(G1348), .ZN(new_n809));
  AOI211_X1 g384(.A(new_n808), .B(new_n809), .C1(new_n742), .C2(new_n741), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n803), .A2(new_n804), .A3(new_n805), .A4(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n793), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g387(.A(KEYINPUT31), .B(G11), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n794), .A2(G22), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(G166), .B2(new_n794), .ZN(new_n815));
  INV_X1    g390(.A(G1971), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n794), .A2(G23), .ZN(new_n818));
  INV_X1    g393(.A(new_n598), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n818), .B1(new_n819), .B2(new_n794), .ZN(new_n820));
  XNOR2_X1  g395(.A(KEYINPUT33), .B(G1976), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT94), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n820), .B(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n794), .A2(G6), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(new_n608), .B2(new_n794), .ZN(new_n825));
  XOR2_X1   g400(.A(KEYINPUT32), .B(G1981), .Z(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n817), .A2(new_n823), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n828), .A2(KEYINPUT34), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT95), .ZN(new_n830));
  MUX2_X1   g405(.A(G24), .B(G290), .S(G16), .Z(new_n831));
  INV_X1    g406(.A(G1986), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  AND3_X1   g408(.A1(new_n829), .A2(new_n830), .A3(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT36), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n828), .A2(KEYINPUT34), .ZN(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(new_n483), .ZN(new_n838));
  INV_X1    g413(.A(G131), .ZN(new_n839));
  OR3_X1    g414(.A1(new_n838), .A2(KEYINPUT93), .A3(new_n839), .ZN(new_n840));
  OR2_X1    g415(.A1(G95), .A2(G2105), .ZN(new_n841));
  INV_X1    g416(.A(G107), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n465), .B1(new_n842), .B2(G2105), .ZN(new_n843));
  AOI22_X1  g418(.A1(new_n485), .A2(G119), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g419(.A(KEYINPUT93), .B1(new_n838), .B2(new_n839), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n840), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  MUX2_X1   g421(.A(G25), .B(new_n846), .S(new_n710), .Z(new_n847));
  XNOR2_X1  g422(.A(KEYINPUT35), .B(G1991), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n847), .B(new_n848), .Z(new_n849));
  NAND4_X1  g424(.A1(new_n834), .A2(new_n835), .A3(new_n837), .A4(new_n849), .ZN(new_n850));
  NAND4_X1  g425(.A1(new_n849), .A2(new_n830), .A3(new_n829), .A4(new_n833), .ZN(new_n851));
  OAI21_X1  g426(.A(KEYINPUT36), .B1(new_n851), .B2(new_n836), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  AND3_X1   g428(.A1(new_n812), .A2(new_n813), .A3(new_n853), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n645), .A2(new_n713), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  OR2_X1    g431(.A1(new_n777), .A2(new_n771), .ZN(new_n857));
  NAND4_X1  g432(.A1(new_n854), .A2(KEYINPUT103), .A3(new_n856), .A4(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT103), .ZN(new_n859));
  NAND4_X1  g434(.A1(new_n812), .A2(new_n853), .A3(new_n857), .A4(new_n813), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n859), .B1(new_n860), .B2(new_n855), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n858), .A2(new_n861), .ZN(G311));
  NAND3_X1  g437(.A1(new_n854), .A2(new_n856), .A3(new_n857), .ZN(G150));
  OAI211_X1 g438(.A(G67), .B(new_n509), .C1(new_n512), .C2(new_n513), .ZN(new_n864));
  NAND2_X1  g439(.A1(G80), .A2(G543), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  AOI22_X1  g441(.A1(new_n866), .A2(G651), .B1(G55), .B2(new_n519), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n522), .A2(G93), .A3(new_n527), .ZN(new_n868));
  AND3_X1   g443(.A1(new_n867), .A2(KEYINPUT104), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(KEYINPUT104), .B1(new_n867), .B2(new_n868), .ZN(new_n870));
  OR2_X1    g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n872), .A2(G860), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(KEYINPUT105), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT37), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n557), .B1(new_n869), .B2(new_n870), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n867), .A2(new_n868), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n558), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(KEYINPUT39), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n635), .A2(G559), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(KEYINPUT38), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n880), .B(new_n882), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n875), .B1(new_n883), .B2(G860), .ZN(G145));
  AND3_X1   g459(.A1(new_n492), .A2(new_n478), .A3(new_n493), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n478), .B1(new_n492), .B2(new_n493), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n645), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(G162), .A2(G160), .ZN(new_n888));
  INV_X1    g463(.A(new_n645), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n492), .A2(new_n478), .A3(new_n493), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  AND3_X1   g466(.A1(new_n887), .A2(new_n891), .A3(new_n765), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n765), .B1(new_n887), .B2(new_n891), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n483), .A2(G142), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n485), .A2(G130), .ZN(new_n896));
  OR2_X1    g471(.A1(G106), .A2(G2105), .ZN(new_n897));
  OAI211_X1 g472(.A(new_n897), .B(G2104), .C1(G118), .C2(new_n462), .ZN(new_n898));
  NAND4_X1  g473(.A1(new_n753), .A2(new_n895), .A3(new_n896), .A4(new_n898), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n895), .A2(new_n896), .A3(new_n898), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n900), .A2(new_n752), .A3(new_n751), .A4(new_n749), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n902), .A2(new_n724), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n723), .A2(new_n899), .A3(new_n901), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n903), .A2(G164), .A3(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(G164), .B1(new_n903), .B2(new_n904), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n846), .B(new_n649), .ZN(new_n908));
  NOR3_X1   g483(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n908), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n903), .A2(new_n904), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(new_n505), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n910), .B1(new_n912), .B2(new_n905), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n894), .B1(new_n909), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n908), .B1(new_n906), .B2(new_n907), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n912), .A2(new_n905), .A3(new_n910), .ZN(new_n916));
  OAI211_X1 g491(.A(new_n915), .B(new_n916), .C1(new_n893), .C2(new_n892), .ZN(new_n917));
  INV_X1    g492(.A(G37), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n914), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(KEYINPUT106), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT107), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT106), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n914), .A2(new_n917), .A3(new_n922), .A4(new_n918), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n920), .A2(new_n921), .A3(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n921), .B1(new_n920), .B2(new_n923), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT40), .ZN(new_n927));
  NOR3_X1   g502(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n920), .A2(new_n923), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(KEYINPUT107), .ZN(new_n930));
  AOI21_X1  g505(.A(KEYINPUT40), .B1(new_n930), .B2(new_n924), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n928), .A2(new_n931), .ZN(G395));
  XNOR2_X1  g507(.A(G290), .B(new_n819), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n608), .B(new_n529), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n933), .B(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT108), .ZN(new_n936));
  OR3_X1    g511(.A1(new_n935), .A2(new_n936), .A3(KEYINPUT42), .ZN(new_n937));
  OAI21_X1  g512(.A(KEYINPUT42), .B1(new_n935), .B2(new_n936), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT109), .ZN(new_n939));
  INV_X1    g514(.A(new_n935), .ZN(new_n940));
  AOI22_X1  g515(.A1(new_n937), .A2(new_n938), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(G299), .A2(new_n624), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n635), .A2(new_n576), .A3(new_n583), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  NOR2_X1   g521(.A1(G299), .A2(new_n624), .ZN(new_n947));
  AND2_X1   g522(.A1(new_n617), .A2(new_n623), .ZN(new_n948));
  AOI22_X1  g523(.A1(new_n948), .A2(new_n622), .B1(new_n576), .B2(new_n583), .ZN(new_n949));
  OAI21_X1  g524(.A(KEYINPUT41), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT41), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n943), .A2(new_n944), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n879), .B(new_n633), .ZN(new_n954));
  MUX2_X1   g529(.A(new_n946), .B(new_n953), .S(new_n954), .Z(new_n955));
  NAND3_X1  g530(.A1(new_n937), .A2(new_n939), .A3(new_n938), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n942), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n955), .ZN(new_n958));
  INV_X1    g533(.A(new_n956), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n958), .B1(new_n959), .B2(new_n941), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n625), .B1(new_n957), .B2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT110), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n871), .A2(G868), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n962), .A2(new_n963), .A3(new_n965), .ZN(new_n966));
  OAI21_X1  g541(.A(KEYINPUT110), .B1(new_n961), .B2(new_n964), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(G295));
  NAND2_X1  g543(.A1(new_n962), .A2(new_n965), .ZN(G331));
  NAND2_X1  g544(.A1(G301), .A2(G168), .ZN(new_n970));
  OAI211_X1 g545(.A(G286), .B(new_n544), .C1(new_n548), .C2(new_n549), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n970), .A2(new_n878), .A3(new_n876), .A4(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  AOI22_X1  g548(.A1(new_n970), .A2(new_n971), .B1(new_n878), .B2(new_n876), .ZN(new_n974));
  OAI21_X1  g549(.A(KEYINPUT111), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT111), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n972), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n975), .A2(new_n946), .A3(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT112), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n953), .B1(new_n973), .B2(new_n974), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n975), .A2(KEYINPUT112), .A3(new_n946), .A4(new_n977), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n980), .A2(new_n981), .A3(new_n935), .A4(new_n982), .ZN(new_n983));
  AND2_X1   g558(.A1(new_n983), .A2(new_n918), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n945), .A2(KEYINPUT113), .A3(KEYINPUT41), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT113), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n950), .A2(new_n986), .A3(new_n952), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n545), .A2(new_n547), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(KEYINPUT73), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(G286), .B1(new_n991), .B2(new_n544), .ZN(new_n992));
  INV_X1    g567(.A(new_n971), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n879), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n976), .B1(new_n994), .B2(new_n972), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n992), .A2(new_n993), .ZN(new_n996));
  INV_X1    g571(.A(new_n879), .ZN(new_n997));
  AOI21_X1  g572(.A(KEYINPUT111), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  OAI211_X1 g573(.A(new_n985), .B(new_n987), .C1(new_n995), .C2(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n946), .A2(new_n994), .A3(new_n972), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(new_n940), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(KEYINPUT114), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT114), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1001), .A2(new_n1004), .A3(new_n940), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT43), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n984), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n995), .A2(new_n998), .ZN(new_n1009));
  AOI21_X1  g584(.A(KEYINPUT112), .B1(new_n1009), .B2(new_n946), .ZN(new_n1010));
  NOR4_X1   g585(.A1(new_n995), .A2(new_n998), .A3(new_n979), .A4(new_n945), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n935), .B1(new_n1012), .B2(new_n981), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n983), .A2(new_n918), .ZN(new_n1014));
  OAI21_X1  g589(.A(KEYINPUT43), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1008), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT44), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1004), .B1(new_n1001), .B2(new_n940), .ZN(new_n1019));
  AOI211_X1 g594(.A(KEYINPUT114), .B(new_n935), .C1(new_n999), .C2(new_n1000), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n918), .B(new_n983), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1017), .B1(new_n1021), .B2(KEYINPUT43), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n980), .A2(new_n981), .A3(new_n982), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(new_n940), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1024), .A2(new_n1007), .A3(new_n918), .A4(new_n983), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT115), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n984), .A2(KEYINPUT115), .A3(new_n1007), .A4(new_n1024), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1022), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1018), .A2(new_n1029), .ZN(G397));
  INV_X1    g605(.A(G40), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n478), .A2(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g607(.A(KEYINPUT116), .B(G1384), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(KEYINPUT45), .B1(new_n505), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1032), .A2(new_n1035), .ZN(new_n1036));
  XNOR2_X1  g611(.A(new_n723), .B(G2067), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1036), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  XNOR2_X1  g614(.A(new_n1039), .B(KEYINPUT117), .ZN(new_n1040));
  XNOR2_X1  g615(.A(new_n753), .B(G1996), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1040), .B1(new_n1038), .B2(new_n1041), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n846), .A2(new_n848), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(G2067), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n724), .A2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1036), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1047));
  AND2_X1   g622(.A1(new_n846), .A2(new_n848), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1038), .B1(new_n1048), .B2(new_n1043), .ZN(new_n1049));
  NOR3_X1   g624(.A1(new_n1036), .A2(G1986), .A3(G290), .ZN(new_n1050));
  XOR2_X1   g625(.A(new_n1050), .B(KEYINPUT48), .Z(new_n1051));
  AND3_X1   g626(.A1(new_n1042), .A2(new_n1049), .A3(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1038), .B1(new_n1037), .B2(new_n753), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1036), .A2(G1996), .ZN(new_n1054));
  XOR2_X1   g629(.A(new_n1054), .B(KEYINPUT46), .Z(new_n1055));
  NAND2_X1  g630(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1056));
  XOR2_X1   g631(.A(new_n1056), .B(KEYINPUT47), .Z(new_n1057));
  NOR3_X1   g632(.A1(new_n1047), .A2(new_n1052), .A3(new_n1057), .ZN(new_n1058));
  XNOR2_X1  g633(.A(G290), .B(new_n832), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1042), .B(new_n1049), .C1(new_n1036), .C2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(G8), .ZN(new_n1061));
  AOI21_X1  g636(.A(KEYINPUT65), .B1(new_n476), .B2(G2105), .ZN(new_n1062));
  AOI211_X1 g637(.A(new_n460), .B(new_n462), .C1(new_n474), .C2(new_n475), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1064), .A2(G40), .A3(new_n473), .A4(new_n459), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT50), .ZN(new_n1066));
  INV_X1    g641(.A(G1384), .ZN(new_n1067));
  INV_X1    g642(.A(new_n496), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1068), .B1(new_n457), .B2(G126), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n500), .B1(new_n1069), .B2(new_n462), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n503), .A2(new_n504), .ZN(new_n1071));
  OAI211_X1 g646(.A(new_n1066), .B(new_n1067), .C1(new_n1070), .C2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(KEYINPUT118), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT118), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n505), .A2(new_n1074), .A3(new_n1066), .A4(new_n1067), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1065), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1076));
  AND2_X1   g651(.A1(new_n503), .A2(new_n504), .ZN(new_n1077));
  AOI22_X1  g652(.A1(new_n497), .A2(G2105), .B1(G102), .B2(new_n499), .ZN(new_n1078));
  AOI21_X1  g653(.A(G1384), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(KEYINPUT119), .B1(new_n1079), .B2(new_n1066), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1067), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT119), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1081), .A2(new_n1082), .A3(KEYINPUT50), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1080), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(G2090), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1076), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT45), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1081), .A2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n505), .A2(KEYINPUT45), .A3(new_n1034), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1032), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(new_n816), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1061), .B1(new_n1086), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT55), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1093), .B1(G303), .B2(G8), .ZN(new_n1094));
  AOI211_X1 g669(.A(KEYINPUT55), .B(new_n1061), .C1(new_n590), .C2(new_n591), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1092), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(G1976), .B1(new_n599), .B2(new_n601), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n593), .A2(new_n596), .A3(G1976), .A4(new_n597), .ZN(new_n1100));
  OAI211_X1 g675(.A(G8), .B(new_n1100), .C1(new_n1065), .C2(new_n1081), .ZN(new_n1101));
  NOR3_X1   g676(.A1(new_n1099), .A2(new_n1101), .A3(KEYINPUT52), .ZN(new_n1102));
  OAI21_X1  g677(.A(G8), .B1(new_n1065), .B2(new_n1081), .ZN(new_n1103));
  OAI211_X1 g678(.A(G61), .B(new_n509), .C1(new_n512), .C2(new_n513), .ZN(new_n1104));
  NAND2_X1  g679(.A1(G73), .A2(G543), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  AOI22_X1  g681(.A1(new_n1106), .A2(G651), .B1(G48), .B2(new_n519), .ZN(new_n1107));
  INV_X1    g682(.A(G1981), .ZN(new_n1108));
  AND3_X1   g683(.A1(new_n1107), .A2(new_n1108), .A3(new_n603), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1108), .B1(new_n1107), .B2(new_n603), .ZN(new_n1110));
  OAI211_X1 g685(.A(KEYINPUT120), .B(KEYINPUT49), .C1(new_n1109), .C2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g686(.A(G1981), .B1(new_n604), .B2(new_n607), .ZN(new_n1112));
  NAND2_X1  g687(.A1(KEYINPUT120), .A2(KEYINPUT49), .ZN(new_n1113));
  OR2_X1    g688(.A1(KEYINPUT120), .A2(KEYINPUT49), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1107), .A2(new_n1108), .A3(new_n603), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1112), .A2(new_n1113), .A3(new_n1114), .A4(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1103), .B1(new_n1111), .B2(new_n1116), .ZN(new_n1117));
  AND2_X1   g692(.A1(new_n1101), .A2(KEYINPUT52), .ZN(new_n1118));
  NOR3_X1   g693(.A1(new_n1102), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1098), .A2(new_n1119), .ZN(new_n1120));
  OR2_X1    g695(.A1(G288), .A2(G1976), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1111), .A2(new_n1116), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1115), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1032), .A2(new_n1079), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1123), .A2(G8), .A3(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1120), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1076), .A2(new_n1084), .A3(new_n771), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1079), .A2(KEYINPUT45), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1032), .A2(new_n1088), .A3(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(new_n785), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1128), .A2(G168), .A3(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1132), .A2(G8), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(KEYINPUT51), .ZN(new_n1134));
  AOI21_X1  g709(.A(G168), .B1(new_n1128), .B2(new_n1131), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT51), .ZN(new_n1136));
  OAI211_X1 g711(.A(G8), .B(new_n1132), .C1(new_n1135), .C2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT62), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1134), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1081), .A2(KEYINPUT50), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(new_n1072), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1141), .A2(new_n1065), .ZN(new_n1142));
  AOI22_X1  g717(.A1(new_n1142), .A2(new_n1085), .B1(new_n1090), .B2(new_n816), .ZN(new_n1143));
  OAI22_X1  g718(.A1(new_n1143), .A2(new_n1061), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1144));
  AND3_X1   g719(.A1(new_n1119), .A2(new_n1097), .A3(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1076), .A2(new_n1084), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT53), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1032), .A2(new_n781), .A3(new_n1088), .A4(new_n1089), .ZN(new_n1148));
  AOI22_X1  g723(.A1(new_n1146), .A2(new_n742), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1147), .A2(G2078), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1032), .A2(new_n1088), .A3(new_n1129), .A4(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(G301), .B1(new_n1149), .B2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1139), .A2(new_n1145), .A3(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1138), .B1(new_n1134), .B2(new_n1137), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1127), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1133), .A2(G286), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1145), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT63), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  AND2_X1   g734(.A1(new_n1092), .A2(KEYINPUT121), .ZN(new_n1160));
  OR2_X1    g735(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1161), .B1(new_n1092), .B2(KEYINPUT121), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1119), .B1(new_n1160), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1163), .A2(KEYINPUT122), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT122), .ZN(new_n1165));
  OAI211_X1 g740(.A(new_n1165), .B(new_n1119), .C1(new_n1160), .C2(new_n1162), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1098), .A2(new_n1158), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1164), .A2(new_n1156), .A3(new_n1166), .A4(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1155), .B1(new_n1159), .B2(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT54), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1171), .A2(new_n1032), .ZN(new_n1172));
  AOI211_X1 g747(.A(KEYINPUT119), .B(new_n1066), .C1(new_n505), .C2(new_n1067), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1082), .B1(new_n1081), .B2(KEYINPUT50), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n742), .B1(new_n1172), .B2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n476), .A2(G2105), .ZN(new_n1177));
  NAND4_X1  g752(.A1(new_n1089), .A2(G40), .A3(new_n1177), .A4(new_n1150), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n459), .A2(new_n473), .ZN(new_n1179));
  OR3_X1    g754(.A1(new_n1178), .A2(new_n1179), .A3(new_n1035), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1148), .A2(new_n1147), .ZN(new_n1181));
  AND4_X1   g756(.A1(G301), .A2(new_n1176), .A3(new_n1180), .A4(new_n1181), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1170), .B1(new_n1152), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1134), .A2(new_n1137), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1149), .A2(G301), .A3(new_n1151), .ZN(new_n1185));
  AND3_X1   g760(.A1(new_n1176), .A2(new_n1180), .A3(new_n1181), .ZN(new_n1186));
  OAI211_X1 g761(.A(new_n1185), .B(KEYINPUT54), .C1(new_n1186), .C2(G301), .ZN(new_n1187));
  NAND4_X1  g762(.A1(new_n1183), .A2(new_n1145), .A3(new_n1184), .A4(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1188), .A2(KEYINPUT126), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1176), .A2(new_n1151), .A3(new_n1181), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1190), .A2(G171), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1149), .A2(G301), .A3(new_n1180), .ZN(new_n1192));
  AOI21_X1  g767(.A(KEYINPUT54), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1119), .A2(new_n1097), .A3(new_n1144), .ZN(new_n1194));
  NOR2_X1   g769(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g770(.A(KEYINPUT126), .ZN(new_n1196));
  NAND4_X1  g771(.A1(new_n1195), .A2(new_n1196), .A3(new_n1184), .A4(new_n1187), .ZN(new_n1197));
  INV_X1    g772(.A(G1956), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1198), .B1(new_n1141), .B2(new_n1065), .ZN(new_n1199));
  INV_X1    g774(.A(KEYINPUT57), .ZN(new_n1200));
  OAI21_X1  g775(.A(new_n1200), .B1(new_n573), .B2(new_n575), .ZN(new_n1201));
  NAND4_X1  g776(.A1(new_n581), .A2(KEYINPUT57), .A3(new_n574), .A4(new_n568), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  XNOR2_X1  g778(.A(KEYINPUT56), .B(G2072), .ZN(new_n1204));
  NAND4_X1  g779(.A1(new_n1032), .A2(new_n1088), .A3(new_n1089), .A4(new_n1204), .ZN(new_n1205));
  NAND3_X1  g780(.A1(new_n1199), .A2(new_n1203), .A3(new_n1205), .ZN(new_n1206));
  AOI21_X1  g781(.A(new_n1203), .B1(new_n1199), .B2(new_n1205), .ZN(new_n1207));
  INV_X1    g782(.A(KEYINPUT125), .ZN(new_n1208));
  OAI21_X1  g783(.A(new_n1206), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  NAND4_X1  g784(.A1(new_n1199), .A2(KEYINPUT125), .A3(new_n1203), .A4(new_n1205), .ZN(new_n1210));
  NAND3_X1  g785(.A1(new_n1209), .A2(KEYINPUT61), .A3(new_n1210), .ZN(new_n1211));
  AOI21_X1  g786(.A(G1348), .B1(new_n1076), .B2(new_n1084), .ZN(new_n1212));
  INV_X1    g787(.A(new_n1212), .ZN(new_n1213));
  NOR2_X1   g788(.A1(new_n1124), .A2(G2067), .ZN(new_n1214));
  INV_X1    g789(.A(new_n1214), .ZN(new_n1215));
  NAND3_X1  g790(.A1(new_n1213), .A2(KEYINPUT60), .A3(new_n1215), .ZN(new_n1216));
  INV_X1    g791(.A(KEYINPUT60), .ZN(new_n1217));
  OAI21_X1  g792(.A(new_n1217), .B1(new_n1212), .B2(new_n1214), .ZN(new_n1218));
  NAND3_X1  g793(.A1(new_n1216), .A2(new_n635), .A3(new_n1218), .ZN(new_n1219));
  NAND4_X1  g794(.A1(new_n1213), .A2(KEYINPUT60), .A3(new_n624), .A4(new_n1215), .ZN(new_n1220));
  XOR2_X1   g795(.A(KEYINPUT58), .B(G1341), .Z(new_n1221));
  NAND2_X1  g796(.A1(new_n1124), .A2(new_n1221), .ZN(new_n1222));
  OAI21_X1  g797(.A(new_n1222), .B1(G1996), .B2(new_n1090), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1223), .A2(new_n558), .ZN(new_n1224));
  NOR2_X1   g799(.A1(KEYINPUT124), .A2(KEYINPUT59), .ZN(new_n1225));
  NAND2_X1  g800(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  NAND4_X1  g801(.A1(new_n1211), .A2(new_n1219), .A3(new_n1220), .A4(new_n1226), .ZN(new_n1227));
  INV_X1    g802(.A(new_n1206), .ZN(new_n1228));
  OR2_X1    g803(.A1(new_n1228), .A2(KEYINPUT123), .ZN(new_n1229));
  NAND2_X1  g804(.A1(new_n1228), .A2(KEYINPUT123), .ZN(new_n1230));
  AOI21_X1  g805(.A(KEYINPUT61), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  AND2_X1   g806(.A1(KEYINPUT124), .A2(KEYINPUT59), .ZN(new_n1232));
  NOR3_X1   g807(.A1(new_n1224), .A2(new_n1225), .A3(new_n1232), .ZN(new_n1233));
  NOR3_X1   g808(.A1(new_n1227), .A2(new_n1231), .A3(new_n1233), .ZN(new_n1234));
  NAND2_X1  g809(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1235));
  OAI21_X1  g810(.A(new_n635), .B1(new_n1212), .B2(new_n1214), .ZN(new_n1236));
  INV_X1    g811(.A(new_n1207), .ZN(new_n1237));
  AOI21_X1  g812(.A(new_n1235), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  OAI211_X1 g813(.A(new_n1189), .B(new_n1197), .C1(new_n1234), .C2(new_n1238), .ZN(new_n1239));
  AOI211_X1 g814(.A(KEYINPUT127), .B(new_n1060), .C1(new_n1169), .C2(new_n1239), .ZN(new_n1240));
  INV_X1    g815(.A(KEYINPUT127), .ZN(new_n1241));
  INV_X1    g816(.A(new_n1155), .ZN(new_n1242));
  NAND2_X1  g817(.A1(new_n1168), .A2(new_n1159), .ZN(new_n1243));
  NAND2_X1  g818(.A1(new_n1189), .A2(new_n1197), .ZN(new_n1244));
  NOR2_X1   g819(.A1(new_n1227), .A2(new_n1231), .ZN(new_n1245));
  INV_X1    g820(.A(new_n1233), .ZN(new_n1246));
  AOI21_X1  g821(.A(new_n1238), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  OAI211_X1 g822(.A(new_n1242), .B(new_n1243), .C1(new_n1244), .C2(new_n1247), .ZN(new_n1248));
  INV_X1    g823(.A(new_n1060), .ZN(new_n1249));
  AOI21_X1  g824(.A(new_n1241), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  OAI21_X1  g825(.A(new_n1058), .B1(new_n1240), .B2(new_n1250), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g826(.A(G319), .ZN(new_n1253));
  NOR2_X1   g827(.A1(G401), .A2(new_n1253), .ZN(new_n1254));
  NOR2_X1   g828(.A1(G227), .A2(G229), .ZN(new_n1255));
  AND4_X1   g829(.A1(new_n929), .A2(new_n1016), .A3(new_n1254), .A4(new_n1255), .ZN(G308));
  NAND4_X1  g830(.A1(new_n1016), .A2(new_n929), .A3(new_n1254), .A4(new_n1255), .ZN(G225));
endmodule


