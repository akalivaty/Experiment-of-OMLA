//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 0 1 1 0 1 0 1 1 1 1 0 1 0 1 1 0 1 1 1 0 1 1 1 1 0 0 1 1 0 0 1 1 0 1 0 0 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n749,
    new_n750, new_n751, new_n752, new_n754, new_n755, new_n756, new_n757,
    new_n759, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n944, new_n945, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985;
  INV_X1    g000(.A(KEYINPUT34), .ZN(new_n202));
  OAI21_X1  g001(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n203));
  AND2_X1   g002(.A1(G183gat), .A2(G190gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G169gat), .A2(G176gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(G183gat), .A2(G190gat), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n206), .B1(new_n207), .B2(KEYINPUT24), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n205), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT23), .ZN(new_n210));
  INV_X1    g009(.A(G169gat), .ZN(new_n211));
  INV_X1    g010(.A(G176gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n210), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  OAI21_X1  g012(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  AOI21_X1  g014(.A(KEYINPUT25), .B1(new_n209), .B2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT24), .ZN(new_n217));
  AOI22_X1  g016(.A1(new_n204), .A2(new_n217), .B1(G169gat), .B2(G176gat), .ZN(new_n218));
  OR2_X1    g017(.A1(G183gat), .A2(G190gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n219), .A2(KEYINPUT24), .A3(new_n207), .ZN(new_n220));
  AND4_X1   g019(.A1(KEYINPUT25), .A2(new_n218), .A3(new_n215), .A4(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(KEYINPUT64), .B1(new_n216), .B2(new_n221), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n218), .A2(new_n215), .A3(new_n220), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT25), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT64), .ZN(new_n226));
  NAND4_X1  g025(.A1(new_n218), .A2(new_n215), .A3(new_n220), .A4(KEYINPUT25), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  OAI21_X1  g027(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n229));
  OR2_X1    g028(.A1(new_n229), .A2(KEYINPUT66), .ZN(new_n230));
  AOI22_X1  g029(.A1(new_n229), .A2(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n231));
  NOR4_X1   g030(.A1(KEYINPUT67), .A2(KEYINPUT26), .A3(G169gat), .A4(G176gat), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT67), .ZN(new_n233));
  NOR2_X1   g032(.A1(G169gat), .A2(G176gat), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT26), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n233), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  OAI211_X1 g035(.A(new_n230), .B(new_n231), .C1(new_n232), .C2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT27), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n238), .A2(G183gat), .ZN(new_n239));
  INV_X1    g038(.A(G183gat), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n240), .A2(KEYINPUT27), .ZN(new_n241));
  OAI21_X1  g040(.A(KEYINPUT65), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n240), .A2(KEYINPUT27), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT65), .ZN(new_n244));
  AOI21_X1  g043(.A(G190gat), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  AOI21_X1  g044(.A(KEYINPUT28), .B1(new_n242), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n238), .A2(G183gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n243), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT28), .ZN(new_n249));
  NOR3_X1   g048(.A1(new_n248), .A2(new_n249), .A3(G190gat), .ZN(new_n250));
  OAI211_X1 g049(.A(new_n237), .B(new_n207), .C1(new_n246), .C2(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n222), .A2(new_n228), .A3(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(G127gat), .B(G134gat), .ZN(new_n253));
  OR2_X1    g052(.A1(new_n253), .A2(KEYINPUT69), .ZN(new_n254));
  XNOR2_X1  g053(.A(G113gat), .B(G120gat), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n253), .A2(KEYINPUT69), .ZN(new_n257));
  XOR2_X1   g056(.A(KEYINPUT70), .B(KEYINPUT1), .Z(new_n258));
  NAND4_X1  g057(.A1(new_n254), .A2(new_n256), .A3(new_n257), .A4(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(G127gat), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n260), .A2(KEYINPUT68), .A3(G134gat), .ZN(new_n261));
  INV_X1    g060(.A(new_n253), .ZN(new_n262));
  OAI221_X1 g061(.A(new_n261), .B1(new_n255), .B2(KEYINPUT1), .C1(new_n262), .C2(KEYINPUT68), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n259), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n252), .A2(new_n265), .ZN(new_n266));
  NAND4_X1  g065(.A1(new_n222), .A2(new_n264), .A3(new_n251), .A4(new_n228), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(G227gat), .A2(G233gat), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n202), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT71), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n268), .A2(new_n202), .A3(new_n269), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n270), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(new_n269), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n266), .A2(new_n274), .A3(new_n267), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT33), .ZN(new_n276));
  XOR2_X1   g075(.A(G15gat), .B(G43gat), .Z(new_n277));
  XNOR2_X1  g076(.A(G71gat), .B(G99gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n277), .B(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  OAI211_X1 g079(.A(new_n275), .B(KEYINPUT32), .C1(new_n276), .C2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n275), .A2(KEYINPUT32), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n275), .A2(new_n276), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n282), .A2(new_n283), .A3(new_n279), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n268), .A2(KEYINPUT71), .A3(new_n202), .A4(new_n269), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n273), .A2(new_n281), .A3(new_n284), .A4(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n284), .A2(new_n281), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n272), .A2(new_n271), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n268), .A2(new_n269), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(KEYINPUT34), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n288), .A2(new_n285), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n287), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT80), .ZN(new_n293));
  NAND2_X1  g092(.A1(G228gat), .A2(G233gat), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  AND2_X1   g094(.A1(G155gat), .A2(G162gat), .ZN(new_n296));
  NOR2_X1   g095(.A1(G155gat), .A2(G162gat), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(G141gat), .B(G148gat), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT2), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n300), .B1(G155gat), .B2(G162gat), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n298), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(G141gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(G148gat), .ZN(new_n304));
  INV_X1    g103(.A(G148gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(G141gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(G155gat), .B(G162gat), .ZN(new_n308));
  INV_X1    g107(.A(G155gat), .ZN(new_n309));
  INV_X1    g108(.A(G162gat), .ZN(new_n310));
  OAI21_X1  g109(.A(KEYINPUT2), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n307), .A2(new_n308), .A3(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT3), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n302), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT29), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(G211gat), .A2(G218gat), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  NOR2_X1   g118(.A1(G211gat), .A2(G218gat), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT73), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT22), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n318), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(G197gat), .ZN(new_n325));
  INV_X1    g124(.A(G204gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(G197gat), .A2(G204gat), .ZN(new_n328));
  AOI22_X1  g127(.A1(new_n322), .A2(new_n324), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  AOI21_X1  g128(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(KEYINPUT73), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n321), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT74), .ZN(new_n333));
  AND2_X1   g132(.A1(G197gat), .A2(G204gat), .ZN(new_n334));
  NOR2_X1   g133(.A1(G197gat), .A2(G204gat), .ZN(new_n335));
  OAI22_X1  g134(.A1(new_n330), .A2(KEYINPUT73), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n324), .A2(new_n322), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n333), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  AOI22_X1  g137(.A1(new_n332), .A2(new_n333), .B1(new_n338), .B2(new_n321), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n295), .B1(new_n317), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n302), .A2(new_n312), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  OR2_X1    g141(.A1(new_n319), .A2(new_n320), .ZN(new_n343));
  OAI211_X1 g142(.A(new_n333), .B(new_n343), .C1(new_n336), .C2(new_n337), .ZN(new_n344));
  AOI21_X1  g143(.A(KEYINPUT74), .B1(new_n329), .B2(new_n331), .ZN(new_n345));
  OAI211_X1 g144(.A(new_n315), .B(new_n344), .C1(new_n345), .C2(new_n343), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n342), .B1(new_n346), .B2(new_n313), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n340), .A2(new_n347), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n343), .B1(new_n336), .B2(new_n337), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n324), .A2(new_n322), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n327), .A2(new_n328), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n350), .A2(new_n321), .A3(new_n331), .A4(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n349), .A2(new_n315), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(new_n313), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(new_n341), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n338), .A2(new_n321), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(new_n344), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(new_n316), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n295), .B1(new_n355), .B2(new_n358), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n293), .B1(new_n348), .B2(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n342), .B1(new_n353), .B2(new_n313), .ZN(new_n361));
  AOI22_X1  g160(.A1(new_n356), .A2(new_n344), .B1(new_n314), .B2(new_n315), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n294), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  OAI211_X1 g162(.A(new_n363), .B(KEYINPUT80), .C1(new_n347), .C2(new_n340), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n360), .A2(G22gat), .A3(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n348), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT81), .ZN(new_n367));
  INV_X1    g166(.A(G22gat), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n366), .A2(new_n367), .A3(new_n368), .A4(new_n363), .ZN(new_n369));
  XNOR2_X1  g168(.A(G78gat), .B(G106gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(new_n370), .B(KEYINPUT31), .ZN(new_n371));
  INV_X1    g170(.A(G50gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n371), .B(new_n372), .ZN(new_n373));
  OAI211_X1 g172(.A(new_n363), .B(new_n368), .C1(new_n347), .C2(new_n340), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n373), .B1(new_n374), .B2(KEYINPUT81), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n365), .A2(new_n369), .A3(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n368), .B1(new_n366), .B2(new_n363), .ZN(new_n377));
  INV_X1    g176(.A(new_n374), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n373), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n286), .A2(new_n292), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(KEYINPUT85), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT85), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n286), .A2(new_n292), .A3(new_n380), .A4(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n225), .A2(new_n227), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n251), .A2(new_n386), .ZN(new_n387));
  AND2_X1   g186(.A1(G226gat), .A2(G233gat), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n388), .B1(new_n252), .B2(new_n315), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n389), .B1(new_n390), .B2(KEYINPUT75), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT75), .ZN(new_n392));
  AOI211_X1 g191(.A(new_n392), .B(new_n388), .C1(new_n252), .C2(new_n315), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n357), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n388), .A2(KEYINPUT29), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n387), .A2(new_n395), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n222), .A2(new_n388), .A3(new_n251), .A4(new_n228), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT76), .B1(new_n398), .B2(new_n339), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT76), .ZN(new_n400));
  AOI211_X1 g199(.A(new_n400), .B(new_n357), .C1(new_n396), .C2(new_n397), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n394), .A2(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(G8gat), .B(G36gat), .ZN(new_n404));
  XNOR2_X1  g203(.A(new_n404), .B(G64gat), .ZN(new_n405));
  INV_X1    g204(.A(G92gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n405), .B(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n403), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(KEYINPUT77), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT77), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n403), .A2(new_n411), .A3(new_n408), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n394), .A2(new_n402), .A3(new_n407), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT30), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND4_X1  g215(.A1(new_n394), .A2(new_n402), .A3(KEYINPUT30), .A4(new_n407), .ZN(new_n417));
  AND2_X1   g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  XOR2_X1   g217(.A(KEYINPUT79), .B(KEYINPUT0), .Z(new_n419));
  XNOR2_X1  g218(.A(G1gat), .B(G29gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n419), .B(new_n420), .ZN(new_n421));
  XNOR2_X1  g220(.A(G57gat), .B(G85gat), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n421), .B(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n342), .A2(new_n259), .A3(new_n263), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(KEYINPUT4), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT4), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n342), .A2(new_n259), .A3(new_n263), .A4(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(G225gat), .A2(G233gat), .ZN(new_n430));
  AOI22_X1  g229(.A1(new_n259), .A2(new_n263), .B1(new_n341), .B2(KEYINPUT3), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(new_n314), .ZN(new_n432));
  XOR2_X1   g231(.A(KEYINPUT78), .B(KEYINPUT5), .Z(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n429), .A2(new_n430), .A3(new_n432), .A4(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n264), .A2(new_n341), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(new_n425), .ZN(new_n437));
  INV_X1    g236(.A(new_n430), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n435), .A2(new_n439), .ZN(new_n440));
  AOI22_X1  g239(.A1(new_n426), .A2(new_n428), .B1(new_n314), .B2(new_n431), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n434), .B1(new_n441), .B2(new_n430), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n424), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT6), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n429), .A2(new_n430), .A3(new_n432), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(new_n433), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n446), .A2(new_n423), .A3(new_n439), .A4(new_n435), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n443), .A2(new_n444), .A3(new_n447), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n440), .A2(new_n442), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n449), .A2(KEYINPUT6), .A3(new_n423), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n413), .A2(new_n418), .A3(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(KEYINPUT35), .B1(new_n385), .B2(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n411), .B1(new_n403), .B2(new_n408), .ZN(new_n454));
  AOI211_X1 g253(.A(KEYINPUT77), .B(new_n407), .C1(new_n394), .C2(new_n402), .ZN(new_n455));
  OAI211_X1 g254(.A(new_n416), .B(new_n417), .C1(new_n454), .C2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n451), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT35), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n380), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT72), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n286), .A2(new_n292), .A3(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n287), .A2(new_n291), .A3(KEYINPUT72), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n460), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n458), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n453), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n429), .A2(new_n432), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT39), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n467), .A2(new_n468), .A3(new_n438), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT82), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n470), .B1(new_n437), .B2(new_n438), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n436), .A2(KEYINPUT82), .A3(new_n430), .A4(new_n425), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n471), .A2(KEYINPUT39), .A3(new_n472), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n441), .A2(new_n430), .ZN(new_n474));
  OAI211_X1 g273(.A(new_n469), .B(new_n424), .C1(new_n473), .C2(new_n474), .ZN(new_n475));
  XOR2_X1   g274(.A(KEYINPUT83), .B(KEYINPUT40), .Z(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(new_n447), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT84), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT40), .ZN(new_n480));
  OR3_X1    g279(.A1(new_n475), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n479), .B1(new_n475), .B2(new_n480), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n478), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n456), .A2(new_n483), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n339), .B1(new_n391), .B2(new_n393), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT37), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n486), .B1(new_n398), .B2(new_n357), .ZN(new_n487));
  AOI21_X1  g286(.A(KEYINPUT38), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  OAI211_X1 g287(.A(new_n488), .B(new_n408), .C1(KEYINPUT37), .C2(new_n403), .ZN(new_n489));
  AND3_X1   g288(.A1(new_n448), .A2(new_n414), .A3(new_n450), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n486), .B1(new_n394), .B2(new_n402), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n408), .A2(KEYINPUT37), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n491), .B1(new_n409), .B2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT38), .ZN(new_n494));
  OAI211_X1 g293(.A(new_n489), .B(new_n490), .C1(new_n493), .C2(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n484), .A2(new_n495), .A3(new_n380), .ZN(new_n496));
  INV_X1    g295(.A(new_n380), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n497), .B1(new_n456), .B2(new_n457), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT36), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n462), .A2(new_n499), .A3(new_n463), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n286), .A2(new_n292), .A3(KEYINPUT36), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n496), .A2(new_n498), .A3(new_n502), .ZN(new_n503));
  AND3_X1   g302(.A1(new_n466), .A2(KEYINPUT86), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(KEYINPUT86), .B1(new_n466), .B2(new_n503), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(G15gat), .B(G22gat), .ZN(new_n507));
  INV_X1    g306(.A(G1gat), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n507), .A2(KEYINPUT16), .A3(new_n508), .ZN(new_n509));
  OAI221_X1 g308(.A(new_n509), .B1(KEYINPUT89), .B2(G8gat), .C1(new_n508), .C2(new_n507), .ZN(new_n510));
  NAND2_X1  g309(.A1(KEYINPUT89), .A2(G8gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n510), .B(new_n511), .ZN(new_n512));
  XOR2_X1   g311(.A(G71gat), .B(G78gat), .Z(new_n513));
  INV_X1    g312(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(G71gat), .A2(G78gat), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT9), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  XOR2_X1   g316(.A(G57gat), .B(G64gat), .Z(new_n518));
  NAND3_X1  g317(.A1(new_n514), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n517), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(new_n513), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n512), .B1(KEYINPUT21), .B2(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n524), .B(new_n240), .ZN(new_n525));
  XNOR2_X1  g324(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n526));
  NAND2_X1  g325(.A1(G231gat), .A2(G233gat), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n526), .B(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n525), .B(new_n528), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n523), .A2(KEYINPUT21), .ZN(new_n530));
  XNOR2_X1  g329(.A(G127gat), .B(G155gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n530), .B(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n532), .B(G211gat), .ZN(new_n533));
  OR2_X1    g332(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n529), .A2(new_n533), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AND2_X1   g335(.A1(G232gat), .A2(G233gat), .ZN(new_n537));
  OR2_X1    g336(.A1(new_n537), .A2(KEYINPUT41), .ZN(new_n538));
  XNOR2_X1  g337(.A(G134gat), .B(G162gat), .ZN(new_n539));
  XOR2_X1   g338(.A(new_n538), .B(new_n539), .Z(new_n540));
  OR2_X1    g339(.A1(new_n372), .A2(G43gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n372), .A2(G43gat), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n541), .A2(KEYINPUT15), .A3(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(KEYINPUT87), .B(G43gat), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(new_n372), .ZN(new_n545));
  AOI21_X1  g344(.A(KEYINPUT15), .B1(new_n545), .B2(new_n541), .ZN(new_n546));
  INV_X1    g345(.A(G29gat), .ZN(new_n547));
  INV_X1    g346(.A(G36gat), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n547), .A2(new_n548), .A3(KEYINPUT14), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT14), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n550), .B1(G29gat), .B2(G36gat), .ZN(new_n551));
  OAI211_X1 g350(.A(new_n549), .B(new_n551), .C1(new_n547), .C2(new_n548), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n543), .B1(new_n546), .B2(new_n552), .ZN(new_n553));
  OR2_X1    g352(.A1(new_n552), .A2(new_n543), .ZN(new_n554));
  AND2_X1   g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT88), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n555), .A2(new_n556), .A3(KEYINPUT17), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT17), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n553), .A2(new_n554), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n558), .B1(new_n559), .B2(KEYINPUT88), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(G85gat), .A2(G92gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(KEYINPUT7), .ZN(new_n563));
  NAND2_X1  g362(.A1(G99gat), .A2(G106gat), .ZN(new_n564));
  INV_X1    g363(.A(G85gat), .ZN(new_n565));
  AOI22_X1  g364(.A1(KEYINPUT8), .A2(new_n564), .B1(new_n565), .B2(new_n406), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  XOR2_X1   g366(.A(G99gat), .B(G106gat), .Z(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n567), .B(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(KEYINPUT92), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT92), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n567), .A2(new_n568), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n567), .A2(new_n568), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n572), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n571), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n561), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(G190gat), .B(G218gat), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(KEYINPUT93), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n537), .A2(KEYINPUT41), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n583), .B1(new_n577), .B2(new_n555), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n579), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n580), .A2(KEYINPUT93), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  OAI211_X1 g386(.A(new_n579), .B(new_n584), .C1(KEYINPUT93), .C2(new_n580), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n540), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n587), .A2(new_n540), .A3(new_n588), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n536), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(G230gat), .A2(G233gat), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  NOR3_X1   g394(.A1(new_n574), .A2(new_n572), .A3(new_n575), .ZN(new_n596));
  AND2_X1   g395(.A1(new_n563), .A2(new_n566), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(new_n569), .ZN(new_n598));
  AOI21_X1  g397(.A(KEYINPUT92), .B1(new_n598), .B2(new_n573), .ZN(new_n599));
  OAI211_X1 g398(.A(KEYINPUT10), .B(new_n523), .C1(new_n596), .C2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n570), .A2(new_n523), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT10), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n522), .B1(new_n574), .B2(new_n575), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n595), .B1(new_n600), .B2(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n594), .B1(new_n601), .B2(new_n603), .ZN(new_n606));
  XNOR2_X1  g405(.A(G120gat), .B(G148gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(G176gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(new_n326), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  OR3_X1    g409(.A1(new_n605), .A2(new_n606), .A3(new_n610), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n610), .B1(new_n605), .B2(new_n606), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(G113gat), .B(G141gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(KEYINPUT11), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(new_n211), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(new_n325), .ZN(new_n617));
  XOR2_X1   g416(.A(new_n617), .B(KEYINPUT12), .Z(new_n618));
  INV_X1    g417(.A(new_n512), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n561), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(G229gat), .A2(G233gat), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n512), .A2(new_n555), .ZN(new_n622));
  NAND4_X1  g421(.A1(new_n620), .A2(KEYINPUT18), .A3(new_n621), .A4(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(KEYINPUT90), .ZN(new_n624));
  INV_X1    g423(.A(new_n622), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n625), .B1(new_n619), .B2(new_n561), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT90), .ZN(new_n627));
  NAND4_X1  g426(.A1(new_n626), .A2(new_n627), .A3(KEYINPUT18), .A4(new_n621), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n624), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n626), .A2(new_n621), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT18), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n512), .B(new_n555), .ZN(new_n632));
  XOR2_X1   g431(.A(new_n621), .B(KEYINPUT13), .Z(new_n633));
  AOI22_X1  g432(.A1(new_n630), .A2(new_n631), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n618), .B1(new_n629), .B2(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n629), .A2(new_n634), .A3(new_n618), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(KEYINPUT91), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT91), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n629), .A2(new_n634), .A3(new_n638), .A4(new_n618), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n635), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  NOR3_X1   g439(.A1(new_n593), .A2(new_n613), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n506), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n642), .A2(new_n451), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(new_n508), .ZN(G1324gat));
  NAND2_X1  g443(.A1(new_n416), .A2(new_n417), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n645), .B1(new_n410), .B2(new_n412), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n642), .A2(new_n646), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n647), .A2(KEYINPUT42), .ZN(new_n648));
  NOR2_X1   g447(.A1(KEYINPUT94), .A2(KEYINPUT42), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(KEYINPUT16), .ZN(new_n650));
  NOR3_X1   g449(.A1(new_n642), .A2(new_n646), .A3(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n648), .B1(G8gat), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n653), .B1(G8gat), .B2(new_n652), .ZN(G1325gat));
  INV_X1    g453(.A(KEYINPUT95), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n502), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n500), .A2(KEYINPUT95), .A3(new_n501), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(G15gat), .B1(new_n642), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n462), .A2(new_n463), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  OR2_X1    g461(.A1(new_n662), .A2(G15gat), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n660), .B1(new_n642), .B2(new_n663), .ZN(G1326gat));
  OR3_X1    g463(.A1(new_n642), .A2(KEYINPUT96), .A3(new_n380), .ZN(new_n665));
  OAI21_X1  g464(.A(KEYINPUT96), .B1(new_n642), .B2(new_n380), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  OR2_X1    g466(.A1(new_n667), .A2(KEYINPUT97), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(KEYINPUT97), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(KEYINPUT43), .B(G22gat), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n668), .A2(new_n671), .A3(new_n669), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(G1327gat));
  NOR3_X1   g474(.A1(new_n504), .A2(new_n505), .A3(new_n592), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n640), .A2(new_n536), .A3(new_n613), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NOR3_X1   g477(.A1(new_n678), .A2(G29gat), .A3(new_n451), .ZN(new_n679));
  XOR2_X1   g478(.A(new_n679), .B(KEYINPUT45), .Z(new_n680));
  INV_X1    g479(.A(KEYINPUT99), .ZN(new_n681));
  INV_X1    g480(.A(new_n591), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n681), .B1(new_n682), .B2(new_n589), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n590), .A2(KEYINPUT99), .A3(new_n591), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  NAND4_X1  g485(.A1(new_n656), .A2(new_n496), .A3(new_n498), .A4(new_n657), .ZN(new_n687));
  AOI211_X1 g486(.A(KEYINPUT44), .B(new_n686), .C1(new_n687), .C2(new_n466), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n689), .B1(new_n676), .B2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT100), .ZN(new_n692));
  XOR2_X1   g491(.A(new_n677), .B(KEYINPUT98), .Z(new_n693));
  NAND3_X1  g492(.A1(new_n691), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT86), .ZN(new_n695));
  AND3_X1   g494(.A1(new_n484), .A2(new_n495), .A3(new_n380), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n498), .A2(new_n502), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND4_X1  g497(.A1(new_n646), .A2(new_n451), .A3(new_n382), .A4(new_n384), .ZN(new_n699));
  AOI22_X1  g498(.A1(new_n699), .A2(KEYINPUT35), .B1(new_n458), .B2(new_n464), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n695), .B1(new_n698), .B2(new_n700), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n466), .A2(new_n503), .A3(KEYINPUT86), .ZN(new_n702));
  INV_X1    g501(.A(new_n592), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n701), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n688), .B1(new_n704), .B2(KEYINPUT44), .ZN(new_n705));
  INV_X1    g504(.A(new_n693), .ZN(new_n706));
  OAI21_X1  g505(.A(KEYINPUT100), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n694), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(KEYINPUT101), .B1(new_n708), .B2(new_n451), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(G29gat), .ZN(new_n710));
  NOR3_X1   g509(.A1(new_n708), .A2(KEYINPUT101), .A3(new_n451), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n680), .B1(new_n710), .B2(new_n711), .ZN(G1328gat));
  OAI21_X1  g511(.A(G36gat), .B1(new_n708), .B2(new_n646), .ZN(new_n713));
  NOR3_X1   g512(.A1(new_n678), .A2(G36gat), .A3(new_n646), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT46), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n713), .A2(new_n715), .ZN(G1329gat));
  OR2_X1    g515(.A1(new_n662), .A2(new_n544), .ZN(new_n717));
  OR2_X1    g516(.A1(new_n678), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT102), .ZN(new_n719));
  OR2_X1    g518(.A1(new_n719), .A2(KEYINPUT47), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n691), .A2(new_n693), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n721), .A2(new_n659), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n544), .A2(KEYINPUT47), .ZN(new_n723));
  OAI211_X1 g522(.A(new_n718), .B(new_n720), .C1(new_n722), .C2(new_n723), .ZN(new_n724));
  NOR3_X1   g523(.A1(new_n678), .A2(new_n719), .A3(new_n717), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n694), .A2(new_n707), .A3(new_n658), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n725), .B1(new_n726), .B2(new_n544), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n724), .B1(new_n727), .B2(KEYINPUT47), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT103), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  OAI211_X1 g529(.A(KEYINPUT103), .B(new_n724), .C1(new_n727), .C2(KEYINPUT47), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(G1330gat));
  OAI21_X1  g531(.A(G50gat), .B1(new_n721), .B2(new_n380), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT104), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n678), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n676), .A2(KEYINPUT104), .A3(new_n677), .ZN(new_n736));
  NAND4_X1  g535(.A1(new_n735), .A2(new_n372), .A3(new_n497), .A4(new_n736), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n733), .A2(KEYINPUT48), .A3(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(G50gat), .B1(new_n708), .B2(new_n380), .ZN(new_n739));
  AND2_X1   g538(.A1(new_n739), .A2(new_n737), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n738), .B1(new_n740), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g540(.A1(new_n687), .A2(new_n466), .ZN(new_n742));
  INV_X1    g541(.A(new_n640), .ZN(new_n743));
  INV_X1    g542(.A(new_n613), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n743), .A2(new_n593), .A3(new_n744), .ZN(new_n745));
  AND2_X1   g544(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(new_n457), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g547(.A(new_n646), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n746), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(KEYINPUT105), .ZN(new_n751));
  NOR2_X1   g550(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n751), .B(new_n752), .ZN(G1333gat));
  NAND3_X1  g552(.A1(new_n746), .A2(G71gat), .A3(new_n658), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(KEYINPUT106), .ZN(new_n755));
  AOI21_X1  g554(.A(G71gat), .B1(new_n746), .B2(new_n661), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  XOR2_X1   g556(.A(new_n757), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g557(.A1(new_n746), .A2(new_n497), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g559(.A1(new_n743), .A2(new_n536), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n742), .A2(new_n703), .A3(new_n761), .ZN(new_n762));
  XOR2_X1   g561(.A(new_n762), .B(KEYINPUT51), .Z(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(KEYINPUT107), .ZN(new_n764));
  NAND4_X1  g563(.A1(new_n764), .A2(new_n565), .A3(new_n457), .A4(new_n613), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n691), .A2(new_n613), .A3(new_n761), .ZN(new_n766));
  OAI21_X1  g565(.A(G85gat), .B1(new_n766), .B2(new_n451), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n765), .A2(new_n767), .ZN(G1336gat));
  OAI21_X1  g567(.A(G92gat), .B1(new_n766), .B2(new_n646), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n763), .A2(new_n613), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n456), .A2(new_n406), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n769), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(KEYINPUT52), .ZN(G1337gat));
  NOR3_X1   g572(.A1(new_n662), .A2(G99gat), .A3(new_n744), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n764), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(G99gat), .B1(new_n766), .B2(new_n659), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(G1338gat));
  NOR2_X1   g576(.A1(new_n766), .A2(new_n380), .ZN(new_n778));
  INV_X1    g577(.A(G106gat), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n770), .A2(G106gat), .A3(new_n380), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT108), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT109), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n782), .B1(new_n783), .B2(KEYINPUT53), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n780), .A2(new_n781), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n781), .A2(KEYINPUT108), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n786), .B(new_n783), .C1(new_n779), .C2(new_n778), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT53), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n785), .B1(new_n787), .B2(new_n788), .ZN(G1339gat));
  INV_X1    g588(.A(KEYINPUT114), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n637), .A2(new_n639), .ZN(new_n791));
  XNOR2_X1  g590(.A(KEYINPUT111), .B(KEYINPUT54), .ZN(new_n792));
  AND3_X1   g591(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n523), .A2(KEYINPUT10), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n794), .B1(new_n571), .B2(new_n576), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n594), .B(new_n792), .C1(new_n793), .C2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(new_n610), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n600), .A2(new_n595), .A3(new_n604), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(KEYINPUT110), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT110), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n600), .A2(new_n604), .A3(new_n800), .A4(new_n595), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT54), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n605), .A2(new_n803), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n797), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  AND3_X1   g604(.A1(new_n805), .A2(KEYINPUT112), .A3(KEYINPUT55), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n611), .B1(new_n805), .B2(KEYINPUT55), .ZN(new_n807));
  AOI21_X1  g606(.A(KEYINPUT112), .B1(new_n805), .B2(KEYINPUT55), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n806), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  OAI22_X1  g608(.A1(new_n626), .A2(new_n621), .B1(new_n632), .B2(new_n633), .ZN(new_n810));
  INV_X1    g609(.A(new_n617), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n791), .A2(new_n809), .A3(new_n685), .A4(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(KEYINPUT113), .ZN(new_n814));
  AOI22_X1  g613(.A1(new_n637), .A2(new_n639), .B1(new_n811), .B2(new_n810), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT113), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n815), .A2(new_n816), .A3(new_n685), .A4(new_n809), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n791), .A2(new_n613), .A3(new_n812), .ZN(new_n819));
  INV_X1    g618(.A(new_n809), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n819), .B1(new_n640), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(new_n686), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n536), .B1(new_n818), .B2(new_n822), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n640), .A2(new_n536), .A3(new_n592), .A4(new_n744), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n790), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  AOI22_X1  g625(.A1(new_n814), .A2(new_n817), .B1(new_n821), .B2(new_n686), .ZN(new_n827));
  OAI211_X1 g626(.A(KEYINPUT114), .B(new_n824), .C1(new_n827), .C2(new_n536), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n829), .A2(new_n451), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n385), .A2(new_n456), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(G113gat), .B1(new_n833), .B2(new_n743), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n456), .A2(new_n451), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n662), .A2(new_n497), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n826), .A2(new_n828), .A3(new_n835), .A4(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT115), .ZN(new_n838));
  OR2_X1    g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n837), .A2(new_n838), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n743), .A2(G113gat), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n834), .B1(new_n841), .B2(new_n842), .ZN(G1340gat));
  OR3_X1    g642(.A1(new_n832), .A2(G120gat), .A3(new_n744), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n839), .A2(new_n613), .A3(new_n840), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT116), .ZN(new_n846));
  AND3_X1   g645(.A1(new_n845), .A2(new_n846), .A3(G120gat), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n846), .B1(new_n845), .B2(G120gat), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n844), .B1(new_n847), .B2(new_n848), .ZN(G1341gat));
  INV_X1    g648(.A(new_n536), .ZN(new_n850));
  OR3_X1    g649(.A1(new_n832), .A2(KEYINPUT117), .A3(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(KEYINPUT117), .B1(new_n832), .B2(new_n850), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n851), .A2(new_n260), .A3(new_n852), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n841), .A2(G127gat), .A3(new_n536), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n853), .A2(new_n854), .ZN(G1342gat));
  NOR2_X1   g654(.A1(new_n592), .A2(G134gat), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(KEYINPUT56), .B1(new_n832), .B2(new_n857), .ZN(new_n858));
  OR3_X1    g657(.A1(new_n832), .A2(KEYINPUT56), .A3(new_n857), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n839), .A2(new_n703), .A3(new_n840), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT118), .ZN(new_n861));
  AND3_X1   g660(.A1(new_n860), .A2(new_n861), .A3(G134gat), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n861), .B1(new_n860), .B2(G134gat), .ZN(new_n863));
  OAI211_X1 g662(.A(new_n858), .B(new_n859), .C1(new_n862), .C2(new_n863), .ZN(G1343gat));
  NOR2_X1   g663(.A1(new_n658), .A2(new_n380), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n866), .A2(new_n456), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n830), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n743), .A2(new_n303), .ZN(new_n869));
  XNOR2_X1  g668(.A(new_n869), .B(KEYINPUT120), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n871), .A2(KEYINPUT58), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT121), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT57), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n826), .A2(new_n874), .A3(new_n497), .A4(new_n828), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n658), .A2(new_n451), .A3(new_n456), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n821), .A2(new_n592), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n536), .B1(new_n818), .B2(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT119), .ZN(new_n879));
  OR2_X1    g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n825), .B1(new_n878), .B2(new_n879), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n380), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  OAI211_X1 g681(.A(new_n875), .B(new_n876), .C1(new_n882), .C2(new_n874), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n873), .B1(new_n883), .B2(new_n640), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(G141gat), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n883), .A2(new_n873), .A3(new_n640), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n872), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(new_n883), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n303), .B1(new_n888), .B2(new_n743), .ZN(new_n889));
  OAI21_X1  g688(.A(KEYINPUT58), .B1(new_n889), .B2(new_n871), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n887), .A2(new_n890), .ZN(G1344gat));
  INV_X1    g690(.A(new_n868), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n892), .A2(new_n305), .A3(new_n613), .ZN(new_n893));
  AOI211_X1 g692(.A(KEYINPUT59), .B(new_n305), .C1(new_n888), .C2(new_n613), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT59), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n497), .A2(new_n874), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n815), .A2(new_n809), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n877), .B1(new_n592), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(new_n850), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n896), .B1(new_n899), .B2(new_n824), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n826), .A2(new_n497), .A3(new_n828), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n900), .B1(new_n901), .B2(KEYINPUT57), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n902), .A2(new_n613), .A3(new_n876), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n895), .B1(new_n903), .B2(G148gat), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n893), .B1(new_n894), .B2(new_n904), .ZN(G1345gat));
  OAI21_X1  g704(.A(G155gat), .B1(new_n883), .B2(new_n850), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n536), .A2(new_n309), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n906), .B1(new_n868), .B2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT122), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OAI211_X1 g709(.A(new_n906), .B(KEYINPUT122), .C1(new_n868), .C2(new_n907), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(G1346gat));
  NAND3_X1  g711(.A1(new_n892), .A2(new_n310), .A3(new_n703), .ZN(new_n913));
  OAI21_X1  g712(.A(G162gat), .B1(new_n883), .B2(new_n686), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(G1347gat));
  NOR2_X1   g714(.A1(new_n646), .A2(new_n457), .ZN(new_n916));
  NAND4_X1  g715(.A1(new_n826), .A2(new_n828), .A3(new_n836), .A4(new_n916), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n917), .B(KEYINPUT123), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n918), .A2(G169gat), .A3(new_n743), .ZN(new_n919));
  INV_X1    g718(.A(new_n829), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n385), .A2(new_n646), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n920), .A2(new_n451), .A3(new_n921), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n211), .B1(new_n922), .B2(new_n640), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n919), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(KEYINPUT124), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT124), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n919), .A2(new_n926), .A3(new_n923), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n925), .A2(new_n927), .ZN(G1348gat));
  NOR4_X1   g727(.A1(new_n829), .A2(new_n457), .A3(new_n646), .A4(new_n385), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n929), .A2(new_n212), .A3(new_n613), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT123), .ZN(new_n931));
  AND2_X1   g730(.A1(new_n917), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n917), .A2(new_n931), .ZN(new_n933));
  NOR3_X1   g732(.A1(new_n932), .A2(new_n933), .A3(new_n744), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n930), .B1(new_n934), .B2(new_n212), .ZN(G1349gat));
  NOR2_X1   g734(.A1(new_n850), .A2(new_n248), .ZN(new_n936));
  AOI21_X1  g735(.A(KEYINPUT125), .B1(new_n929), .B2(new_n936), .ZN(new_n937));
  NOR3_X1   g736(.A1(new_n932), .A2(new_n933), .A3(new_n850), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n937), .B1(new_n938), .B2(new_n240), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(KEYINPUT60), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT60), .ZN(new_n941));
  OAI211_X1 g740(.A(new_n937), .B(new_n941), .C1(new_n938), .C2(new_n240), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n940), .A2(new_n942), .ZN(G1350gat));
  OR3_X1    g742(.A1(new_n922), .A2(G190gat), .A3(new_n686), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n918), .A2(new_n703), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT61), .ZN(new_n946));
  AND3_X1   g745(.A1(new_n945), .A2(new_n946), .A3(G190gat), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n946), .B1(new_n945), .B2(G190gat), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n944), .B1(new_n947), .B2(new_n948), .ZN(G1351gat));
  NOR2_X1   g748(.A1(new_n866), .A2(new_n646), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n920), .A2(new_n451), .A3(new_n950), .ZN(new_n951));
  INV_X1    g750(.A(new_n951), .ZN(new_n952));
  AOI21_X1  g751(.A(G197gat), .B1(new_n952), .B2(new_n743), .ZN(new_n953));
  NOR3_X1   g752(.A1(new_n658), .A2(new_n457), .A3(new_n646), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n954), .B1(new_n902), .B2(KEYINPUT126), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT126), .ZN(new_n956));
  AOI211_X1 g755(.A(new_n956), .B(new_n900), .C1(new_n901), .C2(KEYINPUT57), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n640), .A2(new_n325), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n953), .B1(new_n958), .B2(new_n959), .ZN(G1352gat));
  NAND2_X1  g759(.A1(new_n958), .A2(new_n613), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n961), .A2(G204gat), .ZN(new_n962));
  NOR3_X1   g761(.A1(new_n951), .A2(G204gat), .A3(new_n744), .ZN(new_n963));
  XNOR2_X1  g762(.A(new_n963), .B(KEYINPUT62), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n962), .A2(new_n964), .ZN(G1353gat));
  OR3_X1    g764(.A1(new_n951), .A2(G211gat), .A3(new_n850), .ZN(new_n966));
  INV_X1    g765(.A(new_n902), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n954), .A2(new_n536), .ZN(new_n968));
  OAI21_X1  g767(.A(G211gat), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT63), .ZN(new_n970));
  AND2_X1   g769(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n969), .A2(new_n970), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n966), .B1(new_n971), .B2(new_n972), .ZN(G1354gat));
  INV_X1    g772(.A(KEYINPUT127), .ZN(new_n974));
  INV_X1    g773(.A(G218gat), .ZN(new_n975));
  NOR2_X1   g774(.A1(new_n592), .A2(new_n975), .ZN(new_n976));
  INV_X1    g775(.A(new_n976), .ZN(new_n977));
  NOR3_X1   g776(.A1(new_n955), .A2(new_n957), .A3(new_n977), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n975), .B1(new_n951), .B2(new_n686), .ZN(new_n979));
  INV_X1    g778(.A(new_n979), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n974), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n967), .A2(new_n956), .ZN(new_n982));
  INV_X1    g781(.A(new_n957), .ZN(new_n983));
  NAND4_X1  g782(.A1(new_n982), .A2(new_n983), .A3(new_n954), .A4(new_n976), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n984), .A2(KEYINPUT127), .A3(new_n979), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n981), .A2(new_n985), .ZN(G1355gat));
endmodule


