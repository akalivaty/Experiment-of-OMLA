//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 0 1 1 1 1 1 1 0 0 0 0 0 1 1 1 0 0 0 0 1 1 0 0 0 0 1 0 0 1 1 0 1 0 0 0 1 0 1 0 1 1 0 1 1 1 0 1 0 1 0 0 1 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:26 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n672, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT25), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT16), .ZN(new_n192));
  INV_X1    g006(.A(G125), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n192), .B1(new_n193), .B2(G140), .ZN(new_n194));
  XNOR2_X1  g008(.A(G125), .B(G140), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT74), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT74), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n197), .A2(new_n193), .A3(G140), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n194), .B1(new_n199), .B2(new_n192), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G146), .ZN(new_n201));
  INV_X1    g015(.A(G146), .ZN(new_n202));
  OAI211_X1 g016(.A(new_n202), .B(new_n194), .C1(new_n199), .C2(new_n192), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G128), .ZN(new_n205));
  OAI21_X1  g019(.A(KEYINPUT23), .B1(new_n205), .B2(G119), .ZN(new_n206));
  INV_X1    g020(.A(G119), .ZN(new_n207));
  OAI21_X1  g021(.A(KEYINPUT73), .B1(new_n207), .B2(G128), .ZN(new_n208));
  XNOR2_X1  g022(.A(new_n206), .B(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G110), .ZN(new_n211));
  XOR2_X1   g025(.A(G119), .B(G128), .Z(new_n212));
  XNOR2_X1  g026(.A(KEYINPUT24), .B(G110), .ZN(new_n213));
  OAI211_X1 g027(.A(new_n204), .B(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(new_n213), .ZN(new_n215));
  XNOR2_X1  g029(.A(new_n215), .B(KEYINPUT75), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n216), .B1(G110), .B2(new_n210), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n195), .A2(new_n202), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n217), .A2(new_n201), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n214), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G953), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n221), .A2(G221), .A3(G234), .ZN(new_n222));
  XNOR2_X1  g036(.A(new_n222), .B(KEYINPUT76), .ZN(new_n223));
  XNOR2_X1  g037(.A(KEYINPUT22), .B(G137), .ZN(new_n224));
  XNOR2_X1  g038(.A(new_n223), .B(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  XNOR2_X1  g040(.A(new_n220), .B(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n191), .B1(new_n228), .B2(G902), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n227), .A2(KEYINPUT25), .A3(new_n188), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n190), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n189), .A2(G902), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n231), .B1(new_n227), .B2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n207), .A2(G116), .ZN(new_n235));
  INV_X1    g049(.A(G116), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G119), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g052(.A(KEYINPUT2), .B(G113), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G113), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(KEYINPUT2), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT2), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G113), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  XNOR2_X1  g059(.A(G116), .B(G119), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT68), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n240), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n238), .A2(new_n239), .A3(KEYINPUT68), .ZN(new_n250));
  AND2_X1   g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT70), .ZN(new_n252));
  AND2_X1   g066(.A1(KEYINPUT64), .A2(G143), .ZN(new_n253));
  NOR2_X1   g067(.A1(KEYINPUT64), .A2(G143), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n202), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(G143), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G146), .ZN(new_n257));
  OAI21_X1  g071(.A(KEYINPUT1), .B1(new_n256), .B2(G146), .ZN(new_n258));
  AOI22_X1  g072(.A1(new_n255), .A2(new_n257), .B1(G128), .B2(new_n258), .ZN(new_n259));
  OR2_X1    g073(.A1(KEYINPUT64), .A2(G143), .ZN(new_n260));
  NAND2_X1  g074(.A1(KEYINPUT64), .A2(G143), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n260), .A2(KEYINPUT65), .A3(G146), .A4(new_n261), .ZN(new_n262));
  NOR3_X1   g076(.A1(new_n253), .A2(new_n254), .A3(new_n202), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT65), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n264), .B1(new_n256), .B2(G146), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n262), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT1), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G128), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n259), .B1(new_n266), .B2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(G134), .ZN(new_n271));
  OR3_X1    g085(.A1(new_n271), .A2(KEYINPUT67), .A3(G137), .ZN(new_n272));
  INV_X1    g086(.A(G137), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n273), .A2(G134), .ZN(new_n274));
  OAI21_X1  g088(.A(KEYINPUT67), .B1(new_n271), .B2(G137), .ZN(new_n275));
  OAI211_X1 g089(.A(new_n272), .B(G131), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n274), .ZN(new_n277));
  INV_X1    g091(.A(G131), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n273), .A2(KEYINPUT11), .A3(G134), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT11), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n280), .B1(new_n271), .B2(G137), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n277), .A2(new_n278), .A3(new_n279), .A4(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n276), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n252), .B1(new_n270), .B2(new_n283), .ZN(new_n284));
  AND2_X1   g098(.A1(new_n276), .A2(new_n282), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n260), .A2(G146), .A3(new_n261), .ZN(new_n286));
  INV_X1    g100(.A(new_n265), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n268), .B1(new_n288), .B2(new_n262), .ZN(new_n289));
  OAI211_X1 g103(.A(new_n285), .B(KEYINPUT70), .C1(new_n259), .C2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n284), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n277), .A2(new_n279), .A3(new_n281), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(G131), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n282), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n255), .A2(new_n257), .ZN(new_n295));
  NAND2_X1  g109(.A1(KEYINPUT0), .A2(G128), .ZN(new_n296));
  OR2_X1    g110(.A1(KEYINPUT0), .A2(G128), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  AOI211_X1 g112(.A(KEYINPUT66), .B(new_n296), .C1(new_n288), .C2(new_n262), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT66), .ZN(new_n300));
  INV_X1    g114(.A(new_n296), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n300), .B1(new_n266), .B2(new_n301), .ZN(new_n302));
  OAI211_X1 g116(.A(new_n294), .B(new_n298), .C1(new_n299), .C2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT69), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n253), .A2(new_n254), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n265), .B1(new_n306), .B2(G146), .ZN(new_n307));
  NOR4_X1   g121(.A1(new_n253), .A2(new_n254), .A3(new_n264), .A4(new_n202), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n301), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(KEYINPUT66), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n266), .A2(new_n300), .A3(new_n301), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n312), .A2(KEYINPUT69), .A3(new_n294), .A4(new_n298), .ZN(new_n313));
  AOI211_X1 g127(.A(new_n251), .B(new_n291), .C1(new_n305), .C2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(new_n270), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(new_n285), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT30), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n303), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n291), .B1(new_n305), .B2(new_n313), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n318), .B1(new_n319), .B2(new_n317), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n314), .B1(new_n320), .B2(new_n251), .ZN(new_n321));
  XOR2_X1   g135(.A(KEYINPUT26), .B(G101), .Z(new_n322));
  INV_X1    g136(.A(G237), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n323), .A2(new_n221), .A3(G210), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n322), .B(new_n324), .ZN(new_n325));
  XNOR2_X1  g139(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n325), .B(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n321), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n303), .A2(new_n316), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(new_n251), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT28), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n331), .B1(new_n329), .B2(new_n251), .ZN(new_n332));
  INV_X1    g146(.A(new_n251), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n319), .A2(new_n333), .ZN(new_n334));
  OAI211_X1 g148(.A(new_n330), .B(new_n332), .C1(new_n334), .C2(new_n331), .ZN(new_n335));
  INV_X1    g149(.A(new_n327), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(KEYINPUT29), .B1(new_n328), .B2(new_n337), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n319), .A2(new_n333), .ZN(new_n339));
  OAI21_X1  g153(.A(KEYINPUT28), .B1(new_n339), .B2(new_n314), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n340), .A2(KEYINPUT29), .A3(new_n336), .A4(new_n332), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(new_n188), .ZN(new_n342));
  OAI21_X1  g156(.A(G472), .B1(new_n338), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT72), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  OAI211_X1 g159(.A(KEYINPUT72), .B(G472), .C1(new_n338), .C2(new_n342), .ZN(new_n346));
  AND2_X1   g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n335), .A2(new_n327), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n320), .A2(new_n251), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n350), .A2(new_n336), .A3(new_n334), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT31), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n321), .A2(KEYINPUT31), .A3(new_n336), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n349), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NOR2_X1   g169(.A1(G472), .A2(G902), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(KEYINPUT32), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  AND3_X1   g172(.A1(new_n321), .A2(KEYINPUT31), .A3(new_n336), .ZN(new_n359));
  AOI21_X1  g173(.A(KEYINPUT31), .B1(new_n321), .B2(new_n336), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n348), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT32), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n361), .A2(new_n362), .A3(new_n356), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n358), .A2(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n234), .B1(new_n347), .B2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(G478), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n366), .A2(KEYINPUT15), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n260), .A2(new_n261), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n368), .A2(new_n205), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n256), .A2(G128), .ZN(new_n370));
  OAI21_X1  g184(.A(G134), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n306), .A2(G128), .ZN(new_n372));
  OAI211_X1 g186(.A(new_n372), .B(new_n271), .C1(G128), .C2(new_n256), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  XNOR2_X1  g188(.A(KEYINPUT88), .B(G122), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n375), .A2(new_n236), .ZN(new_n376));
  AND2_X1   g190(.A1(new_n236), .A2(G122), .ZN(new_n377));
  OR2_X1    g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT14), .ZN(new_n379));
  OAI21_X1  g193(.A(G107), .B1(new_n376), .B2(new_n379), .ZN(new_n380));
  AND2_X1   g194(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n378), .A2(new_n380), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n374), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT89), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT13), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n370), .A2(new_n385), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n384), .B1(new_n369), .B2(new_n386), .ZN(new_n387));
  OAI211_X1 g201(.A(new_n372), .B(KEYINPUT89), .C1(new_n385), .C2(new_n370), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT90), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n369), .A2(new_n389), .A3(KEYINPUT13), .ZN(new_n390));
  OAI21_X1  g204(.A(KEYINPUT90), .B1(new_n372), .B2(new_n385), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n387), .A2(new_n388), .A3(new_n390), .A4(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT91), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n392), .A2(new_n393), .A3(G134), .ZN(new_n394));
  INV_X1    g208(.A(G107), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n378), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n395), .B1(new_n376), .B2(new_n377), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n373), .A2(new_n397), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n394), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n393), .B1(new_n392), .B2(G134), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n383), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  XNOR2_X1  g216(.A(KEYINPUT9), .B(G234), .ZN(new_n403));
  NOR3_X1   g217(.A1(new_n403), .A2(new_n187), .A3(G953), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  OAI211_X1 g220(.A(new_n383), .B(new_n404), .C1(new_n400), .C2(new_n401), .ZN(new_n407));
  AOI21_X1  g221(.A(G902), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n408), .A2(KEYINPUT92), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT92), .ZN(new_n410));
  AOI211_X1 g224(.A(new_n410), .B(G902), .C1(new_n406), .C2(new_n407), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n367), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  OAI22_X1  g226(.A1(new_n408), .A2(KEYINPUT92), .B1(KEYINPUT15), .B2(new_n366), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  AND2_X1   g228(.A1(new_n221), .A2(G952), .ZN(new_n415));
  NAND2_X1  g229(.A1(G234), .A2(G237), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  XOR2_X1   g231(.A(KEYINPUT21), .B(G898), .Z(new_n418));
  NAND3_X1  g232(.A1(new_n416), .A2(G902), .A3(G953), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n417), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  XOR2_X1   g234(.A(new_n420), .B(KEYINPUT93), .Z(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(G214), .ZN(new_n423));
  NOR3_X1   g237(.A1(new_n423), .A2(G237), .A3(G953), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(G143), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n425), .B1(new_n368), .B2(new_n424), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(G131), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT17), .ZN(new_n428));
  OAI211_X1 g242(.A(new_n425), .B(new_n278), .C1(new_n368), .C2(new_n424), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n427), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n426), .A2(KEYINPUT17), .A3(G131), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n201), .A2(new_n430), .A3(new_n203), .A4(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(KEYINPUT18), .A2(G131), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n426), .B(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n218), .B1(new_n199), .B2(new_n202), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n432), .A2(new_n436), .ZN(new_n437));
  XNOR2_X1  g251(.A(G113), .B(G122), .ZN(new_n438));
  INV_X1    g252(.A(G104), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n438), .B(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n437), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n432), .A2(new_n440), .A3(new_n436), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n188), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(G475), .ZN(new_n446));
  AOI22_X1  g260(.A1(new_n200), .A2(G146), .B1(new_n427), .B2(new_n429), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT19), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n448), .B1(new_n196), .B2(new_n198), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n195), .A2(KEYINPUT19), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n202), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  AOI22_X1  g265(.A1(new_n447), .A2(new_n451), .B1(new_n434), .B2(new_n435), .ZN(new_n452));
  OAI21_X1  g266(.A(KEYINPUT87), .B1(new_n452), .B2(new_n440), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n427), .A2(new_n429), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n201), .A2(new_n454), .A3(new_n451), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(new_n436), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT87), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n456), .A2(new_n457), .A3(new_n441), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n453), .A2(new_n443), .A3(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT20), .ZN(new_n460));
  NOR2_X1   g274(.A1(G475), .A2(G902), .ZN(new_n461));
  AND3_X1   g275(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n460), .B1(new_n459), .B2(new_n461), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n446), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NOR3_X1   g278(.A1(new_n414), .A2(new_n422), .A3(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(G214), .B1(G237), .B2(G902), .ZN(new_n466));
  XOR2_X1   g280(.A(new_n466), .B(KEYINPUT81), .Z(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(KEYINPUT78), .B1(new_n395), .B2(G104), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT78), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n470), .A2(new_n439), .A3(G107), .ZN(new_n471));
  AND3_X1   g285(.A1(new_n395), .A2(KEYINPUT3), .A3(G104), .ZN(new_n472));
  AOI21_X1  g286(.A(KEYINPUT3), .B1(new_n395), .B2(G104), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n469), .B(new_n471), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(G101), .ZN(new_n475));
  AND2_X1   g289(.A1(new_n469), .A2(new_n471), .ZN(new_n476));
  INV_X1    g290(.A(G101), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT3), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n478), .B1(new_n439), .B2(G107), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n395), .A2(KEYINPUT3), .A3(G104), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n476), .A2(new_n477), .A3(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n475), .A2(KEYINPUT4), .A3(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n477), .B1(new_n476), .B2(new_n481), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT4), .ZN(new_n485));
  AOI21_X1  g299(.A(KEYINPUT79), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  AND4_X1   g300(.A1(KEYINPUT79), .A2(new_n474), .A3(new_n485), .A4(G101), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n251), .B(new_n483), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT82), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  XNOR2_X1  g304(.A(G110), .B(G122), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n474), .A2(new_n485), .A3(G101), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT79), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n484), .A2(KEYINPUT79), .A3(new_n485), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n496), .A2(KEYINPUT82), .A3(new_n251), .A4(new_n483), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n439), .A2(G107), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n395), .A2(G104), .ZN(new_n499));
  OAI21_X1  g313(.A(G101), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n482), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(G113), .B1(new_n235), .B2(KEYINPUT5), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n503), .B1(KEYINPUT5), .B2(new_n246), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n504), .B1(new_n246), .B2(new_n245), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n490), .A2(new_n491), .A3(new_n497), .A4(new_n506), .ZN(new_n507));
  XOR2_X1   g321(.A(KEYINPUT84), .B(KEYINPUT8), .Z(new_n508));
  XNOR2_X1  g322(.A(new_n508), .B(new_n491), .ZN(new_n509));
  INV_X1    g323(.A(new_n506), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n502), .A2(new_n505), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NOR3_X1   g326(.A1(new_n289), .A2(G125), .A3(new_n259), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n221), .A2(G224), .ZN(new_n514));
  XOR2_X1   g328(.A(new_n514), .B(KEYINPUT83), .Z(new_n515));
  INV_X1    g329(.A(KEYINPUT7), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n298), .B1(new_n299), .B2(new_n302), .ZN(new_n518));
  AOI211_X1 g332(.A(new_n513), .B(new_n517), .C1(new_n518), .C2(G125), .ZN(new_n519));
  INV_X1    g333(.A(new_n517), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n518), .A2(G125), .ZN(new_n521));
  INV_X1    g335(.A(new_n513), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n507), .B(new_n512), .C1(new_n519), .C2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(new_n188), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT85), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n491), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n497), .A2(new_n506), .ZN(new_n529));
  AND2_X1   g343(.A1(new_n488), .A2(new_n489), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n531), .A2(KEYINPUT6), .A3(new_n507), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT6), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n533), .B(new_n528), .C1(new_n529), .C2(new_n530), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n521), .A2(new_n522), .ZN(new_n535));
  XNOR2_X1  g349(.A(new_n535), .B(new_n515), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n532), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n524), .A2(KEYINPUT85), .A3(new_n188), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n527), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(G210), .B1(G237), .B2(G902), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n539), .A2(KEYINPUT86), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n539), .A2(new_n541), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT86), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n527), .A2(new_n540), .A3(new_n537), .A4(new_n538), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n465), .A2(new_n468), .A3(new_n542), .A4(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(G469), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n312), .A2(new_n496), .A3(new_n298), .A4(new_n483), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n267), .B1(new_n368), .B2(new_n202), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n288), .B(new_n262), .C1(new_n550), .C2(new_n205), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n266), .A2(new_n269), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(new_n502), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT10), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n294), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n501), .A2(new_n555), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(new_n315), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n549), .A2(new_n556), .A3(new_n557), .A4(new_n559), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n315), .A2(new_n502), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n501), .B1(new_n552), .B2(new_n551), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n294), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(KEYINPUT12), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n221), .A2(G227), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n565), .B(KEYINPUT77), .ZN(new_n566));
  XNOR2_X1  g380(.A(G110), .B(G140), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n566), .B(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT12), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n570), .B(new_n294), .C1(new_n561), .C2(new_n562), .ZN(new_n571));
  AND4_X1   g385(.A1(new_n560), .A2(new_n564), .A3(new_n569), .A4(new_n571), .ZN(new_n572));
  AND4_X1   g386(.A1(new_n312), .A2(new_n496), .A3(new_n298), .A4(new_n483), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n559), .B1(KEYINPUT10), .B2(new_n562), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n294), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n569), .B1(new_n575), .B2(new_n560), .ZN(new_n576));
  OAI211_X1 g390(.A(new_n548), .B(new_n188), .C1(new_n572), .C2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(G469), .A2(G902), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n564), .A2(new_n560), .A3(new_n571), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(new_n568), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n575), .A2(new_n560), .A3(new_n569), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n580), .A2(G469), .A3(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n577), .A2(new_n578), .A3(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(G221), .B1(new_n403), .B2(G902), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT80), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n585), .B(new_n586), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n547), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n365), .A2(new_n588), .ZN(new_n589));
  XNOR2_X1  g403(.A(KEYINPUT94), .B(G101), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n589), .B(new_n590), .ZN(G3));
  OAI21_X1  g405(.A(G472), .B1(new_n355), .B2(G902), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n361), .A2(new_n356), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n587), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n543), .A2(KEYINPUT95), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT95), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n539), .A2(new_n597), .A3(new_n541), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n596), .A2(new_n545), .A3(new_n598), .ZN(new_n599));
  AND2_X1   g413(.A1(new_n599), .A2(new_n466), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT97), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT96), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n602), .B1(new_n408), .B2(G478), .ZN(new_n603));
  INV_X1    g417(.A(new_n407), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n392), .A2(G134), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(KEYINPUT91), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n606), .A2(new_n394), .A3(new_n399), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n404), .B1(new_n607), .B2(new_n383), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n188), .B1(new_n604), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n609), .A2(KEYINPUT96), .A3(new_n366), .ZN(new_n610));
  OAI21_X1  g424(.A(KEYINPUT33), .B1(new_n604), .B2(new_n608), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT33), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n406), .A2(new_n612), .A3(new_n407), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n366), .A2(G902), .ZN(new_n615));
  AOI22_X1  g429(.A1(new_n603), .A2(new_n610), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n464), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n601), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n613), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n612), .B1(new_n406), .B2(new_n407), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n615), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(KEYINPUT96), .B1(new_n609), .B2(new_n366), .ZN(new_n622));
  NOR3_X1   g436(.A1(new_n408), .A2(new_n602), .A3(G478), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n624), .A2(KEYINPUT97), .A3(new_n464), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n422), .B1(new_n618), .B2(new_n625), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n595), .A2(new_n233), .A3(new_n600), .A4(new_n626), .ZN(new_n627));
  XOR2_X1   g441(.A(KEYINPUT34), .B(G104), .Z(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(G6));
  AOI211_X1 g443(.A(new_n422), .B(new_n464), .C1(new_n412), .C2(new_n413), .ZN(new_n630));
  AND2_X1   g444(.A1(new_n233), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n595), .A2(new_n600), .A3(new_n631), .ZN(new_n632));
  XOR2_X1   g446(.A(KEYINPUT35), .B(G107), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G9));
  NOR2_X1   g448(.A1(new_n225), .A2(KEYINPUT36), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n220), .B(new_n635), .ZN(new_n636));
  AND2_X1   g450(.A1(new_n636), .A2(new_n232), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n231), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n547), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n595), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT37), .B(G110), .Z(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G12));
  OR2_X1    g456(.A1(new_n419), .A2(G900), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n417), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n414), .A2(new_n617), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(KEYINPUT98), .ZN(new_n646));
  INV_X1    g460(.A(new_n638), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT98), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n414), .A2(new_n648), .A3(new_n617), .A4(new_n644), .ZN(new_n649));
  AND3_X1   g463(.A1(new_n646), .A2(new_n647), .A3(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n364), .A2(new_n346), .A3(new_n345), .ZN(new_n651));
  INV_X1    g465(.A(new_n587), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n650), .A2(new_n651), .A3(new_n652), .A4(new_n600), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G128), .ZN(G30));
  XOR2_X1   g468(.A(new_n644), .B(KEYINPUT39), .Z(new_n655));
  OR2_X1    g469(.A1(new_n587), .A2(new_n655), .ZN(new_n656));
  OR2_X1    g470(.A1(new_n656), .A2(KEYINPUT40), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n617), .B1(new_n412), .B2(new_n413), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n638), .A2(new_n466), .A3(new_n658), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n659), .B1(new_n656), .B2(KEYINPUT40), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n546), .A2(new_n542), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  OR2_X1    g478(.A1(new_n339), .A2(new_n314), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n188), .B1(new_n665), .B2(new_n336), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n321), .A2(new_n327), .ZN(new_n667));
  OAI21_X1  g481(.A(G472), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n364), .A2(new_n668), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n657), .A2(new_n660), .A3(new_n664), .A4(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(new_n368), .ZN(G45));
  NOR2_X1   g485(.A1(new_n616), .A2(new_n617), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(new_n644), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n673), .A2(new_n638), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n651), .A2(new_n600), .A3(new_n652), .A4(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G146), .ZN(G48));
  INV_X1    g490(.A(new_n584), .ZN(new_n677));
  OR2_X1    g491(.A1(new_n572), .A2(new_n576), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(new_n188), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(G469), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n680), .A2(KEYINPUT100), .A3(new_n577), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT100), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n679), .A2(new_n682), .A3(G469), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n677), .B1(new_n681), .B2(new_n683), .ZN(new_n684));
  AND4_X1   g498(.A1(new_n466), .A2(new_n626), .A3(new_n684), .A4(new_n599), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(new_n365), .ZN(new_n686));
  XNOR2_X1  g500(.A(KEYINPUT41), .B(G113), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G15));
  AND3_X1   g502(.A1(new_n684), .A2(new_n466), .A3(new_n599), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n689), .A2(new_n651), .A3(new_n631), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G116), .ZN(G18));
  AND2_X1   g505(.A1(new_n647), .A2(new_n465), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n689), .A2(new_n651), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G119), .ZN(G21));
  INV_X1    g508(.A(new_n684), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n695), .A2(new_n422), .ZN(new_n696));
  AND2_X1   g510(.A1(new_n340), .A2(new_n332), .ZN(new_n697));
  OAI22_X1  g511(.A1(new_n359), .A2(new_n360), .B1(new_n697), .B2(new_n336), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(new_n356), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n592), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n234), .A2(new_n700), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n696), .A2(new_n701), .A3(new_n600), .A4(new_n658), .ZN(new_n702));
  XOR2_X1   g516(.A(KEYINPUT101), .B(G122), .Z(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(G24));
  NOR3_X1   g518(.A1(new_n700), .A2(new_n638), .A3(new_n673), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n689), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G125), .ZN(G27));
  NOR3_X1   g521(.A1(new_n355), .A2(KEYINPUT32), .A3(new_n357), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n362), .B1(new_n361), .B2(new_n356), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n345), .A2(new_n346), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n233), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(new_n466), .ZN(new_n713));
  AOI211_X1 g527(.A(KEYINPUT104), .B(new_n713), .C1(new_n546), .C2(new_n542), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT104), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n715), .B1(new_n661), .B2(new_n466), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n712), .A2(new_n714), .A3(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(new_n673), .ZN(new_n718));
  OR2_X1    g532(.A1(new_n581), .A2(KEYINPUT102), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n581), .A2(KEYINPUT102), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n719), .A2(new_n580), .A3(new_n720), .ZN(new_n721));
  OAI211_X1 g535(.A(new_n577), .B(new_n578), .C1(new_n721), .C2(new_n548), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(new_n584), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(KEYINPUT103), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT103), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n722), .A2(new_n725), .A3(new_n584), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n717), .A2(KEYINPUT42), .A3(new_n718), .A4(new_n727), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n716), .A2(new_n714), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n365), .A2(new_n729), .A3(new_n718), .A4(new_n727), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT42), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n728), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G131), .ZN(G33));
  AND2_X1   g548(.A1(new_n646), .A2(new_n649), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n365), .A2(new_n729), .A3(new_n735), .A4(new_n727), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G134), .ZN(G36));
  NAND2_X1  g551(.A1(new_n661), .A2(new_n466), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(KEYINPUT104), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n661), .A2(new_n715), .A3(new_n466), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n616), .A2(new_n464), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(KEYINPUT43), .ZN(new_n743));
  INV_X1    g557(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n744), .A2(KEYINPUT105), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT105), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n743), .A2(new_n746), .ZN(new_n747));
  OAI211_X1 g561(.A(new_n594), .B(new_n647), .C1(new_n745), .C2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT44), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n741), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n750), .B1(new_n749), .B2(new_n748), .ZN(new_n751));
  OR2_X1    g565(.A1(new_n751), .A2(KEYINPUT106), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(KEYINPUT106), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT45), .ZN(new_n754));
  OR2_X1    g568(.A1(new_n721), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n580), .A2(new_n581), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n548), .B1(new_n756), .B2(new_n754), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n578), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT46), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(new_n577), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n759), .A2(new_n760), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n584), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n764), .A2(new_n655), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n752), .A2(new_n753), .A3(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G137), .ZN(G39));
  XNOR2_X1  g581(.A(new_n764), .B(KEYINPUT47), .ZN(new_n768));
  NOR4_X1   g582(.A1(new_n741), .A2(new_n233), .A3(new_n651), .A4(new_n673), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n768), .B1(KEYINPUT107), .B2(new_n769), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n770), .B1(KEYINPUT107), .B2(new_n769), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G140), .ZN(G42));
  INV_X1    g586(.A(KEYINPUT54), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT110), .ZN(new_n774));
  AND4_X1   g588(.A1(new_n365), .A2(new_n729), .A3(new_n735), .A4(new_n727), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n705), .A2(new_n727), .ZN(new_n776));
  INV_X1    g590(.A(new_n644), .ZN(new_n777));
  NOR4_X1   g591(.A1(new_n638), .A2(new_n464), .A3(new_n414), .A4(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n651), .A2(new_n652), .A3(new_n778), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n741), .B1(new_n776), .B2(new_n779), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n774), .B1(new_n775), .B2(new_n780), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n587), .B1(new_n347), .B2(new_n364), .ZN(new_n782));
  AOI22_X1  g596(.A1(new_n782), .A2(new_n778), .B1(new_n705), .B2(new_n727), .ZN(new_n783));
  OAI211_X1 g597(.A(KEYINPUT110), .B(new_n736), .C1(new_n783), .C2(new_n741), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n733), .A2(new_n781), .A3(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT109), .ZN(new_n786));
  INV_X1    g600(.A(new_n661), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT108), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n787), .A2(new_n788), .A3(new_n468), .A4(new_n630), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n630), .A2(new_n468), .A3(new_n546), .A4(new_n542), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n790), .A2(KEYINPUT108), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n789), .A2(new_n595), .A3(new_n791), .A4(new_n233), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n786), .B1(new_n792), .B2(new_n640), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  OAI211_X1 g608(.A(new_n689), .B(new_n651), .C1(new_n631), .C2(new_n692), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n672), .A2(new_n421), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n661), .A2(new_n796), .A3(new_n467), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n595), .A2(new_n797), .A3(new_n233), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n795), .A2(new_n702), .A3(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n792), .A2(new_n786), .A3(new_n640), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n365), .B1(new_n685), .B2(new_n588), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n794), .A2(new_n799), .A3(new_n800), .A4(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n785), .A2(new_n802), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n647), .A2(new_n723), .A3(new_n777), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n804), .A2(new_n600), .A3(new_n669), .A4(new_n658), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n653), .A2(new_n706), .A3(new_n805), .A4(new_n675), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT112), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT52), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n806), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n806), .B(KEYINPUT52), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(KEYINPUT112), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n803), .A2(KEYINPUT53), .A3(new_n809), .A4(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT111), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n813), .B1(new_n785), .B2(new_n802), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n736), .B1(new_n783), .B2(new_n741), .ZN(new_n815));
  AOI22_X1  g629(.A1(new_n815), .A2(new_n774), .B1(new_n728), .B2(new_n732), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n801), .A2(new_n702), .A3(new_n795), .A4(new_n798), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n792), .A2(new_n786), .A3(new_n640), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n817), .A2(new_n818), .A3(new_n793), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n816), .A2(new_n819), .A3(KEYINPUT111), .A4(new_n784), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n810), .B1(new_n814), .B2(new_n820), .ZN(new_n821));
  OAI211_X1 g635(.A(new_n773), .B(new_n812), .C1(new_n821), .C2(KEYINPUT53), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT113), .ZN(new_n823));
  OR2_X1    g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n822), .A2(new_n823), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n814), .A2(new_n820), .ZN(new_n826));
  INV_X1    g640(.A(new_n810), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(KEYINPUT53), .ZN(new_n829));
  INV_X1    g643(.A(new_n826), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT53), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n811), .A2(new_n831), .A3(new_n809), .ZN(new_n832));
  OAI211_X1 g646(.A(new_n829), .B(KEYINPUT54), .C1(new_n830), .C2(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n824), .A2(new_n825), .A3(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT114), .ZN(new_n835));
  XNOR2_X1  g649(.A(new_n834), .B(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n741), .A2(new_n695), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n669), .A2(new_n234), .A3(new_n417), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  XOR2_X1   g653(.A(new_n839), .B(KEYINPUT115), .Z(new_n840));
  NAND3_X1  g654(.A1(new_n840), .A2(new_n617), .A3(new_n616), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n681), .A2(new_n683), .ZN(new_n842));
  INV_X1    g656(.A(new_n842), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n768), .B1(new_n584), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n744), .A2(new_n417), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(new_n701), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n846), .A2(new_n741), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n700), .A2(new_n638), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n837), .A2(new_n845), .ZN(new_n849));
  AOI22_X1  g663(.A1(new_n844), .A2(new_n847), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NOR4_X1   g664(.A1(new_n846), .A2(new_n466), .A3(new_n664), .A4(new_n695), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n851), .B(KEYINPUT50), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n841), .A2(new_n850), .A3(new_n852), .ZN(new_n853));
  OR2_X1    g667(.A1(new_n853), .A2(KEYINPUT51), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(KEYINPUT51), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n849), .A2(new_n365), .ZN(new_n856));
  XNOR2_X1  g670(.A(new_n856), .B(KEYINPUT48), .ZN(new_n857));
  XOR2_X1   g671(.A(new_n415), .B(KEYINPUT116), .Z(new_n858));
  INV_X1    g672(.A(new_n689), .ZN(new_n859));
  OAI211_X1 g673(.A(new_n857), .B(new_n858), .C1(new_n859), .C2(new_n846), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n618), .A2(new_n625), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n860), .B1(new_n861), .B2(new_n840), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n854), .A2(new_n855), .A3(new_n862), .ZN(new_n863));
  OAI22_X1  g677(.A1(new_n836), .A2(new_n863), .B1(G952), .B2(G953), .ZN(new_n864));
  XOR2_X1   g678(.A(new_n842), .B(KEYINPUT49), .Z(new_n865));
  NAND4_X1  g679(.A1(new_n233), .A2(new_n584), .A3(new_n468), .A4(new_n742), .ZN(new_n866));
  OR4_X1    g680(.A1(new_n664), .A2(new_n865), .A3(new_n669), .A4(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n864), .A2(new_n867), .ZN(G75));
  NOR2_X1   g682(.A1(new_n221), .A2(G952), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n532), .A2(new_n534), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n870), .B(new_n536), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n871), .B(KEYINPUT55), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n812), .B1(new_n821), .B2(KEYINPUT53), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n873), .A2(G210), .A3(G902), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT56), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n872), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n873), .A2(G902), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(KEYINPUT117), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT117), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n873), .A2(new_n879), .A3(G902), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n878), .A2(new_n541), .A3(new_n880), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n872), .A2(new_n875), .ZN(new_n882));
  AOI211_X1 g696(.A(new_n869), .B(new_n876), .C1(new_n881), .C2(new_n882), .ZN(G51));
  INV_X1    g697(.A(new_n758), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n878), .A2(new_n884), .A3(new_n880), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(KEYINPUT119), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT119), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n878), .A2(new_n887), .A3(new_n884), .A4(new_n880), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n873), .A2(KEYINPUT54), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(new_n822), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n578), .B(KEYINPUT118), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n891), .B(KEYINPUT57), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(new_n678), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n886), .A2(new_n888), .A3(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(new_n869), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT120), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n895), .A2(KEYINPUT120), .A3(new_n896), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(G54));
  INV_X1    g715(.A(new_n459), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n878), .A2(new_n880), .ZN(new_n903));
  NAND2_X1  g717(.A1(KEYINPUT58), .A2(G475), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n902), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(new_n896), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n903), .A2(new_n902), .A3(new_n904), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n906), .A2(new_n907), .ZN(G60));
  NAND2_X1  g722(.A1(G478), .A2(G902), .ZN(new_n909));
  XOR2_X1   g723(.A(new_n909), .B(KEYINPUT59), .Z(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n890), .A2(new_n614), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(new_n896), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n836), .A2(new_n911), .ZN(new_n914));
  INV_X1    g728(.A(new_n614), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n913), .B1(new_n914), .B2(new_n915), .ZN(G63));
  XNOR2_X1  g730(.A(KEYINPUT121), .B(KEYINPUT61), .ZN(new_n917));
  NAND2_X1  g731(.A1(G217), .A2(G902), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n918), .B(KEYINPUT122), .Z(new_n919));
  XOR2_X1   g733(.A(new_n919), .B(KEYINPUT60), .Z(new_n920));
  AND2_X1   g734(.A1(new_n873), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n921), .A2(new_n636), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(new_n896), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n921), .A2(new_n227), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n917), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n924), .B(KEYINPUT123), .Z(new_n926));
  NAND3_X1  g740(.A1(new_n922), .A2(KEYINPUT61), .A3(new_n896), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n925), .B1(new_n926), .B2(new_n927), .ZN(G66));
  AOI21_X1  g742(.A(new_n221), .B1(new_n418), .B2(G224), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n929), .B1(new_n802), .B2(new_n221), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n870), .B1(G898), .B2(new_n221), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n930), .B(new_n931), .Z(G69));
  AND2_X1   g746(.A1(new_n766), .A2(new_n771), .ZN(new_n933));
  AND2_X1   g747(.A1(new_n653), .A2(new_n706), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n670), .A2(new_n675), .A3(new_n934), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n935), .B(KEYINPUT62), .Z(new_n936));
  AOI21_X1  g750(.A(new_n672), .B1(new_n617), .B2(new_n414), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n656), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n717), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n933), .A2(new_n936), .A3(new_n939), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n320), .B(KEYINPUT124), .Z(new_n941));
  NOR2_X1   g755(.A1(new_n449), .A2(new_n450), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n941), .B(new_n942), .Z(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n940), .A2(new_n221), .A3(new_n944), .ZN(new_n945));
  OAI21_X1  g759(.A(G900), .B1(new_n943), .B2(G227), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(G953), .ZN(new_n947));
  NAND4_X1  g761(.A1(new_n765), .A2(new_n365), .A3(new_n600), .A4(new_n658), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n948), .A2(new_n736), .ZN(new_n949));
  AND4_X1   g763(.A1(new_n675), .A2(new_n949), .A3(new_n733), .A4(new_n934), .ZN(new_n950));
  AOI21_X1  g764(.A(G953), .B1(new_n933), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n943), .B1(G227), .B2(new_n221), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n945), .B(new_n947), .C1(new_n951), .C2(new_n952), .ZN(G72));
  NAND3_X1  g767(.A1(new_n933), .A2(new_n819), .A3(new_n950), .ZN(new_n954));
  XNOR2_X1  g768(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n955));
  NAND2_X1  g769(.A1(G472), .A2(G902), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n955), .B(new_n956), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n957), .B(KEYINPUT126), .Z(new_n958));
  NAND2_X1  g772(.A1(new_n954), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n328), .B1(new_n959), .B2(KEYINPUT127), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n960), .B1(KEYINPUT127), .B2(new_n959), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n958), .B1(new_n940), .B2(new_n802), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n869), .B1(new_n962), .B2(new_n667), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n829), .B1(new_n830), .B2(new_n832), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n328), .A2(new_n957), .ZN(new_n966));
  NOR3_X1   g780(.A1(new_n965), .A2(new_n667), .A3(new_n966), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n964), .A2(new_n967), .ZN(G57));
endmodule


