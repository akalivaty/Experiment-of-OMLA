//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 1 1 1 1 0 0 1 1 0 0 0 0 0 0 0 0 1 1 0 0 0 0 1 1 1 0 0 1 0 0 1 0 0 0 0 0 0 1 1 0 1 1 1 1 1 0 1 0 0 1 1 1 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:21 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n445, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n546, new_n547, new_n548, new_n549, new_n550, new_n552,
    new_n554, new_n555, new_n556, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n565, new_n566, new_n567, new_n569, new_n570,
    new_n571, new_n573, new_n574, new_n575, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n587, new_n588,
    new_n591, new_n592, new_n594, new_n595, new_n596, new_n597, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1104, new_n1105, new_n1106,
    new_n1107;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT65), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT66), .Z(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G125), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n461), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n462), .A2(G2105), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n468), .A2(G2105), .B1(G101), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT67), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n472), .A2(new_n462), .A3(KEYINPUT3), .ZN(new_n473));
  AOI21_X1  g048(.A(KEYINPUT67), .B1(new_n464), .B2(G2104), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n464), .A2(G2104), .ZN(new_n475));
  OAI211_X1 g050(.A(new_n471), .B(new_n473), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G137), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n470), .A2(new_n478), .ZN(new_n479));
  XOR2_X1   g054(.A(new_n479), .B(KEYINPUT68), .Z(G160));
  OAI211_X1 g055(.A(G2105), .B(new_n473), .C1(new_n474), .C2(new_n475), .ZN(new_n481));
  INV_X1    g056(.A(G124), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT69), .ZN(new_n484));
  XNOR2_X1  g059(.A(new_n483), .B(new_n484), .ZN(new_n485));
  OAI21_X1  g060(.A(KEYINPUT70), .B1(G100), .B2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  NOR3_X1   g062(.A1(KEYINPUT70), .A2(G100), .A3(G2105), .ZN(new_n488));
  OAI221_X1 g063(.A(G2104), .B1(G112), .B2(new_n471), .C1(new_n487), .C2(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n477), .A2(G136), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n485), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G162));
  OAI21_X1  g067(.A(new_n472), .B1(new_n462), .B2(KEYINPUT3), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(new_n463), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n494), .A2(G138), .A3(new_n471), .A4(new_n473), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n497), .A2(new_n471), .A3(G138), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n466), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(G126), .ZN(new_n502));
  NOR2_X1   g077(.A1(G102), .A2(G2105), .ZN(new_n503));
  OAI21_X1  g078(.A(G2104), .B1(new_n471), .B2(G114), .ZN(new_n504));
  OAI22_X1  g079(.A1(new_n481), .A2(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n501), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(G164));
  INV_X1    g083(.A(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(KEYINPUT5), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT5), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G543), .ZN(new_n512));
  AND2_X1   g087(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n513), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  XOR2_X1   g091(.A(new_n516), .B(KEYINPUT71), .Z(new_n517));
  XNOR2_X1  g092(.A(KEYINPUT6), .B(G651), .ZN(new_n518));
  AND2_X1   g093(.A1(new_n518), .A2(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G50), .ZN(new_n520));
  INV_X1    g095(.A(G88), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n513), .A2(new_n518), .ZN(new_n522));
  OAI211_X1 g097(.A(new_n517), .B(new_n520), .C1(new_n521), .C2(new_n522), .ZN(G303));
  INV_X1    g098(.A(G303), .ZN(G166));
  OR2_X1    g099(.A1(new_n519), .A2(KEYINPUT73), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n519), .A2(KEYINPUT73), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G51), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT7), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n513), .A2(G63), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT72), .ZN(new_n533));
  INV_X1    g108(.A(new_n522), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G89), .ZN(new_n535));
  NAND4_X1  g110(.A1(new_n529), .A2(new_n531), .A3(new_n533), .A4(new_n535), .ZN(G286));
  INV_X1    g111(.A(G286), .ZN(G168));
  NAND2_X1  g112(.A1(new_n513), .A2(G64), .ZN(new_n538));
  INV_X1    g113(.A(G77), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n539), .B2(new_n509), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G651), .ZN(new_n541));
  INV_X1    g116(.A(G90), .ZN(new_n542));
  INV_X1    g117(.A(G52), .ZN(new_n543));
  OAI221_X1 g118(.A(new_n541), .B1(new_n542), .B2(new_n522), .C1(new_n527), .C2(new_n543), .ZN(G301));
  INV_X1    g119(.A(G301), .ZN(G171));
  AND2_X1   g120(.A1(new_n528), .A2(G43), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n513), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n547));
  INV_X1    g122(.A(G81), .ZN(new_n548));
  OAI22_X1  g123(.A1(new_n547), .A2(new_n515), .B1(new_n522), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  AND3_X1   g126(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G36), .ZN(G176));
  XOR2_X1   g128(.A(KEYINPUT74), .B(KEYINPUT8), .Z(new_n554));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n554), .B(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n552), .A2(new_n556), .ZN(G188));
  AND3_X1   g132(.A1(new_n518), .A2(G53), .A3(G543), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT9), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n558), .B(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n534), .A2(G91), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n513), .B(KEYINPUT75), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n562), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n563));
  OAI211_X1 g138(.A(new_n560), .B(new_n561), .C1(new_n563), .C2(new_n515), .ZN(G299));
  NAND2_X1  g139(.A1(new_n534), .A2(G87), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n519), .A2(G49), .ZN(new_n566));
  OAI21_X1  g141(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(G288));
  NAND2_X1  g143(.A1(new_n519), .A2(G48), .ZN(new_n569));
  INV_X1    g144(.A(G86), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n513), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n571));
  OAI221_X1 g146(.A(new_n569), .B1(new_n570), .B2(new_n522), .C1(new_n571), .C2(new_n515), .ZN(G305));
  NAND2_X1  g147(.A1(new_n534), .A2(G85), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n574));
  INV_X1    g149(.A(G47), .ZN(new_n575));
  OAI221_X1 g150(.A(new_n573), .B1(new_n515), .B2(new_n574), .C1(new_n527), .C2(new_n575), .ZN(G290));
  NAND2_X1  g151(.A1(G301), .A2(G868), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n562), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n578), .A2(new_n515), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n579), .B1(G54), .B2(new_n528), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n534), .A2(G92), .ZN(new_n581));
  XOR2_X1   g156(.A(new_n581), .B(KEYINPUT10), .Z(new_n582));
  NAND2_X1  g157(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n577), .B1(new_n584), .B2(G868), .ZN(G284));
  OAI21_X1  g160(.A(new_n577), .B1(new_n584), .B2(G868), .ZN(G321));
  NAND2_X1  g161(.A1(G286), .A2(G868), .ZN(new_n587));
  INV_X1    g162(.A(G299), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(G868), .B2(new_n588), .ZN(G297));
  OAI21_X1  g164(.A(new_n587), .B1(G868), .B2(new_n588), .ZN(G280));
  INV_X1    g165(.A(G559), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n584), .B1(new_n591), .B2(G860), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n592), .B(KEYINPUT76), .ZN(G148));
  NAND2_X1  g168(.A1(new_n584), .A2(new_n591), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(G868), .ZN(new_n595));
  OR2_X1    g170(.A1(new_n595), .A2(KEYINPUT77), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(KEYINPUT77), .ZN(new_n597));
  OAI211_X1 g172(.A(new_n596), .B(new_n597), .C1(G868), .C2(new_n550), .ZN(G323));
  XNOR2_X1  g173(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g174(.A(new_n481), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n600), .A2(G123), .ZN(new_n601));
  XOR2_X1   g176(.A(new_n601), .B(KEYINPUT81), .Z(new_n602));
  NAND2_X1  g177(.A1(new_n477), .A2(G135), .ZN(new_n603));
  NOR2_X1   g178(.A1(G99), .A2(G2105), .ZN(new_n604));
  OAI21_X1  g179(.A(G2104), .B1(new_n471), .B2(G111), .ZN(new_n605));
  OAI211_X1 g180(.A(new_n602), .B(new_n603), .C1(new_n604), .C2(new_n605), .ZN(new_n606));
  XOR2_X1   g181(.A(new_n606), .B(KEYINPUT82), .Z(new_n607));
  OR2_X1    g182(.A1(new_n607), .A2(G2096), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(G2096), .ZN(new_n609));
  XNOR2_X1  g184(.A(KEYINPUT78), .B(KEYINPUT12), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n471), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n610), .B(new_n611), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT13), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n613), .A2(G2100), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT80), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n613), .A2(G2100), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(KEYINPUT79), .Z(new_n617));
  NAND4_X1  g192(.A1(new_n608), .A2(new_n609), .A3(new_n615), .A4(new_n617), .ZN(G156));
  XNOR2_X1  g193(.A(G2451), .B(G2454), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT16), .ZN(new_n620));
  XNOR2_X1  g195(.A(G2443), .B(G2446), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XNOR2_X1  g197(.A(G1341), .B(G1348), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n622), .B(new_n623), .Z(new_n624));
  XOR2_X1   g199(.A(G2427), .B(G2430), .Z(new_n625));
  XNOR2_X1  g200(.A(KEYINPUT15), .B(G2435), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(KEYINPUT84), .B(G2438), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(KEYINPUT83), .B(KEYINPUT14), .Z(new_n630));
  NAND2_X1  g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n624), .B(new_n631), .ZN(new_n632));
  AND2_X1   g207(.A1(new_n632), .A2(G14), .ZN(G401));
  XOR2_X1   g208(.A(G2072), .B(G2078), .Z(new_n634));
  XOR2_X1   g209(.A(G2084), .B(G2090), .Z(new_n635));
  INV_X1    g210(.A(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(G2067), .B(G2678), .Z(new_n637));
  OR2_X1    g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT85), .B(KEYINPUT18), .ZN(new_n639));
  AOI21_X1  g214(.A(new_n634), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(G2096), .Z(new_n641));
  INV_X1    g216(.A(KEYINPUT17), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n642), .B1(new_n636), .B2(new_n637), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n639), .B1(new_n638), .B2(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n641), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT86), .B(G2100), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(G227));
  XNOR2_X1  g222(.A(G1971), .B(G1976), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT87), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(KEYINPUT19), .Z(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(G1956), .B(G2474), .Z(new_n652));
  XOR2_X1   g227(.A(G1961), .B(G1966), .Z(new_n653));
  NAND2_X1  g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n652), .A2(new_n653), .ZN(new_n656));
  OR3_X1    g231(.A1(new_n651), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n650), .A2(new_n654), .ZN(new_n658));
  XOR2_X1   g233(.A(KEYINPUT88), .B(KEYINPUT20), .Z(new_n659));
  AOI22_X1  g234(.A1(new_n658), .A2(new_n659), .B1(new_n651), .B2(new_n656), .ZN(new_n660));
  OAI211_X1 g235(.A(new_n657), .B(new_n660), .C1(new_n658), .C2(new_n659), .ZN(new_n661));
  XOR2_X1   g236(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT89), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n661), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1991), .B(G1996), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1981), .B(G1986), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(G229));
  INV_X1    g243(.A(G16), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n669), .A2(G19), .ZN(new_n670));
  OAI21_X1  g245(.A(new_n670), .B1(new_n550), .B2(new_n669), .ZN(new_n671));
  MUX2_X1   g246(.A(new_n670), .B(new_n671), .S(KEYINPUT92), .Z(new_n672));
  OR2_X1    g247(.A1(new_n672), .A2(G1341), .ZN(new_n673));
  OR2_X1    g248(.A1(G29), .A2(G32), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n477), .A2(G141), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n675), .B(KEYINPUT94), .Z(new_n676));
  NAND3_X1  g251(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(KEYINPUT26), .Z(new_n678));
  AOI22_X1  g253(.A1(new_n600), .A2(G129), .B1(G105), .B2(new_n469), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n676), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(G29), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n674), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT27), .B(G1996), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n682), .A2(new_n683), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n672), .A2(G1341), .ZN(new_n686));
  NAND4_X1  g261(.A1(new_n673), .A2(new_n684), .A3(new_n685), .A4(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n669), .A2(G4), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n688), .B1(new_n584), .B2(new_n669), .ZN(new_n689));
  INV_X1    g264(.A(G1348), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(G115), .A2(G2104), .ZN(new_n692));
  INV_X1    g267(.A(G127), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n692), .B1(new_n466), .B2(new_n693), .ZN(new_n694));
  AOI22_X1  g269(.A1(new_n477), .A2(G139), .B1(new_n694), .B2(G2105), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n469), .A2(G103), .ZN(new_n696));
  XOR2_X1   g271(.A(new_n696), .B(KEYINPUT25), .Z(new_n697));
  NAND2_X1  g272(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  MUX2_X1   g273(.A(G33), .B(new_n698), .S(G29), .Z(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G2072), .ZN(new_n700));
  NOR2_X1   g275(.A1(G5), .A2(G16), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n701), .B1(G171), .B2(G16), .ZN(new_n702));
  OAI211_X1 g277(.A(new_n691), .B(new_n700), .C1(G1961), .C2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(G1956), .ZN(new_n704));
  INV_X1    g279(.A(KEYINPUT23), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(G299), .B2(G16), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n669), .A2(G20), .ZN(new_n707));
  MUX2_X1   g282(.A(new_n705), .B(new_n706), .S(new_n707), .Z(new_n708));
  AOI211_X1 g283(.A(new_n687), .B(new_n703), .C1(new_n704), .C2(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n681), .A2(G27), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(G164), .B2(new_n681), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT99), .ZN(new_n712));
  INV_X1    g287(.A(G2078), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(G2067), .ZN(new_n715));
  AND2_X1   g290(.A1(new_n681), .A2(G26), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n600), .A2(G128), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n477), .A2(G140), .ZN(new_n718));
  NOR2_X1   g293(.A1(G104), .A2(G2105), .ZN(new_n719));
  OAI21_X1  g294(.A(G2104), .B1(new_n471), .B2(G116), .ZN(new_n720));
  OAI211_X1 g295(.A(new_n717), .B(new_n718), .C1(new_n719), .C2(new_n720), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n716), .B1(new_n721), .B2(G29), .ZN(new_n722));
  MUX2_X1   g297(.A(new_n716), .B(new_n722), .S(KEYINPUT28), .Z(new_n723));
  OAI221_X1 g298(.A(new_n714), .B1(new_n704), .B2(new_n708), .C1(new_n715), .C2(new_n723), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(new_n715), .B2(new_n723), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n709), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT31), .B(G11), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT30), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(G28), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n729), .A2(KEYINPUT95), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n681), .B1(new_n728), .B2(G28), .ZN(new_n731));
  AOI22_X1  g306(.A1(new_n731), .A2(KEYINPUT96), .B1(new_n729), .B2(KEYINPUT95), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(KEYINPUT96), .B2(new_n731), .ZN(new_n733));
  OAI221_X1 g308(.A(new_n727), .B1(new_n730), .B2(new_n733), .C1(new_n606), .C2(new_n681), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT97), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n669), .A2(G21), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G168), .B2(new_n669), .ZN(new_n737));
  AOI22_X1  g312(.A1(new_n737), .A2(G1966), .B1(G1961), .B2(new_n702), .ZN(new_n738));
  OAI211_X1 g313(.A(new_n735), .B(new_n738), .C1(G1966), .C2(new_n737), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT98), .Z(new_n740));
  NAND2_X1  g315(.A1(new_n681), .A2(G35), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G162), .B2(new_n681), .ZN(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT29), .B(G2090), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT24), .ZN(new_n745));
  OR2_X1    g320(.A1(new_n745), .A2(G34), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(G34), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n746), .A2(new_n747), .A3(new_n681), .ZN(new_n748));
  INV_X1    g323(.A(G160), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n748), .B1(new_n749), .B2(new_n681), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT93), .ZN(new_n751));
  INV_X1    g326(.A(G2084), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NOR4_X1   g328(.A1(new_n726), .A2(new_n740), .A3(new_n744), .A4(new_n753), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n699), .A2(G2072), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n669), .A2(G22), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G166), .B2(new_n669), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n757), .A2(G1971), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n669), .A2(G23), .ZN(new_n759));
  INV_X1    g334(.A(G288), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n759), .B1(new_n760), .B2(new_n669), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT33), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(G1976), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n757), .A2(G1971), .ZN(new_n764));
  MUX2_X1   g339(.A(G6), .B(G305), .S(G16), .Z(new_n765));
  XOR2_X1   g340(.A(KEYINPUT32), .B(G1981), .Z(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NAND4_X1  g342(.A1(new_n758), .A2(new_n763), .A3(new_n764), .A4(new_n767), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n768), .A2(KEYINPUT34), .ZN(new_n769));
  AND2_X1   g344(.A1(new_n669), .A2(G24), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(G290), .B2(G16), .ZN(new_n771));
  INV_X1    g346(.A(G1986), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n768), .A2(KEYINPUT34), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n681), .A2(G25), .ZN(new_n775));
  INV_X1    g350(.A(G131), .ZN(new_n776));
  NOR2_X1   g351(.A1(G95), .A2(G2105), .ZN(new_n777));
  OAI21_X1  g352(.A(G2104), .B1(new_n471), .B2(G107), .ZN(new_n778));
  OAI22_X1  g353(.A1(new_n476), .A2(new_n776), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G119), .B2(new_n600), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n775), .B1(new_n780), .B2(new_n681), .ZN(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT35), .B(G1991), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(new_n771), .B2(new_n772), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n781), .A2(new_n782), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND4_X1  g361(.A1(new_n769), .A2(new_n773), .A3(new_n774), .A4(new_n786), .ZN(new_n787));
  XOR2_X1   g362(.A(KEYINPUT90), .B(KEYINPUT36), .Z(new_n788));
  OR2_X1    g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n787), .A2(KEYINPUT36), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n789), .A2(KEYINPUT91), .A3(new_n790), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n789), .A2(KEYINPUT91), .ZN(new_n792));
  NAND4_X1  g367(.A1(new_n754), .A2(new_n755), .A3(new_n791), .A4(new_n792), .ZN(G150));
  INV_X1    g368(.A(G150), .ZN(G311));
  AND2_X1   g369(.A1(new_n528), .A2(G55), .ZN(new_n795));
  AOI22_X1  g370(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n796));
  INV_X1    g371(.A(G93), .ZN(new_n797));
  OAI22_X1  g372(.A1(new_n796), .A2(new_n515), .B1(new_n522), .B2(new_n797), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n795), .A2(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  XOR2_X1   g375(.A(KEYINPUT101), .B(G860), .Z(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(KEYINPUT37), .Z(new_n803));
  NOR2_X1   g378(.A1(new_n583), .A2(new_n591), .ZN(new_n804));
  XNOR2_X1  g379(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n800), .A2(KEYINPUT100), .ZN(new_n807));
  INV_X1    g382(.A(new_n550), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT100), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n799), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n807), .A2(new_n808), .A3(new_n810), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n550), .A2(new_n799), .A3(new_n809), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n806), .B(new_n813), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n803), .B1(new_n814), .B2(new_n801), .ZN(G145));
  XNOR2_X1  g390(.A(new_n491), .B(KEYINPUT102), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(G160), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(new_n612), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n600), .A2(G130), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n477), .A2(G142), .ZN(new_n820));
  NOR2_X1   g395(.A1(G106), .A2(G2105), .ZN(new_n821));
  OAI21_X1  g396(.A(G2104), .B1(new_n471), .B2(G118), .ZN(new_n822));
  OAI211_X1 g397(.A(new_n819), .B(new_n820), .C1(new_n821), .C2(new_n822), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(new_n780), .Z(new_n824));
  XNOR2_X1  g399(.A(new_n818), .B(new_n824), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n507), .B(new_n721), .Z(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(new_n680), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n698), .A2(KEYINPUT103), .ZN(new_n828));
  AND2_X1   g403(.A1(new_n698), .A2(KEYINPUT103), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n827), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n830), .B1(new_n828), .B2(new_n827), .ZN(new_n831));
  XOR2_X1   g406(.A(new_n831), .B(new_n606), .Z(new_n832));
  XNOR2_X1  g407(.A(new_n825), .B(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT104), .ZN(new_n834));
  OR3_X1    g409(.A1(new_n833), .A2(new_n834), .A3(G37), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n834), .B1(new_n833), .B2(G37), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g413(.A(new_n813), .B(new_n594), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n583), .B(new_n588), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(KEYINPUT41), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n841), .B1(new_n839), .B2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(G305), .B(G288), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(G290), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(G166), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT42), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n843), .B(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(G868), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n849), .B1(G868), .B2(new_n799), .ZN(G295));
  OAI21_X1  g425(.A(new_n849), .B1(G868), .B2(new_n799), .ZN(G331));
  INV_X1    g426(.A(G37), .ZN(new_n852));
  XNOR2_X1  g427(.A(G286), .B(G171), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n813), .B(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(new_n840), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n855), .B1(new_n842), .B2(new_n854), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n852), .B1(new_n856), .B2(new_n846), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n857), .B1(new_n846), .B2(new_n856), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n858), .A2(KEYINPUT43), .ZN(new_n859));
  INV_X1    g434(.A(new_n846), .ZN(new_n860));
  INV_X1    g435(.A(new_n854), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT41), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n840), .A2(KEYINPUT105), .A3(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n842), .ZN(new_n864));
  OAI211_X1 g439(.A(new_n861), .B(new_n863), .C1(new_n864), .C2(KEYINPUT105), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n860), .B1(new_n865), .B2(new_n855), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT43), .ZN(new_n867));
  NOR3_X1   g442(.A1(new_n866), .A2(new_n857), .A3(new_n867), .ZN(new_n868));
  OAI21_X1  g443(.A(KEYINPUT44), .B1(new_n859), .B2(new_n868), .ZN(new_n869));
  OR2_X1    g444(.A1(new_n858), .A2(new_n867), .ZN(new_n870));
  OR3_X1    g445(.A1(new_n866), .A2(new_n857), .A3(KEYINPUT43), .ZN(new_n871));
  AND2_X1   g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n869), .B1(new_n872), .B2(KEYINPUT44), .ZN(G397));
  NAND2_X1  g448(.A1(G303), .A2(G8), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT55), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(G1384), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n499), .B1(new_n495), .B2(KEYINPUT4), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n877), .B1(new_n878), .B2(new_n505), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT45), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n470), .A2(G40), .A3(new_n478), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  OAI211_X1 g458(.A(KEYINPUT45), .B(new_n877), .C1(new_n878), .C2(new_n505), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n881), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(G1971), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n879), .A2(KEYINPUT50), .ZN(new_n888));
  XOR2_X1   g463(.A(KEYINPUT108), .B(KEYINPUT50), .Z(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  OAI211_X1 g465(.A(new_n877), .B(new_n890), .C1(new_n878), .C2(new_n505), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n888), .A2(new_n883), .A3(new_n891), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n887), .B1(G2090), .B2(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(KEYINPUT109), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n876), .A2(G8), .A3(new_n894), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n879), .A2(new_n882), .ZN(new_n896));
  INV_X1    g471(.A(G8), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(G1976), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n898), .B1(new_n899), .B2(G288), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT52), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n901), .B1(new_n760), .B2(G1976), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  AND2_X1   g478(.A1(new_n900), .A2(KEYINPUT52), .ZN(new_n904));
  XNOR2_X1  g479(.A(G305), .B(G1981), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT49), .ZN(new_n906));
  AND2_X1   g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n898), .B1(new_n905), .B2(new_n906), .ZN(new_n908));
  OR3_X1    g483(.A1(new_n907), .A2(new_n908), .A3(KEYINPUT110), .ZN(new_n909));
  OAI21_X1  g484(.A(KEYINPUT110), .B1(new_n907), .B2(new_n908), .ZN(new_n910));
  AOI211_X1 g485(.A(new_n903), .B(new_n904), .C1(new_n909), .C2(new_n910), .ZN(new_n911));
  AND2_X1   g486(.A1(new_n895), .A2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n879), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n913), .A2(new_n890), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n883), .B1(new_n879), .B2(KEYINPUT50), .ZN(new_n915));
  NOR3_X1   g490(.A1(new_n914), .A2(new_n915), .A3(G2090), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n916), .B1(new_n886), .B2(new_n885), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n875), .B1(new_n897), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n912), .A2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT61), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT57), .ZN(new_n921));
  XNOR2_X1  g496(.A(G299), .B(new_n921), .ZN(new_n922));
  XNOR2_X1  g497(.A(KEYINPUT56), .B(G2072), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n881), .A2(new_n883), .A3(new_n884), .A4(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT114), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n924), .B(new_n925), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n704), .B1(new_n914), .B2(new_n915), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n922), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  AND2_X1   g503(.A1(new_n881), .A2(new_n884), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n929), .A2(new_n925), .A3(new_n883), .A4(new_n923), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n924), .A2(KEYINPUT114), .ZN(new_n931));
  AND4_X1   g506(.A1(new_n922), .A2(new_n930), .A3(new_n927), .A4(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n920), .B1(new_n928), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n892), .A2(new_n690), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n896), .A2(KEYINPUT115), .A3(new_n715), .ZN(new_n935));
  AND2_X1   g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n896), .A2(new_n715), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT115), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n583), .B1(new_n936), .B2(new_n939), .ZN(new_n940));
  AND4_X1   g515(.A1(new_n583), .A2(new_n939), .A3(new_n934), .A4(new_n935), .ZN(new_n941));
  OAI21_X1  g516(.A(KEYINPUT60), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n930), .A2(new_n927), .A3(new_n931), .ZN(new_n943));
  INV_X1    g518(.A(new_n922), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n922), .A2(new_n930), .A3(new_n927), .A4(new_n931), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n945), .A2(KEYINPUT61), .A3(new_n946), .ZN(new_n947));
  XNOR2_X1  g522(.A(KEYINPUT58), .B(G1341), .ZN(new_n948));
  OAI22_X1  g523(.A1(new_n885), .A2(G1996), .B1(new_n896), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(new_n550), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(KEYINPUT59), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT59), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n949), .A2(new_n952), .A3(new_n550), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT60), .ZN(new_n954));
  AND4_X1   g529(.A1(new_n954), .A2(new_n934), .A3(new_n939), .A4(new_n935), .ZN(new_n955));
  AOI22_X1  g530(.A1(new_n951), .A2(new_n953), .B1(new_n955), .B2(new_n584), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n933), .A2(new_n942), .A3(new_n947), .A4(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n940), .A2(new_n946), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n957), .A2(new_n958), .A3(new_n945), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n929), .A2(new_n713), .A3(new_n883), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT53), .ZN(new_n961));
  INV_X1    g536(.A(G1961), .ZN(new_n962));
  AOI22_X1  g537(.A1(new_n960), .A2(new_n961), .B1(new_n962), .B2(new_n892), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT124), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT122), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n470), .A2(new_n478), .A3(new_n965), .A4(G40), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n882), .A2(KEYINPUT122), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n881), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n961), .B1(new_n968), .B2(KEYINPUT123), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT123), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n881), .A2(new_n970), .A3(new_n967), .A4(new_n966), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n969), .A2(new_n713), .A3(new_n884), .A4(new_n971), .ZN(new_n972));
  AND3_X1   g547(.A1(new_n963), .A2(new_n964), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n964), .B1(new_n963), .B2(new_n972), .ZN(new_n974));
  NOR3_X1   g549(.A1(new_n973), .A2(new_n974), .A3(G301), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n885), .A2(G2078), .ZN(new_n976));
  OR2_X1    g551(.A1(new_n976), .A2(KEYINPUT121), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n976), .A2(KEYINPUT121), .A3(KEYINPUT53), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n963), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(G301), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(KEYINPUT54), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n979), .A2(G171), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT54), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  AND3_X1   g559(.A1(new_n963), .A2(G301), .A3(new_n972), .ZN(new_n985));
  OAI22_X1  g560(.A1(new_n975), .A2(new_n981), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  AND2_X1   g561(.A1(new_n959), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(G1966), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n885), .A2(new_n988), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n888), .A2(new_n752), .A3(new_n883), .A4(new_n891), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT117), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n991), .A2(new_n992), .A3(G8), .ZN(new_n993));
  NAND2_X1  g568(.A1(G286), .A2(G8), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n897), .B1(new_n989), .B2(new_n990), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n996), .A2(new_n992), .ZN(new_n997));
  OAI21_X1  g572(.A(KEYINPUT51), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT118), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT51), .ZN(new_n1001));
  INV_X1    g576(.A(new_n892), .ZN(new_n1002));
  AOI22_X1  g577(.A1(new_n1002), .A2(new_n752), .B1(new_n885), .B2(new_n988), .ZN(new_n1003));
  OAI211_X1 g578(.A(new_n1001), .B(new_n994), .C1(new_n1003), .C2(new_n897), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT119), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n996), .A2(KEYINPUT51), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1007), .A2(KEYINPUT119), .A3(new_n994), .ZN(new_n1008));
  AND2_X1   g583(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  AOI22_X1  g584(.A1(new_n996), .A2(new_n992), .B1(G8), .B2(G286), .ZN(new_n1010));
  OAI21_X1  g585(.A(KEYINPUT117), .B1(new_n1003), .B2(new_n897), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1001), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(KEYINPUT118), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1000), .A2(new_n1009), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT120), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1003), .A2(new_n994), .ZN(new_n1016));
  XOR2_X1   g591(.A(new_n1016), .B(KEYINPUT116), .Z(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  AND3_X1   g593(.A1(new_n1014), .A2(new_n1015), .A3(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1015), .B1(new_n1014), .B2(new_n1018), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n987), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n996), .A2(G168), .ZN(new_n1022));
  XNOR2_X1  g597(.A(new_n1022), .B(KEYINPUT113), .ZN(new_n1023));
  AND3_X1   g598(.A1(new_n895), .A2(new_n911), .A3(KEYINPUT63), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n894), .A2(G8), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(new_n875), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1023), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n919), .B1(new_n1021), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1023), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1024), .A2(new_n1030), .A3(new_n1026), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(KEYINPUT63), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n904), .B1(new_n909), .B2(new_n910), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1033), .B1(new_n900), .B2(new_n902), .ZN(new_n1034));
  OR2_X1    g609(.A1(new_n1034), .A2(new_n895), .ZN(new_n1035));
  AOI211_X1 g610(.A(G1976), .B(G288), .C1(new_n909), .C2(new_n910), .ZN(new_n1036));
  NOR2_X1   g611(.A1(G305), .A2(G1981), .ZN(new_n1037));
  XNOR2_X1  g612(.A(new_n1037), .B(KEYINPUT111), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n898), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1035), .A2(KEYINPUT112), .A3(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(KEYINPUT112), .B1(new_n1035), .B2(new_n1039), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1032), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g618(.A(KEYINPUT125), .B1(new_n1029), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT125), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1035), .A2(new_n1039), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT112), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  AOI22_X1  g623(.A1(new_n1048), .A2(new_n1040), .B1(new_n1031), .B2(KEYINPUT63), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1012), .A2(KEYINPUT118), .ZN(new_n1050));
  AOI211_X1 g625(.A(new_n999), .B(new_n1001), .C1(new_n1010), .C2(new_n1011), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1052));
  NOR3_X1   g627(.A1(new_n1050), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  OAI21_X1  g628(.A(KEYINPUT120), .B1(new_n1053), .B2(new_n1017), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1014), .A2(new_n1015), .A3(new_n1018), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1027), .B1(new_n1056), .B2(new_n987), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n1045), .B(new_n1049), .C1(new_n1057), .C2(new_n919), .ZN(new_n1058));
  OAI21_X1  g633(.A(KEYINPUT62), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT62), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1054), .A2(new_n1060), .A3(new_n1055), .ZN(new_n1061));
  INV_X1    g636(.A(new_n919), .ZN(new_n1062));
  INV_X1    g637(.A(new_n982), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1059), .A2(new_n1061), .A3(new_n1062), .A4(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT126), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n919), .B1(new_n1056), .B2(KEYINPUT62), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1067), .A2(KEYINPUT126), .A3(new_n1063), .A4(new_n1061), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1044), .A2(new_n1058), .A3(new_n1066), .A4(new_n1068), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n881), .A2(new_n882), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1070), .ZN(new_n1071));
  OR2_X1    g646(.A1(new_n1071), .A2(G1996), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1072), .A2(new_n680), .ZN(new_n1073));
  XOR2_X1   g648(.A(new_n1073), .B(KEYINPUT106), .Z(new_n1074));
  XNOR2_X1  g649(.A(new_n1070), .B(KEYINPUT107), .ZN(new_n1075));
  AND2_X1   g650(.A1(new_n1075), .A2(new_n680), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(G1996), .ZN(new_n1077));
  XNOR2_X1  g652(.A(new_n721), .B(G2067), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1075), .A2(new_n1078), .ZN(new_n1079));
  AND3_X1   g654(.A1(new_n1074), .A2(new_n1077), .A3(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(new_n782), .ZN(new_n1081));
  XNOR2_X1  g656(.A(new_n780), .B(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1075), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1080), .A2(new_n1083), .ZN(new_n1084));
  XNOR2_X1  g659(.A(G290), .B(G1986), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1084), .B1(new_n1070), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1069), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT46), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1076), .B1(new_n1088), .B2(new_n1072), .ZN(new_n1089));
  OAI211_X1 g664(.A(new_n1089), .B(new_n1079), .C1(new_n1088), .C2(new_n1072), .ZN(new_n1090));
  XOR2_X1   g665(.A(new_n1090), .B(KEYINPUT47), .Z(new_n1091));
  AND2_X1   g666(.A1(new_n1084), .A2(KEYINPUT127), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1084), .A2(KEYINPUT127), .ZN(new_n1093));
  OR3_X1    g668(.A1(new_n1071), .A2(G1986), .A3(G290), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT48), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  AND2_X1   g671(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1097));
  NOR4_X1   g672(.A1(new_n1092), .A2(new_n1093), .A3(new_n1096), .A4(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1080), .A2(new_n1081), .A3(new_n780), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1099), .B1(G2067), .B2(new_n721), .ZN(new_n1100));
  AOI211_X1 g675(.A(new_n1091), .B(new_n1098), .C1(new_n1075), .C2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1087), .A2(new_n1101), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g677(.A(G319), .ZN(new_n1104));
  OR2_X1    g678(.A1(G227), .A2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g679(.A(new_n1105), .B1(new_n870), .B2(new_n871), .ZN(new_n1106));
  NOR2_X1   g680(.A1(G229), .A2(G401), .ZN(new_n1107));
  AND3_X1   g681(.A1(new_n1106), .A2(new_n837), .A3(new_n1107), .ZN(G308));
  NAND3_X1  g682(.A1(new_n1106), .A2(new_n837), .A3(new_n1107), .ZN(G225));
endmodule


