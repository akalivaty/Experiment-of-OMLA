

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792;

  INV_X1 U379 ( .A(G478), .ZN(n357) );
  XNOR2_X2 U380 ( .A(n358), .B(n357), .ZN(n587) );
  OR2_X2 U381 ( .A1(n746), .A2(G902), .ZN(n358) );
  XNOR2_X1 U382 ( .A(n550), .B(n401), .ZN(n400) );
  NAND2_X2 U383 ( .A1(n759), .A2(n473), .ZN(n471) );
  OR2_X2 U384 ( .A1(n689), .A2(n592), .ZN(n377) );
  INV_X2 U385 ( .A(KEYINPUT4), .ZN(n421) );
  AND2_X2 U386 ( .A1(n576), .A2(n371), .ZN(n366) );
  XNOR2_X2 U387 ( .A(n378), .B(n426), .ZN(n792) );
  XNOR2_X2 U388 ( .A(n549), .B(n538), .ZN(n774) );
  XNOR2_X2 U389 ( .A(n553), .B(G134), .ZN(n549) );
  AND2_X2 U390 ( .A1(n789), .A2(KEYINPUT68), .ZN(n633) );
  NOR2_X1 U391 ( .A1(G953), .A2(G237), .ZN(n537) );
  XNOR2_X2 U392 ( .A(n632), .B(n631), .ZN(n789) );
  OR2_X2 U393 ( .A1(n731), .A2(n730), .ZN(n440) );
  AND2_X1 U394 ( .A1(n695), .A2(n454), .ZN(n453) );
  NOR2_X1 U395 ( .A1(n735), .A2(n754), .ZN(n409) );
  XNOR2_X1 U396 ( .A(n377), .B(n570), .ZN(n787) );
  NOR2_X1 U397 ( .A1(n388), .A2(n389), .ZN(n434) );
  AND2_X1 U398 ( .A1(n416), .A2(n413), .ZN(n389) );
  XNOR2_X1 U399 ( .A(n545), .B(n544), .ZN(n588) );
  XNOR2_X1 U400 ( .A(n774), .B(G146), .ZN(n498) );
  XNOR2_X1 U401 ( .A(n533), .B(n380), .ZN(n379) );
  INV_X2 U402 ( .A(KEYINPUT3), .ZN(n420) );
  XNOR2_X1 U403 ( .A(KEYINPUT8), .B(KEYINPUT69), .ZN(n514) );
  XNOR2_X1 U404 ( .A(G113), .B(G104), .ZN(n533) );
  AND2_X2 U405 ( .A1(n471), .A2(n472), .ZN(n359) );
  XNOR2_X1 U406 ( .A(n780), .B(KEYINPUT74), .ZN(n360) );
  AND2_X1 U407 ( .A1(n455), .A2(n453), .ZN(n452) );
  NAND2_X1 U408 ( .A1(n419), .A2(n621), .ZN(n648) );
  INV_X1 U409 ( .A(n621), .ZN(n361) );
  NOR2_X1 U410 ( .A1(n745), .A2(n754), .ZN(n410) );
  NOR2_X1 U411 ( .A1(n662), .A2(n754), .ZN(n663) );
  XNOR2_X1 U412 ( .A(n780), .B(KEYINPUT74), .ZN(n375) );
  OR2_X1 U413 ( .A1(G237), .A2(G902), .ZN(n568) );
  XNOR2_X1 U414 ( .A(n387), .B(n386), .ZN(n381) );
  INV_X1 U415 ( .A(KEYINPUT101), .ZN(n386) );
  INV_X1 U416 ( .A(G122), .ZN(n380) );
  OR2_X1 U417 ( .A1(n591), .A2(n468), .ZN(n460) );
  AND2_X1 U418 ( .A1(n466), .A2(n462), .ZN(n461) );
  XNOR2_X1 U419 ( .A(n376), .B(n575), .ZN(n599) );
  NOR2_X1 U420 ( .A1(n792), .A2(n787), .ZN(n376) );
  AND2_X1 U421 ( .A1(n473), .A2(n457), .ZN(n422) );
  INV_X1 U422 ( .A(KEYINPUT48), .ZN(n600) );
  INV_X1 U423 ( .A(KEYINPUT44), .ZN(n635) );
  XNOR2_X1 U424 ( .A(G146), .B(G125), .ZN(n564) );
  XOR2_X1 U425 ( .A(G107), .B(KEYINPUT76), .Z(n487) );
  XNOR2_X1 U426 ( .A(n691), .B(n403), .ZN(n402) );
  INV_X1 U427 ( .A(KEYINPUT85), .ZN(n403) );
  XNOR2_X1 U428 ( .A(n565), .B(n567), .ZN(n476) );
  XOR2_X1 U429 ( .A(G116), .B(G107), .Z(n554) );
  XOR2_X1 U430 ( .A(KEYINPUT24), .B(KEYINPUT84), .Z(n508) );
  XNOR2_X1 U431 ( .A(n554), .B(KEYINPUT7), .ZN(n401) );
  XNOR2_X1 U432 ( .A(n369), .B(n379), .ZN(n407) );
  XNOR2_X1 U433 ( .A(G143), .B(G140), .ZN(n534) );
  XOR2_X1 U434 ( .A(KEYINPUT98), .B(KEYINPUT11), .Z(n535) );
  XNOR2_X1 U435 ( .A(n373), .B(n571), .ZN(n372) );
  AND2_X1 U436 ( .A1(n707), .A2(n572), .ZN(n371) );
  NOR2_X1 U437 ( .A1(G902), .A2(n742), .ZN(n545) );
  INV_X1 U438 ( .A(G475), .ZN(n542) );
  NAND2_X1 U439 ( .A1(n587), .A2(n588), .ZN(n589) );
  INV_X1 U440 ( .A(G953), .ZN(n437) );
  NOR2_X1 U441 ( .A1(n629), .A2(n468), .ZN(n464) );
  NAND2_X1 U442 ( .A1(n461), .A2(n459), .ZN(n595) );
  BUF_X1 U443 ( .A(n721), .Z(n411) );
  XNOR2_X1 U444 ( .A(G902), .B(KEYINPUT15), .ZN(n485) );
  XOR2_X1 U445 ( .A(KEYINPUT5), .B(KEYINPUT72), .Z(n501) );
  XOR2_X1 U446 ( .A(KEYINPUT96), .B(G137), .Z(n496) );
  NAND2_X1 U447 ( .A1(n450), .A2(KEYINPUT65), .ZN(n449) );
  INV_X1 U448 ( .A(n695), .ZN(n450) );
  NAND2_X1 U449 ( .A1(G234), .A2(G237), .ZN(n523) );
  INV_X1 U450 ( .A(G472), .ZN(n458) );
  XNOR2_X1 U451 ( .A(n442), .B(n600), .ZN(n441) );
  AND2_X1 U452 ( .A1(n397), .A2(n653), .ZN(n654) );
  XNOR2_X1 U453 ( .A(n490), .B(n489), .ZN(n491) );
  NOR2_X1 U454 ( .A1(n394), .A2(n586), .ZN(n431) );
  NAND2_X1 U455 ( .A1(n429), .A2(KEYINPUT34), .ZN(n428) );
  XNOR2_X1 U456 ( .A(KEYINPUT22), .B(KEYINPUT71), .ZN(n618) );
  INV_X1 U457 ( .A(KEYINPUT19), .ZN(n474) );
  AND2_X1 U458 ( .A1(n522), .A2(n374), .ZN(n707) );
  XNOR2_X1 U459 ( .A(n557), .B(n556), .ZN(n764) );
  XNOR2_X1 U460 ( .A(n512), .B(n382), .ZN(n752) );
  XOR2_X1 U461 ( .A(KEYINPUT9), .B(KEYINPUT100), .Z(n548) );
  XNOR2_X1 U462 ( .A(n541), .B(n540), .ZN(n742) );
  NOR2_X1 U463 ( .A1(G952), .A2(n437), .ZN(n754) );
  XNOR2_X1 U464 ( .A(n574), .B(n427), .ZN(n426) );
  OR2_X2 U465 ( .A1(n601), .A2(n589), .ZN(n378) );
  INV_X1 U466 ( .A(KEYINPUT105), .ZN(n427) );
  XNOR2_X1 U467 ( .A(n646), .B(n404), .ZN(n683) );
  XNOR2_X1 U468 ( .A(n405), .B(KEYINPUT31), .ZN(n404) );
  INV_X1 U469 ( .A(KEYINPUT97), .ZN(n405) );
  INV_X1 U470 ( .A(KEYINPUT53), .ZN(n435) );
  XNOR2_X1 U471 ( .A(n644), .B(n418), .ZN(n627) );
  AND2_X1 U472 ( .A1(n707), .A2(KEYINPUT33), .ZN(n362) );
  AND2_X1 U473 ( .A1(n444), .A2(KEYINPUT65), .ZN(n363) );
  AND2_X1 U474 ( .A1(n677), .A2(n597), .ZN(n364) );
  NOR2_X1 U475 ( .A1(n704), .A2(n649), .ZN(n365) );
  OR2_X1 U476 ( .A1(n470), .A2(n395), .ZN(n367) );
  AND2_X1 U477 ( .A1(n788), .A2(n608), .ZN(n368) );
  NAND2_X1 U478 ( .A1(G214), .A2(n537), .ZN(n369) );
  INV_X1 U479 ( .A(KEYINPUT34), .ZN(n628) );
  INV_X1 U480 ( .A(KEYINPUT33), .ZN(n417) );
  INV_X1 U481 ( .A(KEYINPUT66), .ZN(n457) );
  INV_X1 U482 ( .A(KEYINPUT2), .ZN(n473) );
  XOR2_X1 U483 ( .A(n484), .B(n483), .Z(n370) );
  NAND2_X1 U484 ( .A1(n576), .A2(n707), .ZN(n642) );
  INV_X1 U485 ( .A(n522), .ZN(n700) );
  AND2_X2 U486 ( .A1(n366), .A2(n372), .ZN(n584) );
  NAND2_X1 U487 ( .A1(n704), .A2(n717), .ZN(n373) );
  INV_X1 U488 ( .A(n699), .ZN(n374) );
  NAND2_X1 U489 ( .A1(n360), .A2(n422), .ZN(n444) );
  AND2_X2 U490 ( .A1(n375), .A2(n473), .ZN(n470) );
  XNOR2_X1 U491 ( .A(n379), .B(n554), .ZN(n557) );
  NOR2_X1 U492 ( .A1(n381), .A2(n699), .ZN(n609) );
  NOR2_X1 U493 ( .A1(n720), .A2(n381), .ZN(n569) );
  NOR2_X1 U494 ( .A1(n719), .A2(n381), .ZN(n723) );
  XNOR2_X1 U495 ( .A(n407), .B(n536), .ZN(n541) );
  XOR2_X1 U496 ( .A(n516), .B(n513), .Z(n382) );
  NAND2_X1 U497 ( .A1(n367), .A2(n446), .ZN(n445) );
  AND2_X1 U498 ( .A1(n363), .A2(n456), .ZN(n446) );
  NOR2_X1 U499 ( .A1(n667), .A2(n683), .ZN(n647) );
  OR2_X1 U500 ( .A1(n591), .A2(n464), .ZN(n463) );
  NAND2_X1 U501 ( .A1(n591), .A2(KEYINPUT80), .ZN(n465) );
  XNOR2_X1 U502 ( .A(n596), .B(KEYINPUT82), .ZN(n408) );
  XNOR2_X1 U503 ( .A(KEYINPUT83), .B(n590), .ZN(n591) );
  BUF_X1 U504 ( .A(n645), .Z(n383) );
  XNOR2_X1 U505 ( .A(n503), .B(n497), .ZN(n398) );
  NOR2_X1 U506 ( .A1(n388), .A2(n389), .ZN(n384) );
  XNOR2_X2 U507 ( .A(n494), .B(n493), .ZN(n385) );
  XNOR2_X1 U508 ( .A(n494), .B(n493), .ZN(n576) );
  XNOR2_X1 U509 ( .A(n739), .B(n738), .ZN(n740) );
  NAND2_X1 U510 ( .A1(n583), .A2(n587), .ZN(n387) );
  XNOR2_X1 U511 ( .A(n564), .B(n563), .ZN(n479) );
  NAND2_X1 U512 ( .A1(n414), .A2(n415), .ZN(n388) );
  NOR2_X2 U513 ( .A1(n737), .A2(G902), .ZN(n494) );
  BUF_X1 U514 ( .A(n732), .Z(n390) );
  XNOR2_X1 U515 ( .A(n477), .B(n764), .ZN(n732) );
  BUF_X1 U516 ( .A(n741), .Z(n750) );
  BUF_X1 U517 ( .A(n789), .Z(n391) );
  INV_X1 U518 ( .A(n580), .ZN(n392) );
  INV_X2 U519 ( .A(n607), .ZN(n580) );
  XNOR2_X1 U520 ( .A(G113), .B(G116), .ZN(n495) );
  BUF_X1 U521 ( .A(n774), .Z(n393) );
  XNOR2_X1 U522 ( .A(G128), .B(KEYINPUT23), .ZN(n507) );
  NOR2_X1 U523 ( .A1(n682), .A2(n679), .ZN(n721) );
  NOR2_X1 U524 ( .A1(n645), .A2(n628), .ZN(n394) );
  NAND2_X1 U525 ( .A1(n359), .A2(KEYINPUT66), .ZN(n395) );
  XNOR2_X1 U526 ( .A(n562), .B(n479), .ZN(n478) );
  NOR2_X1 U527 ( .A1(n395), .A2(n470), .ZN(n455) );
  NAND2_X1 U528 ( .A1(n444), .A2(n456), .ZN(n425) );
  NAND2_X1 U529 ( .A1(n424), .A2(n423), .ZN(n695) );
  XNOR2_X1 U530 ( .A(n475), .B(n474), .ZN(n616) );
  XNOR2_X1 U531 ( .A(n737), .B(n736), .ZN(n738) );
  NOR2_X1 U532 ( .A1(n759), .A2(n473), .ZN(n424) );
  AND2_X1 U533 ( .A1(n706), .A2(n362), .ZN(n413) );
  XNOR2_X1 U534 ( .A(n478), .B(n561), .ZN(n477) );
  XNOR2_X2 U535 ( .A(n399), .B(n499), .ZN(n562) );
  INV_X1 U536 ( .A(n658), .ZN(n472) );
  BUF_X1 U537 ( .A(n429), .Z(n396) );
  NAND2_X1 U538 ( .A1(n640), .A2(n671), .ZN(n397) );
  XNOR2_X2 U539 ( .A(n626), .B(n625), .ZN(n791) );
  INV_X1 U540 ( .A(n627), .ZN(n416) );
  XNOR2_X1 U541 ( .A(n398), .B(n498), .ZN(n659) );
  NAND2_X1 U542 ( .A1(n643), .A2(n417), .ZN(n414) );
  INV_X1 U543 ( .A(n762), .ZN(n399) );
  XNOR2_X2 U544 ( .A(n421), .B(G101), .ZN(n499) );
  XNOR2_X1 U545 ( .A(n400), .B(n551), .ZN(n746) );
  NAND2_X1 U546 ( .A1(n451), .A2(n449), .ZN(n448) );
  NAND2_X1 U547 ( .A1(n471), .A2(n472), .ZN(n412) );
  XNOR2_X1 U548 ( .A(n492), .B(n491), .ZN(n737) );
  NOR2_X1 U549 ( .A1(n643), .A2(n644), .ZN(n713) );
  NAND2_X1 U550 ( .A1(n402), .A2(n693), .ZN(n694) );
  XNOR2_X2 U551 ( .A(n657), .B(n656), .ZN(n759) );
  NAND2_X1 U552 ( .A1(n406), .A2(n645), .ZN(n619) );
  XNOR2_X1 U553 ( .A(n609), .B(KEYINPUT102), .ZN(n406) );
  XNOR2_X1 U554 ( .A(n661), .B(n660), .ZN(n662) );
  NOR2_X1 U555 ( .A1(n408), .A2(n685), .ZN(n598) );
  XNOR2_X1 U556 ( .A(n409), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U557 ( .A(n410), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U558 ( .A1(n465), .A2(n463), .ZN(n462) );
  NAND2_X1 U559 ( .A1(n412), .A2(n457), .ZN(n456) );
  NAND2_X1 U560 ( .A1(n706), .A2(n707), .ZN(n643) );
  NAND2_X1 U561 ( .A1(n627), .A2(n417), .ZN(n415) );
  INV_X1 U562 ( .A(KEYINPUT6), .ZN(n418) );
  NAND2_X1 U563 ( .A1(n624), .A2(n419), .ZN(n625) );
  XNOR2_X2 U564 ( .A(n619), .B(n618), .ZN(n419) );
  XNOR2_X2 U565 ( .A(n420), .B(G119), .ZN(n762) );
  NAND2_X1 U566 ( .A1(n453), .A2(n425), .ZN(n451) );
  INV_X1 U567 ( .A(n780), .ZN(n423) );
  XNOR2_X2 U568 ( .A(n573), .B(KEYINPUT39), .ZN(n601) );
  NAND2_X2 U569 ( .A1(n430), .A2(n428), .ZN(n632) );
  INV_X1 U570 ( .A(n384), .ZN(n429) );
  AND2_X2 U571 ( .A1(n432), .A2(n431), .ZN(n430) );
  NAND2_X1 U572 ( .A1(n434), .A2(n433), .ZN(n432) );
  AND2_X1 U573 ( .A1(n645), .A2(n628), .ZN(n433) );
  XNOR2_X1 U574 ( .A(n436), .B(n435), .ZN(G75) );
  NAND2_X1 U575 ( .A1(n438), .A2(n437), .ZN(n436) );
  XNOR2_X1 U576 ( .A(n440), .B(n439), .ZN(n438) );
  INV_X1 U577 ( .A(KEYINPUT118), .ZN(n439) );
  NAND2_X1 U578 ( .A1(n607), .A2(n717), .ZN(n475) );
  XNOR2_X2 U579 ( .A(G143), .B(G128), .ZN(n553) );
  NAND2_X2 U580 ( .A1(n441), .A2(n368), .ZN(n780) );
  NAND2_X1 U581 ( .A1(n443), .A2(n598), .ZN(n442) );
  NOR2_X1 U582 ( .A1(n599), .A2(n364), .ZN(n443) );
  NAND2_X2 U583 ( .A1(n447), .A2(n445), .ZN(n741) );
  NOR2_X2 U584 ( .A1(n452), .A2(n448), .ZN(n447) );
  INV_X1 U585 ( .A(KEYINPUT65), .ZN(n454) );
  INV_X1 U586 ( .A(n704), .ZN(n644) );
  XNOR2_X2 U587 ( .A(n504), .B(n458), .ZN(n704) );
  AND2_X1 U588 ( .A1(n469), .A2(n629), .ZN(n675) );
  OR2_X1 U589 ( .A1(n469), .A2(n460), .ZN(n459) );
  NAND2_X1 U590 ( .A1(n469), .A2(n467), .ZN(n466) );
  AND2_X1 U591 ( .A1(n629), .A2(n468), .ZN(n467) );
  INV_X1 U592 ( .A(KEYINPUT80), .ZN(n468) );
  XNOR2_X1 U593 ( .A(n585), .B(KEYINPUT104), .ZN(n469) );
  XNOR2_X1 U594 ( .A(n663), .B(n370), .ZN(G57) );
  XNOR2_X2 U595 ( .A(n566), .B(n476), .ZN(n607) );
  XNOR2_X1 U596 ( .A(n636), .B(n635), .ZN(n655) );
  AND2_X2 U597 ( .A1(n620), .A2(n365), .ZN(n637) );
  NOR2_X2 U598 ( .A1(n616), .A2(n615), .ZN(n617) );
  XOR2_X1 U599 ( .A(G119), .B(G110), .Z(n480) );
  XNOR2_X1 U600 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n481) );
  XNOR2_X1 U601 ( .A(KEYINPUT119), .B(KEYINPUT59), .ZN(n482) );
  XNOR2_X1 U602 ( .A(n562), .B(n502), .ZN(n503) );
  XNOR2_X1 U603 ( .A(n480), .B(n510), .ZN(n511) );
  INV_X1 U604 ( .A(G469), .ZN(n493) );
  XNOR2_X1 U605 ( .A(n770), .B(n511), .ZN(n512) );
  XNOR2_X1 U606 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U607 ( .A(n742), .B(n482), .ZN(n743) );
  XNOR2_X1 U608 ( .A(n746), .B(KEYINPUT120), .ZN(n747) );
  XNOR2_X1 U609 ( .A(n630), .B(KEYINPUT35), .ZN(n631) );
  XNOR2_X1 U610 ( .A(n748), .B(n747), .ZN(n749) );
  XOR2_X1 U611 ( .A(KEYINPUT88), .B(KEYINPUT108), .Z(n484) );
  XNOR2_X1 U612 ( .A(KEYINPUT89), .B(KEYINPUT63), .ZN(n483) );
  XNOR2_X1 U613 ( .A(n485), .B(KEYINPUT90), .ZN(n658) );
  XOR2_X1 U614 ( .A(KEYINPUT106), .B(KEYINPUT42), .Z(n570) );
  XOR2_X1 U615 ( .A(G131), .B(KEYINPUT70), .Z(n538) );
  XNOR2_X1 U616 ( .A(n498), .B(G104), .ZN(n492) );
  INV_X2 U617 ( .A(G953), .ZN(n783) );
  NAND2_X1 U618 ( .A1(G227), .A2(n783), .ZN(n486) );
  XNOR2_X1 U619 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U620 ( .A(G137), .B(G140), .ZN(n509) );
  XNOR2_X1 U621 ( .A(KEYINPUT95), .B(n509), .ZN(n769) );
  XOR2_X1 U622 ( .A(n488), .B(n769), .Z(n490) );
  XOR2_X1 U623 ( .A(KEYINPUT73), .B(G110), .Z(n555) );
  XNOR2_X1 U624 ( .A(n499), .B(n555), .ZN(n489) );
  XNOR2_X1 U625 ( .A(n496), .B(n495), .ZN(n497) );
  NAND2_X1 U626 ( .A1(n537), .A2(G210), .ZN(n500) );
  XNOR2_X1 U627 ( .A(n501), .B(n500), .ZN(n502) );
  NOR2_X1 U628 ( .A1(n659), .A2(G902), .ZN(n504) );
  NAND2_X1 U629 ( .A1(n658), .A2(G234), .ZN(n505) );
  XNOR2_X1 U630 ( .A(KEYINPUT20), .B(n505), .ZN(n517) );
  NAND2_X1 U631 ( .A1(G221), .A2(n517), .ZN(n506) );
  XNOR2_X1 U632 ( .A(n506), .B(KEYINPUT21), .ZN(n699) );
  XNOR2_X1 U633 ( .A(n508), .B(n507), .ZN(n513) );
  XNOR2_X1 U634 ( .A(KEYINPUT10), .B(n564), .ZN(n770) );
  INV_X1 U635 ( .A(n509), .ZN(n510) );
  NAND2_X1 U636 ( .A1(n783), .A2(G234), .ZN(n515) );
  XNOR2_X1 U637 ( .A(n515), .B(n514), .ZN(n546) );
  NAND2_X1 U638 ( .A1(G221), .A2(n546), .ZN(n516) );
  NOR2_X1 U639 ( .A1(G902), .A2(n752), .ZN(n521) );
  XOR2_X1 U640 ( .A(KEYINPUT25), .B(KEYINPUT75), .Z(n519) );
  NAND2_X1 U641 ( .A1(G217), .A2(n517), .ZN(n518) );
  XNOR2_X1 U642 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U643 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U644 ( .A(n523), .B(KEYINPUT14), .ZN(n526) );
  NAND2_X1 U645 ( .A1(n526), .A2(G952), .ZN(n524) );
  XNOR2_X1 U646 ( .A(n524), .B(KEYINPUT92), .ZN(n729) );
  NOR2_X1 U647 ( .A1(G953), .A2(n729), .ZN(n525) );
  XOR2_X1 U648 ( .A(KEYINPUT93), .B(n525), .Z(n614) );
  INV_X1 U649 ( .A(n614), .ZN(n529) );
  NAND2_X1 U650 ( .A1(G902), .A2(n526), .ZN(n610) );
  NOR2_X1 U651 ( .A1(G900), .A2(n610), .ZN(n527) );
  NAND2_X1 U652 ( .A1(G953), .A2(n527), .ZN(n528) );
  NAND2_X1 U653 ( .A1(n529), .A2(n528), .ZN(n572) );
  NAND2_X1 U654 ( .A1(n700), .A2(n572), .ZN(n530) );
  NOR2_X1 U655 ( .A1(n699), .A2(n530), .ZN(n577) );
  AND2_X1 U656 ( .A1(n704), .A2(n577), .ZN(n531) );
  XNOR2_X1 U657 ( .A(KEYINPUT28), .B(n531), .ZN(n532) );
  NAND2_X1 U658 ( .A1(n385), .A2(n532), .ZN(n592) );
  XNOR2_X1 U659 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U660 ( .A(n538), .B(KEYINPUT12), .ZN(n539) );
  XNOR2_X1 U661 ( .A(n539), .B(n770), .ZN(n540) );
  XNOR2_X1 U662 ( .A(KEYINPUT13), .B(KEYINPUT99), .ZN(n543) );
  INV_X1 U663 ( .A(n588), .ZN(n583) );
  NAND2_X1 U664 ( .A1(G217), .A2(n546), .ZN(n547) );
  XNOR2_X1 U665 ( .A(n548), .B(n547), .ZN(n551) );
  XNOR2_X1 U666 ( .A(n549), .B(G122), .ZN(n550) );
  INV_X1 U667 ( .A(n553), .ZN(n563) );
  XNOR2_X1 U668 ( .A(KEYINPUT16), .B(n555), .ZN(n556) );
  XOR2_X1 U669 ( .A(KEYINPUT18), .B(KEYINPUT91), .Z(n559) );
  NAND2_X1 U670 ( .A1(G224), .A2(n783), .ZN(n558) );
  XNOR2_X1 U671 ( .A(n559), .B(n558), .ZN(n560) );
  XOR2_X1 U672 ( .A(n560), .B(KEYINPUT17), .Z(n561) );
  NAND2_X1 U673 ( .A1(n732), .A2(n658), .ZN(n566) );
  NAND2_X1 U674 ( .A1(G210), .A2(n568), .ZN(n565) );
  INV_X1 U675 ( .A(KEYINPUT78), .ZN(n567) );
  XNOR2_X2 U676 ( .A(n580), .B(KEYINPUT38), .ZN(n718) );
  NAND2_X1 U677 ( .A1(G214), .A2(n568), .ZN(n717) );
  NAND2_X1 U678 ( .A1(n718), .A2(n717), .ZN(n720) );
  XNOR2_X1 U679 ( .A(KEYINPUT41), .B(n569), .ZN(n689) );
  INV_X1 U680 ( .A(KEYINPUT30), .ZN(n571) );
  AND2_X2 U681 ( .A1(n584), .A2(n718), .ZN(n573) );
  INV_X1 U682 ( .A(KEYINPUT40), .ZN(n574) );
  XNOR2_X1 U683 ( .A(KEYINPUT46), .B(KEYINPUT87), .ZN(n575) );
  XNOR2_X2 U684 ( .A(n385), .B(KEYINPUT1), .ZN(n706) );
  INV_X1 U685 ( .A(n706), .ZN(n621) );
  NAND2_X1 U686 ( .A1(n577), .A2(n717), .ZN(n578) );
  NOR2_X1 U687 ( .A1(n589), .A2(n578), .ZN(n579) );
  NAND2_X1 U688 ( .A1(n416), .A2(n579), .ZN(n604) );
  NOR2_X1 U689 ( .A1(n580), .A2(n604), .ZN(n581) );
  XOR2_X1 U690 ( .A(KEYINPUT36), .B(n581), .Z(n582) );
  NOR2_X1 U691 ( .A1(n621), .A2(n582), .ZN(n685) );
  NOR2_X1 U692 ( .A1(n587), .A2(n583), .ZN(n629) );
  INV_X1 U693 ( .A(n629), .ZN(n586) );
  AND2_X1 U694 ( .A1(n392), .A2(n584), .ZN(n585) );
  NOR2_X1 U695 ( .A1(n588), .A2(n587), .ZN(n682) );
  INV_X1 U696 ( .A(n589), .ZN(n679) );
  NAND2_X1 U697 ( .A1(KEYINPUT47), .A2(n721), .ZN(n590) );
  NOR2_X1 U698 ( .A1(n592), .A2(n616), .ZN(n677) );
  INV_X1 U699 ( .A(n677), .ZN(n593) );
  NAND2_X1 U700 ( .A1(KEYINPUT47), .A2(n593), .ZN(n594) );
  NAND2_X1 U701 ( .A1(n595), .A2(n594), .ZN(n596) );
  NOR2_X1 U702 ( .A1(KEYINPUT47), .A2(n411), .ZN(n597) );
  INV_X1 U703 ( .A(n682), .ZN(n602) );
  NOR2_X1 U704 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U705 ( .A(n603), .B(KEYINPUT107), .ZN(n788) );
  NOR2_X1 U706 ( .A1(n361), .A2(n604), .ZN(n605) );
  XNOR2_X1 U707 ( .A(n605), .B(KEYINPUT43), .ZN(n606) );
  NOR2_X1 U708 ( .A1(n392), .A2(n606), .ZN(n687) );
  INV_X1 U709 ( .A(n687), .ZN(n608) );
  INV_X1 U710 ( .A(n610), .ZN(n611) );
  NOR2_X1 U711 ( .A1(G898), .A2(n783), .ZN(n766) );
  NAND2_X1 U712 ( .A1(n611), .A2(n766), .ZN(n612) );
  XOR2_X1 U713 ( .A(KEYINPUT94), .B(n612), .Z(n613) );
  NOR2_X1 U714 ( .A1(n614), .A2(n613), .ZN(n615) );
  XNOR2_X2 U715 ( .A(n617), .B(KEYINPUT0), .ZN(n645) );
  XNOR2_X1 U716 ( .A(n648), .B(KEYINPUT103), .ZN(n620) );
  INV_X1 U717 ( .A(n700), .ZN(n649) );
  XNOR2_X1 U718 ( .A(KEYINPUT67), .B(KEYINPUT32), .ZN(n626) );
  NOR2_X1 U719 ( .A1(n416), .A2(n621), .ZN(n622) );
  NAND2_X1 U720 ( .A1(n700), .A2(n622), .ZN(n623) );
  XNOR2_X1 U721 ( .A(n623), .B(KEYINPUT77), .ZN(n624) );
  NOR2_X1 U722 ( .A1(n637), .A2(n791), .ZN(n634) );
  INV_X1 U723 ( .A(KEYINPUT86), .ZN(n630) );
  NAND2_X1 U724 ( .A1(n634), .A2(n633), .ZN(n636) );
  INV_X1 U725 ( .A(n637), .ZN(n671) );
  NOR2_X1 U726 ( .A1(n789), .A2(KEYINPUT68), .ZN(n639) );
  INV_X1 U727 ( .A(n791), .ZN(n638) );
  AND2_X1 U728 ( .A1(n639), .A2(n638), .ZN(n640) );
  NAND2_X1 U729 ( .A1(n644), .A2(n383), .ZN(n641) );
  NOR2_X1 U730 ( .A1(n642), .A2(n641), .ZN(n667) );
  NAND2_X1 U731 ( .A1(n713), .A2(n383), .ZN(n646) );
  NOR2_X1 U732 ( .A1(n411), .A2(n647), .ZN(n652) );
  NOR2_X1 U733 ( .A1(n416), .A2(n648), .ZN(n650) );
  NAND2_X1 U734 ( .A1(n650), .A2(n649), .ZN(n664) );
  INV_X1 U735 ( .A(n664), .ZN(n651) );
  NOR2_X1 U736 ( .A1(n652), .A2(n651), .ZN(n653) );
  NAND2_X1 U737 ( .A1(n655), .A2(n654), .ZN(n657) );
  XOR2_X1 U738 ( .A(KEYINPUT45), .B(KEYINPUT64), .Z(n656) );
  NAND2_X1 U739 ( .A1(n741), .A2(G472), .ZN(n661) );
  XNOR2_X1 U740 ( .A(n659), .B(KEYINPUT62), .ZN(n660) );
  XNOR2_X1 U741 ( .A(G101), .B(n664), .ZN(G3) );
  XOR2_X1 U742 ( .A(G104), .B(KEYINPUT109), .Z(n666) );
  NAND2_X1 U743 ( .A1(n667), .A2(n679), .ZN(n665) );
  XNOR2_X1 U744 ( .A(n666), .B(n665), .ZN(G6) );
  XOR2_X1 U745 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n669) );
  NAND2_X1 U746 ( .A1(n667), .A2(n682), .ZN(n668) );
  XNOR2_X1 U747 ( .A(n669), .B(n668), .ZN(n670) );
  XNOR2_X1 U748 ( .A(G107), .B(n670), .ZN(G9) );
  INV_X1 U749 ( .A(n671), .ZN(n672) );
  XOR2_X1 U750 ( .A(G110), .B(n672), .Z(G12) );
  XOR2_X1 U751 ( .A(G128), .B(KEYINPUT29), .Z(n674) );
  NAND2_X1 U752 ( .A1(n677), .A2(n682), .ZN(n673) );
  XNOR2_X1 U753 ( .A(n674), .B(n673), .ZN(G30) );
  XOR2_X1 U754 ( .A(n675), .B(G143), .Z(n676) );
  XNOR2_X1 U755 ( .A(KEYINPUT110), .B(n676), .ZN(G45) );
  NAND2_X1 U756 ( .A1(n677), .A2(n679), .ZN(n678) );
  XNOR2_X1 U757 ( .A(n678), .B(G146), .ZN(G48) );
  XOR2_X1 U758 ( .A(G113), .B(KEYINPUT111), .Z(n681) );
  NAND2_X1 U759 ( .A1(n683), .A2(n679), .ZN(n680) );
  XNOR2_X1 U760 ( .A(n681), .B(n680), .ZN(G15) );
  NAND2_X1 U761 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U762 ( .A(n684), .B(G116), .ZN(G18) );
  XNOR2_X1 U763 ( .A(G125), .B(n685), .ZN(n686) );
  XNOR2_X1 U764 ( .A(n686), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U765 ( .A(G140), .B(n687), .Z(n688) );
  XNOR2_X1 U766 ( .A(KEYINPUT112), .B(n688), .ZN(G42) );
  NOR2_X1 U767 ( .A1(n689), .A2(n396), .ZN(n690) );
  XNOR2_X1 U768 ( .A(n690), .B(KEYINPUT117), .ZN(n698) );
  XNOR2_X1 U769 ( .A(KEYINPUT2), .B(KEYINPUT81), .ZN(n692) );
  NAND2_X1 U770 ( .A1(n759), .A2(n692), .ZN(n691) );
  NAND2_X1 U771 ( .A1(n780), .A2(n692), .ZN(n693) );
  XNOR2_X1 U772 ( .A(n694), .B(KEYINPUT79), .ZN(n696) );
  NAND2_X1 U773 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U774 ( .A1(n698), .A2(n697), .ZN(n731) );
  XOR2_X1 U775 ( .A(KEYINPUT49), .B(KEYINPUT113), .Z(n702) );
  NAND2_X1 U776 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U777 ( .A(n702), .B(n701), .ZN(n703) );
  NOR2_X1 U778 ( .A1(n704), .A2(n703), .ZN(n705) );
  XOR2_X1 U779 ( .A(KEYINPUT114), .B(n705), .Z(n710) );
  NOR2_X1 U780 ( .A1(n707), .A2(n361), .ZN(n708) );
  XNOR2_X1 U781 ( .A(KEYINPUT50), .B(n708), .ZN(n709) );
  NOR2_X1 U782 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U783 ( .A(KEYINPUT115), .B(n711), .Z(n712) );
  NOR2_X1 U784 ( .A1(n713), .A2(n712), .ZN(n714) );
  XOR2_X1 U785 ( .A(KEYINPUT116), .B(n714), .Z(n715) );
  XNOR2_X1 U786 ( .A(n715), .B(KEYINPUT51), .ZN(n716) );
  NOR2_X1 U787 ( .A1(n689), .A2(n716), .ZN(n726) );
  NOR2_X1 U788 ( .A1(n718), .A2(n717), .ZN(n719) );
  NOR2_X1 U789 ( .A1(n411), .A2(n720), .ZN(n722) );
  NOR2_X1 U790 ( .A1(n723), .A2(n722), .ZN(n724) );
  NOR2_X1 U791 ( .A1(n724), .A2(n396), .ZN(n725) );
  NOR2_X1 U792 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U793 ( .A(n727), .B(KEYINPUT52), .ZN(n728) );
  NOR2_X1 U794 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U795 ( .A1(n741), .A2(G210), .ZN(n734) );
  XNOR2_X1 U796 ( .A(n390), .B(n481), .ZN(n733) );
  XNOR2_X1 U797 ( .A(n734), .B(n733), .ZN(n735) );
  NAND2_X1 U798 ( .A1(n750), .A2(G469), .ZN(n739) );
  XOR2_X1 U799 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n736) );
  NOR2_X1 U800 ( .A1(n754), .A2(n740), .ZN(G54) );
  NAND2_X1 U801 ( .A1(n741), .A2(G475), .ZN(n744) );
  XNOR2_X1 U802 ( .A(n744), .B(n743), .ZN(n745) );
  NAND2_X1 U803 ( .A1(n750), .A2(G478), .ZN(n748) );
  NOR2_X1 U804 ( .A1(n754), .A2(n749), .ZN(G63) );
  NAND2_X1 U805 ( .A1(G217), .A2(n750), .ZN(n751) );
  XNOR2_X1 U806 ( .A(n752), .B(n751), .ZN(n753) );
  NOR2_X1 U807 ( .A1(n754), .A2(n753), .ZN(G66) );
  XOR2_X1 U808 ( .A(KEYINPUT121), .B(KEYINPUT61), .Z(n756) );
  NAND2_X1 U809 ( .A1(G224), .A2(G953), .ZN(n755) );
  XNOR2_X1 U810 ( .A(n756), .B(n755), .ZN(n757) );
  NAND2_X1 U811 ( .A1(G898), .A2(n757), .ZN(n758) );
  XOR2_X1 U812 ( .A(KEYINPUT122), .B(n758), .Z(n761) );
  NOR2_X1 U813 ( .A1(G953), .A2(n759), .ZN(n760) );
  NOR2_X1 U814 ( .A1(n761), .A2(n760), .ZN(n768) );
  XOR2_X1 U815 ( .A(n762), .B(G101), .Z(n763) );
  XNOR2_X1 U816 ( .A(n764), .B(n763), .ZN(n765) );
  NOR2_X1 U817 ( .A1(n766), .A2(n765), .ZN(n767) );
  XOR2_X1 U818 ( .A(n768), .B(n767), .Z(G69) );
  XOR2_X1 U819 ( .A(KEYINPUT123), .B(n769), .Z(n772) );
  XNOR2_X1 U820 ( .A(KEYINPUT4), .B(n770), .ZN(n771) );
  XNOR2_X1 U821 ( .A(n772), .B(n771), .ZN(n773) );
  XOR2_X1 U822 ( .A(n393), .B(n773), .Z(n781) );
  INV_X1 U823 ( .A(n781), .ZN(n775) );
  XNOR2_X1 U824 ( .A(G227), .B(n775), .ZN(n776) );
  XNOR2_X1 U825 ( .A(n776), .B(KEYINPUT125), .ZN(n777) );
  NAND2_X1 U826 ( .A1(G900), .A2(n777), .ZN(n778) );
  XNOR2_X1 U827 ( .A(KEYINPUT126), .B(n778), .ZN(n779) );
  NAND2_X1 U828 ( .A1(n779), .A2(G953), .ZN(n786) );
  XNOR2_X1 U829 ( .A(KEYINPUT124), .B(n780), .ZN(n782) );
  XNOR2_X1 U830 ( .A(n782), .B(n781), .ZN(n784) );
  NAND2_X1 U831 ( .A1(n784), .A2(n783), .ZN(n785) );
  NAND2_X1 U832 ( .A1(n786), .A2(n785), .ZN(G72) );
  XOR2_X1 U833 ( .A(G137), .B(n787), .Z(G39) );
  XNOR2_X1 U834 ( .A(G134), .B(n788), .ZN(G36) );
  XNOR2_X1 U835 ( .A(G122), .B(KEYINPUT127), .ZN(n790) );
  XOR2_X1 U836 ( .A(n790), .B(n391), .Z(G24) );
  XOR2_X1 U837 ( .A(n791), .B(G119), .Z(G21) );
  XOR2_X1 U838 ( .A(n792), .B(G131), .Z(G33) );
endmodule

