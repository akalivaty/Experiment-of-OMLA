//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 1 0 1 1 0 0 0 0 0 0 1 0 1 1 0 1 0 0 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 0 0 0 0 0 0 1 1 0 1 1 0 0 1 0 1 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:26 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n727, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n761, new_n762, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n994, new_n995, new_n996,
    new_n997, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  INV_X1    g001(.A(G131), .ZN(new_n188));
  INV_X1    g002(.A(G137), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(KEYINPUT67), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT67), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G137), .ZN(new_n192));
  NAND4_X1  g006(.A1(new_n190), .A2(new_n192), .A3(KEYINPUT11), .A4(G134), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT11), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(KEYINPUT66), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT66), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(KEYINPUT11), .ZN(new_n197));
  INV_X1    g011(.A(G134), .ZN(new_n198));
  AOI22_X1  g012(.A1(new_n195), .A2(new_n197), .B1(new_n198), .B2(G137), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n198), .A2(G137), .ZN(new_n200));
  OAI211_X1 g014(.A(new_n188), .B(new_n193), .C1(new_n199), .C2(new_n200), .ZN(new_n201));
  AOI21_X1  g015(.A(G134), .B1(new_n190), .B2(new_n192), .ZN(new_n202));
  OAI21_X1  g016(.A(KEYINPUT68), .B1(new_n198), .B2(G137), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT68), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n204), .A2(new_n189), .A3(G134), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  OAI21_X1  g020(.A(G131), .B1(new_n202), .B2(new_n206), .ZN(new_n207));
  AND2_X1   g021(.A1(new_n201), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT69), .ZN(new_n209));
  INV_X1    g023(.A(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G143), .ZN(new_n211));
  INV_X1    g025(.A(G143), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G146), .ZN(new_n213));
  AOI21_X1  g027(.A(G128), .B1(new_n211), .B2(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n212), .A2(KEYINPUT1), .A3(G146), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n209), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  XNOR2_X1  g031(.A(G143), .B(G146), .ZN(new_n218));
  OAI211_X1 g032(.A(KEYINPUT69), .B(new_n215), .C1(new_n218), .C2(G128), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT1), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n218), .A2(new_n220), .A3(G128), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n217), .A2(new_n219), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n208), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n211), .A2(new_n213), .ZN(new_n224));
  NAND2_X1  g038(.A1(KEYINPUT0), .A2(G128), .ZN(new_n225));
  NOR3_X1   g039(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n226));
  OAI21_X1  g040(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  OAI211_X1 g042(.A(new_n224), .B(new_n225), .C1(new_n226), .C2(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n218), .A2(KEYINPUT0), .A3(G128), .ZN(new_n230));
  AND2_X1   g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n201), .ZN(new_n232));
  INV_X1    g046(.A(new_n200), .ZN(new_n233));
  XNOR2_X1  g047(.A(KEYINPUT66), .B(KEYINPUT11), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n189), .A2(G134), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n233), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n188), .B1(new_n236), .B2(new_n193), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n231), .B1(new_n232), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(G119), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(KEYINPUT71), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT71), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G119), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n240), .A2(new_n242), .A3(G116), .ZN(new_n243));
  INV_X1    g057(.A(G116), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G119), .ZN(new_n245));
  INV_X1    g059(.A(G113), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(KEYINPUT2), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT2), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G113), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  AND3_X1   g064(.A1(new_n243), .A2(new_n245), .A3(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n250), .B1(new_n243), .B2(new_n245), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n223), .A2(new_n238), .A3(new_n253), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n254), .B(KEYINPUT28), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n223), .A2(new_n238), .ZN(new_n256));
  INV_X1    g070(.A(new_n253), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n255), .A2(new_n258), .ZN(new_n259));
  NOR2_X1   g073(.A1(G237), .A2(G953), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G210), .ZN(new_n261));
  XOR2_X1   g075(.A(new_n261), .B(KEYINPUT27), .Z(new_n262));
  XNOR2_X1  g076(.A(KEYINPUT26), .B(G101), .ZN(new_n263));
  XOR2_X1   g077(.A(new_n262), .B(new_n263), .Z(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(KEYINPUT29), .ZN(new_n265));
  INV_X1    g079(.A(new_n254), .ZN(new_n266));
  AND3_X1   g080(.A1(new_n223), .A2(new_n238), .A3(KEYINPUT30), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT65), .ZN(new_n268));
  AND3_X1   g082(.A1(new_n229), .A2(new_n268), .A3(new_n230), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n268), .B1(new_n229), .B2(new_n230), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n193), .B1(new_n199), .B2(new_n200), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(G131), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(new_n201), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n271), .A2(new_n274), .ZN(new_n275));
  AND3_X1   g089(.A1(new_n217), .A2(new_n219), .A3(new_n221), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n201), .A2(new_n207), .ZN(new_n277));
  NOR3_X1   g091(.A1(new_n276), .A2(new_n277), .A3(KEYINPUT70), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT70), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n279), .B1(new_n208), .B2(new_n222), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n275), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT30), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n267), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n266), .B1(new_n283), .B2(new_n257), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n284), .A2(new_n264), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n281), .A2(new_n257), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n255), .A2(new_n286), .A3(new_n264), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT29), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  OAI221_X1 g103(.A(new_n187), .B1(new_n259), .B2(new_n265), .C1(new_n285), .C2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(G472), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n264), .B1(new_n255), .B2(new_n286), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n284), .A2(KEYINPUT72), .A3(KEYINPUT31), .A4(new_n264), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n223), .A2(new_n238), .A3(KEYINPUT30), .ZN(new_n294));
  OAI21_X1  g108(.A(KEYINPUT70), .B1(new_n276), .B2(new_n277), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n208), .A2(new_n279), .A3(new_n222), .ZN(new_n296));
  AOI22_X1  g110(.A1(new_n295), .A2(new_n296), .B1(new_n274), .B2(new_n271), .ZN(new_n297));
  OAI211_X1 g111(.A(new_n257), .B(new_n294), .C1(new_n297), .C2(KEYINPUT30), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n298), .A2(KEYINPUT72), .A3(new_n254), .A4(new_n264), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT31), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n292), .B1(new_n293), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT73), .ZN(new_n303));
  OR3_X1    g117(.A1(new_n303), .A2(G472), .A3(G902), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n303), .B1(G472), .B2(G902), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  NOR3_X1   g121(.A1(new_n302), .A2(KEYINPUT32), .A3(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT32), .ZN(new_n309));
  INV_X1    g123(.A(new_n292), .ZN(new_n310));
  AND2_X1   g124(.A1(new_n299), .A2(new_n300), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n299), .A2(new_n300), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n310), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n309), .B1(new_n313), .B2(new_n306), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n291), .B1(new_n308), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT78), .ZN(new_n316));
  INV_X1    g130(.A(G128), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n239), .A2(new_n317), .ZN(new_n318));
  XNOR2_X1  g132(.A(KEYINPUT71), .B(G119), .ZN(new_n319));
  OAI211_X1 g133(.A(KEYINPUT23), .B(new_n318), .C1(new_n319), .C2(new_n317), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT23), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n321), .B1(new_n319), .B2(G128), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  XOR2_X1   g137(.A(KEYINPUT24), .B(G110), .Z(new_n324));
  OAI21_X1  g138(.A(new_n318), .B1(new_n319), .B2(new_n317), .ZN(new_n325));
  OAI22_X1  g139(.A1(new_n323), .A2(G110), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(G140), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G125), .ZN(new_n328));
  INV_X1    g142(.A(G125), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G140), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT74), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n328), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n329), .A2(KEYINPUT74), .A3(G140), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n332), .A2(KEYINPUT16), .A3(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT16), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n328), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n210), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  AND3_X1   g151(.A1(new_n328), .A2(new_n330), .A3(new_n210), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n326), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n189), .A2(KEYINPUT22), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT22), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(G137), .ZN(new_n343));
  AND3_X1   g157(.A1(new_n341), .A2(new_n343), .A3(KEYINPUT75), .ZN(new_n344));
  AOI21_X1  g158(.A(KEYINPUT75), .B1(new_n341), .B2(new_n343), .ZN(new_n345));
  OAI21_X1  g159(.A(KEYINPUT76), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT75), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n342), .A2(G137), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n189), .A2(KEYINPUT22), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n347), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT76), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n341), .A2(new_n343), .A3(KEYINPUT75), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n350), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(G953), .ZN(new_n354));
  AND3_X1   g168(.A1(new_n354), .A2(G221), .A3(G234), .ZN(new_n355));
  AND3_X1   g169(.A1(new_n346), .A2(new_n353), .A3(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n355), .B1(new_n346), .B2(new_n353), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n323), .A2(G110), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n325), .A2(new_n324), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n334), .A2(new_n210), .A3(new_n336), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  OAI211_X1 g176(.A(new_n359), .B(new_n360), .C1(new_n362), .C2(new_n337), .ZN(new_n363));
  AND3_X1   g177(.A1(new_n340), .A2(new_n358), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n358), .B1(new_n363), .B2(new_n340), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n187), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NOR2_X1   g180(.A1(KEYINPUT77), .A2(KEYINPUT25), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  OAI221_X1 g182(.A(new_n187), .B1(KEYINPUT77), .B2(KEYINPUT25), .C1(new_n364), .C2(new_n365), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(G217), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n371), .B1(G234), .B2(new_n187), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n316), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(new_n372), .ZN(new_n374));
  AOI211_X1 g188(.A(KEYINPUT78), .B(new_n374), .C1(new_n368), .C2(new_n369), .ZN(new_n375));
  OR2_X1    g189(.A1(new_n364), .A2(new_n365), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n372), .A2(G902), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  NOR3_X1   g193(.A1(new_n373), .A2(new_n375), .A3(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT97), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n354), .A2(G227), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n382), .B(KEYINPUT79), .ZN(new_n383));
  XNOR2_X1  g197(.A(G110), .B(G140), .ZN(new_n384));
  XOR2_X1   g198(.A(new_n383), .B(new_n384), .Z(new_n385));
  INV_X1    g199(.A(G104), .ZN(new_n386));
  OAI21_X1  g200(.A(KEYINPUT3), .B1(new_n386), .B2(G107), .ZN(new_n387));
  AOI21_X1  g201(.A(G101), .B1(new_n386), .B2(G107), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT3), .ZN(new_n389));
  INV_X1    g203(.A(G107), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n389), .A2(new_n390), .A3(G104), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n387), .A2(new_n388), .A3(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(G101), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n390), .A2(G104), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n386), .A2(G107), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n393), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n215), .B1(new_n218), .B2(G128), .ZN(new_n398));
  AND4_X1   g212(.A1(new_n220), .A2(new_n211), .A3(new_n213), .A4(G128), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n392), .B(new_n397), .C1(new_n398), .C2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n217), .A2(new_n219), .ZN(new_n401));
  AND3_X1   g215(.A1(new_n387), .A2(new_n388), .A3(new_n391), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n221), .B1(new_n402), .B2(new_n396), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n400), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n404), .A2(KEYINPUT12), .A3(new_n274), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(KEYINPUT81), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT81), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n404), .A2(new_n407), .A3(KEYINPUT12), .A4(new_n274), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n404), .A2(new_n274), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT12), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n406), .A2(new_n408), .A3(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n274), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n402), .A2(new_n396), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n222), .A2(KEYINPUT10), .A3(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n387), .A2(new_n391), .A3(new_n395), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(G101), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n417), .A2(KEYINPUT4), .A3(new_n392), .ZN(new_n418));
  XOR2_X1   g232(.A(KEYINPUT80), .B(KEYINPUT4), .Z(new_n419));
  NAND3_X1  g233(.A1(new_n416), .A2(G101), .A3(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n231), .A2(new_n418), .A3(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT10), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n400), .A2(new_n422), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n413), .A2(new_n415), .A3(new_n421), .A4(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n385), .B1(new_n412), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n385), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n415), .A2(new_n421), .A3(new_n423), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n426), .B1(new_n274), .B2(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(KEYINPUT82), .B1(new_n425), .B2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT82), .ZN(new_n430));
  AND2_X1   g244(.A1(new_n424), .A2(new_n385), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n427), .A2(new_n274), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(new_n424), .ZN(new_n434));
  AOI21_X1  g248(.A(KEYINPUT12), .B1(new_n404), .B2(new_n274), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n435), .B1(KEYINPUT81), .B2(new_n405), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n434), .B1(new_n436), .B2(new_n408), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n430), .B(new_n433), .C1(new_n437), .C2(new_n385), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n429), .A2(new_n438), .A3(G469), .ZN(new_n439));
  INV_X1    g253(.A(G469), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n440), .A2(new_n187), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n412), .A2(new_n431), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n432), .A2(new_n424), .ZN(new_n443));
  INV_X1    g257(.A(new_n385), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(G902), .B1(new_n442), .B2(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n441), .B1(new_n446), .B2(new_n440), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n439), .A2(new_n447), .ZN(new_n448));
  XNOR2_X1  g262(.A(KEYINPUT9), .B(G234), .ZN(new_n449));
  OAI21_X1  g263(.A(G221), .B1(new_n449), .B2(G902), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(G214), .B1(G237), .B2(G902), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  OAI21_X1  g267(.A(G210), .B1(G237), .B2(G902), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n243), .A2(KEYINPUT5), .A3(new_n245), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT5), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n319), .A2(new_n457), .A3(G116), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n456), .A2(G113), .A3(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n243), .A2(new_n245), .A3(new_n250), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n459), .A2(new_n460), .A3(new_n414), .ZN(new_n461));
  AND2_X1   g275(.A1(new_n416), .A2(G101), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n392), .A2(KEYINPUT4), .ZN(new_n463));
  OAI22_X1  g277(.A1(new_n462), .A2(new_n463), .B1(new_n251), .B2(new_n252), .ZN(new_n464));
  INV_X1    g278(.A(new_n420), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n461), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  XNOR2_X1  g280(.A(G110), .B(G122), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n467), .B(new_n461), .C1(new_n464), .C2(new_n465), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n469), .A2(KEYINPUT6), .A3(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT6), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n466), .A2(new_n472), .A3(new_n468), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n229), .A2(new_n230), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(G125), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n217), .A2(new_n329), .A3(new_n219), .A4(new_n221), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(G224), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n478), .A2(G953), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n477), .B(new_n479), .ZN(new_n480));
  AND3_X1   g294(.A1(new_n471), .A2(new_n473), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n459), .A2(new_n460), .ZN(new_n482));
  INV_X1    g296(.A(new_n414), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(new_n461), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n467), .B(KEYINPUT8), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT7), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n477), .B1(new_n488), .B2(new_n479), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n479), .A2(new_n488), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n475), .A2(new_n476), .A3(new_n490), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n487), .A2(new_n489), .A3(new_n470), .A4(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(new_n187), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n455), .B1(new_n481), .B2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(new_n466), .ZN(new_n495));
  AOI22_X1  g309(.A1(new_n495), .A2(new_n467), .B1(new_n485), .B2(new_n486), .ZN(new_n496));
  AND2_X1   g310(.A1(new_n489), .A2(new_n491), .ZN(new_n497));
  AOI21_X1  g311(.A(G902), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n471), .A2(new_n473), .A3(new_n480), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n498), .A2(new_n454), .A3(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n453), .B1(new_n494), .B2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT95), .ZN(new_n502));
  NOR3_X1   g316(.A1(new_n449), .A2(new_n371), .A3(G953), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(G122), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(G116), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n244), .A2(G122), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n506), .A2(new_n507), .A3(new_n390), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT93), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n506), .A2(new_n507), .A3(KEYINPUT93), .A4(new_n390), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n506), .B1(new_n507), .B2(KEYINPUT14), .ZN(new_n512));
  OAI21_X1  g326(.A(KEYINPUT14), .B1(new_n505), .B2(G116), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT94), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n507), .A2(KEYINPUT94), .A3(KEYINPUT14), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n512), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n510), .B(new_n511), .C1(new_n517), .C2(new_n390), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT92), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n212), .A2(G128), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n317), .A2(G143), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n520), .A2(new_n521), .A3(KEYINPUT91), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(KEYINPUT91), .B1(new_n520), .B2(new_n521), .ZN(new_n524));
  NOR3_X1   g338(.A1(new_n523), .A2(new_n524), .A3(new_n198), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n520), .A2(new_n521), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT91), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(G134), .B1(new_n528), .B2(new_n522), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n519), .B1(new_n525), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n198), .B1(new_n523), .B2(new_n524), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n528), .A2(G134), .A3(new_n522), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n531), .A2(new_n532), .A3(KEYINPUT92), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n518), .B1(new_n530), .B2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n508), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n390), .B1(new_n506), .B2(new_n507), .ZN(new_n536));
  OR2_X1    g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n520), .A2(new_n521), .A3(KEYINPUT13), .ZN(new_n538));
  OAI211_X1 g352(.A(new_n538), .B(G134), .C1(KEYINPUT13), .C2(new_n520), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n537), .A2(new_n531), .A3(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n504), .B1(new_n534), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n510), .A2(new_n511), .ZN(new_n543));
  INV_X1    g357(.A(new_n517), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n543), .B1(new_n544), .B2(G107), .ZN(new_n545));
  AND3_X1   g359(.A1(new_n531), .A2(new_n532), .A3(KEYINPUT92), .ZN(new_n546));
  AOI21_X1  g360(.A(KEYINPUT92), .B1(new_n531), .B2(new_n532), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n548), .A2(new_n540), .A3(new_n503), .ZN(new_n549));
  AOI21_X1  g363(.A(G902), .B1(new_n542), .B2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(G478), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n551), .A2(KEYINPUT15), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  AOI211_X1 g368(.A(G902), .B(new_n552), .C1(new_n542), .C2(new_n549), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n502), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NOR3_X1   g370(.A1(new_n534), .A2(new_n541), .A3(new_n504), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n503), .B1(new_n548), .B2(new_n540), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n187), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(new_n552), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n550), .A2(new_n553), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n560), .A2(new_n561), .A3(KEYINPUT95), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n556), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(G952), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n564), .A2(G953), .ZN(new_n565));
  INV_X1    g379(.A(G234), .ZN(new_n566));
  INV_X1    g380(.A(G237), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n565), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  XOR2_X1   g383(.A(KEYINPUT21), .B(G898), .Z(new_n570));
  XNOR2_X1  g384(.A(new_n570), .B(KEYINPUT96), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  AOI211_X1 g386(.A(new_n187), .B(new_n354), .C1(G234), .C2(G237), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n569), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  XOR2_X1   g389(.A(KEYINPUT89), .B(G475), .Z(new_n576));
  XNOR2_X1  g390(.A(G113), .B(G122), .ZN(new_n577));
  XNOR2_X1  g391(.A(KEYINPUT86), .B(G104), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n577), .B(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT87), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n579), .B(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n567), .A2(new_n354), .A3(G214), .ZN(new_n582));
  NOR2_X1   g396(.A1(KEYINPUT84), .A2(G143), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI211_X1 g398(.A(new_n260), .B(G214), .C1(KEYINPUT84), .C2(G143), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(G131), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT17), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n584), .A2(new_n585), .A3(new_n188), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n334), .A2(new_n336), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(G146), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n188), .B1(new_n584), .B2(new_n585), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(KEYINPUT17), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n590), .A2(new_n592), .A3(new_n361), .A4(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n586), .A2(KEYINPUT18), .A3(G131), .ZN(new_n596));
  NAND2_X1  g410(.A1(KEYINPUT18), .A2(G131), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n584), .A2(new_n585), .A3(new_n597), .ZN(new_n598));
  AND3_X1   g412(.A1(new_n332), .A2(G146), .A3(new_n333), .ZN(new_n599));
  OAI211_X1 g413(.A(new_n596), .B(new_n598), .C1(new_n599), .C2(new_n338), .ZN(new_n600));
  AND3_X1   g414(.A1(new_n581), .A2(new_n595), .A3(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n579), .B1(new_n595), .B2(new_n600), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n187), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n576), .B1(new_n603), .B2(KEYINPUT90), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT90), .ZN(new_n605));
  OAI211_X1 g419(.A(new_n605), .B(new_n187), .C1(new_n601), .C2(new_n602), .ZN(new_n606));
  XOR2_X1   g420(.A(KEYINPUT83), .B(KEYINPUT20), .Z(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT85), .ZN(new_n609));
  INV_X1    g423(.A(new_n589), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n609), .B1(new_n610), .B2(new_n593), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n587), .A2(KEYINPUT85), .A3(new_n589), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT19), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n613), .B1(new_n332), .B2(new_n333), .ZN(new_n614));
  AOI21_X1  g428(.A(KEYINPUT19), .B1(new_n328), .B2(new_n330), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n210), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n611), .A2(new_n612), .A3(new_n592), .A4(new_n616), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n579), .B1(new_n617), .B2(new_n600), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n601), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(G475), .A2(G902), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n608), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  OR2_X1    g436(.A1(new_n621), .A2(KEYINPUT88), .ZN(new_n623));
  AOI21_X1  g437(.A(KEYINPUT20), .B1(new_n621), .B2(KEYINPUT88), .ZN(new_n624));
  OAI211_X1 g438(.A(new_n623), .B(new_n624), .C1(new_n601), .C2(new_n618), .ZN(new_n625));
  AOI22_X1  g439(.A1(new_n604), .A2(new_n606), .B1(new_n622), .B2(new_n625), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n501), .A2(new_n563), .A3(new_n575), .A4(new_n626), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n381), .B1(new_n451), .B2(new_n627), .ZN(new_n628));
  NOR3_X1   g442(.A1(new_n554), .A2(new_n555), .A3(new_n502), .ZN(new_n629));
  AOI21_X1  g443(.A(KEYINPUT95), .B1(new_n560), .B2(new_n561), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n626), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NOR3_X1   g445(.A1(new_n481), .A2(new_n493), .A3(new_n455), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n454), .B1(new_n498), .B2(new_n499), .ZN(new_n633));
  OAI211_X1 g447(.A(new_n575), .B(new_n452), .C1(new_n632), .C2(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n450), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n636), .B1(new_n439), .B2(new_n447), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n635), .A2(KEYINPUT97), .A3(new_n637), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n315), .A2(new_n380), .A3(new_n628), .A4(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(G101), .ZN(G3));
  OAI21_X1  g454(.A(G472), .B1(new_n302), .B2(G902), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n313), .A2(new_n306), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n641), .A2(new_n642), .A3(new_n637), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  OAI21_X1  g458(.A(KEYINPUT33), .B1(new_n557), .B2(new_n558), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT33), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n542), .A2(new_n549), .A3(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n645), .A2(G478), .A3(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n551), .A2(new_n187), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n649), .B1(new_n550), .B2(new_n551), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n626), .A2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n373), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n370), .A2(new_n316), .A3(new_n372), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n653), .A2(new_n654), .A3(new_n378), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n655), .A2(new_n634), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n644), .A2(new_n652), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(KEYINPUT98), .ZN(new_n658));
  XNOR2_X1  g472(.A(KEYINPUT34), .B(G104), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G6));
  NAND2_X1  g474(.A1(new_n617), .A2(new_n600), .ZN(new_n661));
  INV_X1    g475(.A(new_n579), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n581), .A2(new_n595), .A3(new_n600), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n621), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(new_n608), .ZN(new_n666));
  OR2_X1    g480(.A1(new_n666), .A2(KEYINPUT99), .ZN(new_n667));
  AOI22_X1  g481(.A1(new_n666), .A2(KEYINPUT99), .B1(new_n606), .B2(new_n604), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n629), .A2(new_n630), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  NOR3_X1   g484(.A1(new_n670), .A2(new_n655), .A3(new_n634), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n644), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT35), .B(G107), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G9));
  NOR2_X1   g488(.A1(new_n358), .A2(KEYINPUT36), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n340), .A2(new_n363), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n377), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT100), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n653), .A2(new_n680), .A3(new_n654), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n641), .A2(new_n642), .A3(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT101), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n641), .A2(new_n642), .A3(new_n681), .A4(KEYINPUT101), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n684), .A2(new_n628), .A3(new_n638), .A4(new_n685), .ZN(new_n686));
  XOR2_X1   g500(.A(KEYINPUT37), .B(G110), .Z(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G12));
  NAND2_X1  g502(.A1(new_n681), .A2(new_n501), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n573), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n568), .B1(new_n691), .B2(G900), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n667), .A2(new_n668), .A3(new_n669), .A4(new_n692), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n693), .A2(new_n451), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n315), .A2(new_n690), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G128), .ZN(G30));
  NOR2_X1   g510(.A1(new_n632), .A2(new_n633), .ZN(new_n697));
  XNOR2_X1  g511(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n698));
  OR2_X1    g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n697), .A2(new_n698), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n625), .B1(new_n665), .B2(new_n607), .ZN(new_n702));
  INV_X1    g516(.A(new_n576), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n595), .A2(new_n600), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n662), .ZN(new_n705));
  AOI21_X1  g519(.A(G902), .B1(new_n705), .B2(new_n664), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n703), .B1(new_n706), .B2(new_n605), .ZN(new_n707));
  INV_X1    g521(.A(new_n606), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n702), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n669), .A2(new_n709), .ZN(new_n710));
  NOR4_X1   g524(.A1(new_n701), .A2(new_n453), .A3(new_n681), .A4(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n692), .B(KEYINPUT39), .ZN(new_n712));
  AND2_X1   g526(.A1(new_n637), .A2(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT40), .ZN(new_n714));
  OR2_X1    g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(new_n264), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n284), .A2(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(new_n258), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n716), .A2(new_n254), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n187), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  OAI21_X1  g534(.A(G472), .B1(new_n717), .B2(new_n720), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n721), .B1(new_n308), .B2(new_n314), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n713), .A2(new_n714), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n711), .A2(new_n715), .A3(new_n722), .A4(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G143), .ZN(G45));
  AND2_X1   g539(.A1(new_n648), .A2(new_n650), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n726), .A2(new_n709), .A3(new_n692), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n451), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n315), .A2(new_n690), .A3(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G146), .ZN(G48));
  AOI22_X1  g544(.A1(new_n412), .A2(new_n431), .B1(new_n443), .B2(new_n444), .ZN(new_n731));
  OAI21_X1  g545(.A(G469), .B1(new_n731), .B2(G902), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n426), .B1(new_n436), .B2(new_n408), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n385), .B1(new_n432), .B2(new_n424), .ZN(new_n734));
  OAI211_X1 g548(.A(new_n440), .B(new_n187), .C1(new_n733), .C2(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n732), .A2(new_n450), .A3(new_n735), .ZN(new_n736));
  NOR4_X1   g550(.A1(new_n634), .A2(new_n736), .A3(new_n626), .A4(new_n651), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n315), .A2(new_n380), .A3(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(KEYINPUT41), .B(G113), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(KEYINPUT103), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n738), .B(new_n740), .ZN(G15));
  OAI21_X1  g555(.A(KEYINPUT32), .B1(new_n302), .B2(new_n307), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n313), .A2(new_n309), .A3(new_n306), .ZN(new_n743));
  AOI22_X1  g557(.A1(new_n742), .A2(new_n743), .B1(G472), .B2(new_n290), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n744), .A2(new_n736), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(new_n671), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G116), .ZN(G18));
  AND2_X1   g561(.A1(new_n635), .A2(new_n681), .ZN(new_n748));
  AND2_X1   g562(.A1(new_n745), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(new_n239), .ZN(G21));
  NAND2_X1  g564(.A1(new_n259), .A2(new_n716), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n751), .B1(new_n311), .B2(new_n312), .ZN(new_n752));
  XOR2_X1   g566(.A(new_n306), .B(KEYINPUT104), .Z(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  AND2_X1   g568(.A1(new_n641), .A2(new_n754), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n452), .B1(new_n632), .B2(new_n633), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n710), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n736), .A2(new_n574), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n755), .A2(new_n380), .A3(new_n757), .A4(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G122), .ZN(G24));
  NOR3_X1   g574(.A1(new_n727), .A2(new_n756), .A3(new_n736), .ZN(new_n761));
  AND4_X1   g575(.A1(new_n641), .A2(new_n761), .A3(new_n681), .A4(new_n754), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(new_n329), .ZN(G27));
  NAND2_X1  g577(.A1(new_n742), .A2(new_n743), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n655), .B1(new_n764), .B2(new_n291), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(KEYINPUT105), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT105), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n767), .B1(new_n744), .B2(new_n655), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n425), .A2(new_n428), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(G469), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n447), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n636), .A2(new_n453), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n771), .A2(new_n697), .A3(new_n772), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n773), .A2(new_n727), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n766), .A2(new_n768), .A3(KEYINPUT42), .A4(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(new_n727), .ZN(new_n776));
  INV_X1    g590(.A(new_n773), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n765), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT42), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n775), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G131), .ZN(G33));
  NOR4_X1   g596(.A1(new_n744), .A2(new_n655), .A3(new_n693), .A4(new_n773), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(new_n198), .ZN(G36));
  NAND2_X1  g598(.A1(new_n697), .A2(new_n452), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n626), .A2(new_n726), .ZN(new_n786));
  XNOR2_X1  g600(.A(KEYINPUT107), .B(KEYINPUT43), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT43), .ZN(new_n789));
  OAI22_X1  g603(.A1(new_n788), .A2(KEYINPUT108), .B1(new_n789), .B2(new_n786), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n788), .A2(KEYINPUT108), .ZN(new_n791));
  OR2_X1    g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n641), .A2(new_n642), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n792), .A2(new_n793), .A3(new_n681), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT44), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n785), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n792), .A2(KEYINPUT44), .A3(new_n793), .A4(new_n681), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n429), .A2(new_n438), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT45), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n440), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(KEYINPUT106), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT106), .ZN(new_n803));
  AOI21_X1  g617(.A(KEYINPUT45), .B1(new_n429), .B2(new_n438), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n803), .B1(new_n804), .B2(new_n440), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n769), .A2(KEYINPUT45), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n802), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n441), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT46), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n441), .A2(new_n810), .ZN(new_n812));
  AOI22_X1  g626(.A1(new_n807), .A2(new_n812), .B1(new_n440), .B2(new_n446), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n636), .B1(new_n811), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(new_n712), .ZN(new_n815));
  INV_X1    g629(.A(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n798), .A2(new_n816), .ZN(new_n817));
  XOR2_X1   g631(.A(KEYINPUT109), .B(G137), .Z(new_n818));
  XNOR2_X1  g632(.A(new_n817), .B(new_n818), .ZN(G39));
  NAND2_X1  g633(.A1(new_n807), .A2(new_n812), .ZN(new_n820));
  AOI22_X1  g634(.A1(new_n801), .A2(KEYINPUT106), .B1(KEYINPUT45), .B2(new_n769), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n441), .B1(new_n821), .B2(new_n805), .ZN(new_n822));
  OAI211_X1 g636(.A(new_n820), .B(new_n735), .C1(new_n822), .C2(KEYINPUT46), .ZN(new_n823));
  NAND2_X1  g637(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n823), .A2(new_n450), .A3(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n824), .ZN(new_n826));
  NOR2_X1   g640(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n825), .B1(new_n814), .B2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(new_n785), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n744), .A2(new_n655), .A3(new_n776), .A4(new_n830), .ZN(new_n831));
  OR2_X1    g645(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n832), .B(G140), .ZN(G42));
  INV_X1    g647(.A(KEYINPUT50), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n792), .A2(new_n380), .A3(new_n569), .A4(new_n755), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n452), .B1(new_n699), .B2(new_n700), .ZN(new_n836));
  INV_X1    g650(.A(new_n736), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(KEYINPUT117), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT117), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n836), .A2(new_n840), .A3(new_n837), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n834), .B1(new_n835), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n569), .B1(new_n790), .B2(new_n791), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n755), .A2(new_n380), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n846), .A2(KEYINPUT50), .A3(new_n841), .A4(new_n839), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n843), .A2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(new_n722), .ZN(new_n849));
  NOR4_X1   g663(.A1(new_n655), .A2(new_n785), .A3(new_n568), .A4(new_n736), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n726), .A2(new_n709), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n785), .A2(new_n736), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n569), .B(new_n853), .C1(new_n790), .C2(new_n791), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n755), .A2(new_n681), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n852), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n848), .A2(new_n857), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n732), .A2(new_n735), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(new_n636), .ZN(new_n860));
  AOI211_X1 g674(.A(new_n636), .B(new_n826), .C1(new_n811), .C2(new_n813), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n828), .B1(new_n823), .B2(new_n450), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n860), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n835), .A2(new_n785), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n858), .B1(new_n865), .B2(KEYINPUT116), .ZN(new_n866));
  INV_X1    g680(.A(new_n864), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n867), .B1(new_n829), .B2(new_n860), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT116), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(KEYINPUT51), .B1(new_n866), .B2(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n846), .A2(new_n501), .A3(new_n837), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n849), .A2(new_n652), .A3(new_n850), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n872), .A2(new_n565), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n766), .A2(new_n768), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT48), .ZN(new_n876));
  OR3_X1    g690(.A1(new_n875), .A2(new_n876), .A3(new_n854), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n876), .B1(new_n875), .B2(new_n854), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n874), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n857), .A2(KEYINPUT118), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT118), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n882), .B1(new_n852), .B2(new_n856), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n848), .A2(new_n881), .A3(KEYINPUT51), .A4(new_n883), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n880), .B1(new_n884), .B2(new_n868), .ZN(new_n885));
  OAI21_X1  g699(.A(KEYINPUT119), .B1(new_n871), .B2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT51), .ZN(new_n887));
  OAI211_X1 g701(.A(new_n848), .B(new_n857), .C1(new_n868), .C2(new_n869), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n865), .A2(KEYINPUT116), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n887), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT119), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n884), .A2(new_n868), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n892), .A2(new_n879), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n890), .A2(new_n891), .A3(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT113), .ZN(new_n895));
  INV_X1    g709(.A(new_n634), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT112), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n897), .B1(new_n626), .B2(new_n651), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n726), .A2(new_n709), .A3(KEYINPUT112), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n380), .A2(new_n896), .A3(new_n898), .A4(new_n899), .ZN(new_n900));
  OR2_X1    g714(.A1(new_n643), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n895), .B1(new_n639), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n709), .B1(new_n560), .B2(new_n561), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n644), .A2(new_n656), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n686), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n639), .A2(new_n895), .A3(new_n901), .ZN(new_n907));
  AOI21_X1  g721(.A(KEYINPUT114), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n639), .A2(new_n901), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(KEYINPUT113), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n686), .A2(new_n904), .ZN(new_n911));
  AND4_X1   g725(.A1(KEYINPUT114), .A2(new_n910), .A3(new_n911), .A4(new_n907), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n908), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n755), .A2(new_n681), .A3(new_n761), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n771), .A2(new_n669), .A3(new_n501), .A4(new_n709), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n692), .A2(new_n450), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n915), .A2(new_n681), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n722), .A2(new_n917), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n695), .A2(new_n729), .A3(new_n914), .A4(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT52), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n689), .B1(new_n764), .B2(new_n291), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n762), .B1(new_n922), .B2(new_n694), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n923), .A2(KEYINPUT52), .A3(new_n729), .A4(new_n918), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n921), .A2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(new_n670), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n765), .A2(new_n926), .A3(new_n692), .A4(new_n777), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n667), .A2(new_n668), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n560), .A2(new_n561), .A3(new_n692), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n930), .A2(new_n637), .A3(new_n681), .A4(new_n830), .ZN(new_n931));
  OR2_X1    g745(.A1(new_n931), .A2(new_n744), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT115), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n774), .A2(new_n641), .A3(new_n681), .A4(new_n754), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n927), .A2(new_n932), .A3(new_n933), .A4(new_n934), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n934), .B1(new_n931), .B2(new_n744), .ZN(new_n936));
  OAI21_X1  g750(.A(KEYINPUT115), .B1(new_n783), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  OAI211_X1 g752(.A(new_n315), .B(new_n837), .C1(new_n671), .C2(new_n748), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n939), .A2(new_n738), .A3(new_n759), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n940), .B1(new_n775), .B2(new_n780), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n925), .A2(new_n938), .A3(new_n941), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n923), .A2(new_n920), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n943), .A2(KEYINPUT53), .ZN(new_n944));
  NOR3_X1   g758(.A1(new_n913), .A2(new_n942), .A3(new_n944), .ZN(new_n945));
  AND3_X1   g759(.A1(new_n925), .A2(new_n938), .A3(new_n941), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT114), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n643), .A2(new_n900), .ZN(new_n948));
  NOR3_X1   g762(.A1(new_n451), .A2(new_n627), .A3(new_n381), .ZN(new_n949));
  AOI21_X1  g763(.A(KEYINPUT97), .B1(new_n635), .B2(new_n637), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n948), .B1(new_n951), .B2(new_n765), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n686), .B(new_n904), .C1(new_n952), .C2(new_n895), .ZN(new_n953));
  INV_X1    g767(.A(new_n907), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n947), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n906), .A2(KEYINPUT114), .A3(new_n907), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(KEYINPUT53), .B1(new_n946), .B2(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(KEYINPUT54), .B1(new_n945), .B2(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT53), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n960), .B1(new_n913), .B2(new_n942), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT54), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n943), .A2(new_n960), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n946), .A2(new_n957), .A3(new_n963), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n961), .A2(new_n962), .A3(new_n964), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n886), .A2(new_n894), .A3(new_n959), .A4(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n564), .A2(new_n354), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n859), .B(KEYINPUT49), .ZN(new_n969));
  NOR4_X1   g783(.A1(new_n655), .A2(new_n453), .A3(new_n636), .A4(new_n786), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n849), .A2(new_n701), .A3(new_n969), .A4(new_n970), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n971), .B(KEYINPUT111), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n968), .A2(new_n972), .ZN(G75));
  AND3_X1   g787(.A1(new_n946), .A2(new_n957), .A3(new_n963), .ZN(new_n974));
  OAI211_X1 g788(.A(G210), .B(G902), .C1(new_n974), .C2(new_n958), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n471), .A2(new_n473), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n976), .B(new_n480), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n977), .B(KEYINPUT55), .ZN(new_n978));
  XOR2_X1   g792(.A(KEYINPUT120), .B(KEYINPUT56), .Z(new_n979));
  AND3_X1   g793(.A1(new_n975), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT56), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n978), .B1(new_n975), .B2(new_n981), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n354), .A2(G952), .ZN(new_n983));
  NOR3_X1   g797(.A1(new_n980), .A2(new_n982), .A3(new_n983), .ZN(G51));
  XNOR2_X1  g798(.A(new_n441), .B(KEYINPUT57), .ZN(new_n985));
  NOR3_X1   g799(.A1(new_n974), .A2(new_n958), .A3(KEYINPUT54), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n962), .B1(new_n961), .B2(new_n964), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n985), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(new_n731), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n961), .A2(new_n964), .ZN(new_n991));
  NAND4_X1  g805(.A1(new_n991), .A2(G902), .A3(new_n805), .A4(new_n821), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n983), .B1(new_n990), .B2(new_n992), .ZN(G54));
  AND2_X1   g807(.A1(KEYINPUT58), .A2(G475), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n991), .A2(G902), .A3(new_n994), .ZN(new_n995));
  AND2_X1   g809(.A1(new_n995), .A2(new_n619), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n995), .A2(new_n619), .ZN(new_n997));
  NOR3_X1   g811(.A1(new_n996), .A2(new_n997), .A3(new_n983), .ZN(G60));
  INV_X1    g812(.A(new_n983), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n986), .A2(new_n987), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n645), .A2(new_n647), .ZN(new_n1001));
  XOR2_X1   g815(.A(new_n649), .B(KEYINPUT59), .Z(new_n1002));
  NAND2_X1  g816(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n999), .B1(new_n1000), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n959), .A2(new_n965), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n1001), .B1(new_n1005), .B2(new_n1002), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n1004), .A2(new_n1006), .ZN(G63));
  NAND2_X1  g821(.A1(G217), .A2(G902), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1008), .B(KEYINPUT60), .ZN(new_n1009));
  INV_X1    g823(.A(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n677), .B(KEYINPUT121), .ZN(new_n1011));
  OAI211_X1 g825(.A(new_n1010), .B(new_n1011), .C1(new_n974), .C2(new_n958), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1009), .B1(new_n961), .B2(new_n964), .ZN(new_n1013));
  OAI211_X1 g827(.A(new_n1012), .B(new_n999), .C1(new_n1013), .C2(new_n376), .ZN(new_n1014));
  OAI211_X1 g828(.A(KEYINPUT122), .B(new_n999), .C1(new_n1013), .C2(new_n376), .ZN(new_n1015));
  INV_X1    g829(.A(KEYINPUT61), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n1014), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n1010), .B1(new_n974), .B2(new_n958), .ZN(new_n1018));
  INV_X1    g832(.A(new_n376), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n983), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  OAI211_X1 g834(.A(new_n1020), .B(new_n1012), .C1(KEYINPUT122), .C2(KEYINPUT61), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1017), .A2(new_n1021), .ZN(G66));
  INV_X1    g836(.A(new_n940), .ZN(new_n1023));
  AOI21_X1  g837(.A(G953), .B1(new_n957), .B2(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g838(.A(new_n1024), .B(KEYINPUT123), .ZN(new_n1025));
  OAI21_X1  g839(.A(G953), .B1(new_n572), .B2(new_n478), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g841(.A(new_n976), .B1(G898), .B2(new_n354), .ZN(new_n1028));
  XNOR2_X1  g842(.A(new_n1027), .B(new_n1028), .ZN(G69));
  NAND3_X1  g843(.A1(new_n724), .A2(new_n923), .A3(new_n729), .ZN(new_n1030));
  INV_X1    g844(.A(KEYINPUT124), .ZN(new_n1031));
  OR3_X1    g845(.A1(new_n1030), .A2(new_n1031), .A3(KEYINPUT62), .ZN(new_n1032));
  OAI21_X1  g846(.A(new_n1031), .B1(new_n1030), .B2(KEYINPUT62), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  AND2_X1   g848(.A1(new_n898), .A2(new_n899), .ZN(new_n1035));
  OAI211_X1 g849(.A(new_n713), .B(new_n830), .C1(new_n1035), .C2(new_n903), .ZN(new_n1036));
  NOR3_X1   g850(.A1(new_n1036), .A2(new_n744), .A3(new_n655), .ZN(new_n1037));
  AOI21_X1  g851(.A(new_n1037), .B1(new_n798), .B2(new_n816), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n1030), .A2(KEYINPUT62), .ZN(new_n1039));
  NAND4_X1  g853(.A1(new_n1034), .A2(new_n1038), .A3(new_n832), .A4(new_n1039), .ZN(new_n1040));
  NAND2_X1  g854(.A1(new_n1040), .A2(new_n354), .ZN(new_n1041));
  NOR2_X1   g855(.A1(new_n614), .A2(new_n615), .ZN(new_n1042));
  XNOR2_X1  g856(.A(new_n283), .B(new_n1042), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g858(.A(new_n1043), .B1(G900), .B2(G953), .ZN(new_n1045));
  INV_X1    g859(.A(new_n875), .ZN(new_n1046));
  INV_X1    g860(.A(KEYINPUT126), .ZN(new_n1047));
  NAND4_X1  g861(.A1(new_n816), .A2(new_n1046), .A3(new_n1047), .A4(new_n757), .ZN(new_n1048));
  NAND2_X1  g862(.A1(new_n1046), .A2(new_n757), .ZN(new_n1049));
  OAI21_X1  g863(.A(KEYINPUT126), .B1(new_n1049), .B2(new_n815), .ZN(new_n1050));
  NAND2_X1  g864(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1051));
  AND4_X1   g865(.A1(new_n729), .A2(new_n781), .A3(new_n927), .A4(new_n923), .ZN(new_n1052));
  NAND4_X1  g866(.A1(new_n1051), .A2(new_n817), .A3(new_n832), .A4(new_n1052), .ZN(new_n1053));
  OAI21_X1  g867(.A(new_n1045), .B1(new_n1053), .B2(G953), .ZN(new_n1054));
  NAND3_X1  g868(.A1(new_n1044), .A2(KEYINPUT125), .A3(new_n1054), .ZN(new_n1055));
  AOI21_X1  g869(.A(new_n354), .B1(G227), .B2(G900), .ZN(new_n1056));
  XNOR2_X1  g870(.A(new_n1055), .B(new_n1056), .ZN(G72));
  NAND2_X1  g871(.A1(G472), .A2(G902), .ZN(new_n1058));
  XOR2_X1   g872(.A(new_n1058), .B(KEYINPUT63), .Z(new_n1059));
  NAND2_X1  g873(.A1(new_n957), .A2(new_n1023), .ZN(new_n1060));
  OAI21_X1  g874(.A(new_n1059), .B1(new_n1040), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g875(.A1(new_n1061), .A2(new_n717), .ZN(new_n1062));
  INV_X1    g876(.A(new_n285), .ZN(new_n1063));
  NAND2_X1  g877(.A1(new_n284), .A2(new_n264), .ZN(new_n1064));
  NAND2_X1  g878(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  OAI211_X1 g879(.A(new_n1059), .B(new_n1065), .C1(new_n945), .C2(new_n958), .ZN(new_n1066));
  NAND3_X1  g880(.A1(new_n1062), .A2(new_n999), .A3(new_n1066), .ZN(new_n1067));
  OAI21_X1  g881(.A(new_n1059), .B1(new_n1053), .B2(new_n1060), .ZN(new_n1068));
  INV_X1    g882(.A(KEYINPUT127), .ZN(new_n1069));
  XNOR2_X1  g883(.A(new_n1068), .B(new_n1069), .ZN(new_n1070));
  AOI21_X1  g884(.A(new_n719), .B1(new_n283), .B2(new_n257), .ZN(new_n1071));
  AOI21_X1  g885(.A(new_n1067), .B1(new_n1070), .B2(new_n1071), .ZN(G57));
endmodule


