

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590;

  XNOR2_X1 U318 ( .A(n372), .B(n371), .ZN(n375) );
  XNOR2_X1 U319 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U320 ( .A(n421), .B(KEYINPUT119), .ZN(n422) );
  INV_X1 U321 ( .A(KEYINPUT48), .ZN(n400) );
  XNOR2_X1 U322 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U323 ( .A(n400), .B(KEYINPUT109), .ZN(n401) );
  XNOR2_X1 U324 ( .A(n402), .B(n401), .ZN(n530) );
  XNOR2_X1 U325 ( .A(KEYINPUT55), .B(KEYINPUT120), .ZN(n441) );
  XNOR2_X1 U326 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U327 ( .A(n442), .B(n441), .ZN(n457) );
  XNOR2_X1 U328 ( .A(n383), .B(n382), .ZN(n391) );
  XOR2_X1 U329 ( .A(n456), .B(n455), .Z(n532) );
  XOR2_X1 U330 ( .A(n472), .B(KEYINPUT28), .Z(n534) );
  XNOR2_X1 U331 ( .A(n458), .B(KEYINPUT58), .ZN(n459) );
  XNOR2_X1 U332 ( .A(n460), .B(n459), .ZN(G1351GAT) );
  XOR2_X1 U333 ( .A(KEYINPUT10), .B(KEYINPUT66), .Z(n287) );
  XNOR2_X1 U334 ( .A(G134GAT), .B(KEYINPUT11), .ZN(n286) );
  XNOR2_X1 U335 ( .A(n287), .B(n286), .ZN(n305) );
  XOR2_X1 U336 ( .A(KEYINPUT76), .B(G106GAT), .Z(n289) );
  XNOR2_X1 U337 ( .A(G36GAT), .B(G190GAT), .ZN(n288) );
  XOR2_X1 U338 ( .A(n289), .B(n288), .Z(n298) );
  INV_X1 U339 ( .A(n298), .ZN(n297) );
  INV_X1 U340 ( .A(G85GAT), .ZN(n290) );
  NAND2_X1 U341 ( .A1(G99GAT), .A2(n290), .ZN(n293) );
  INV_X1 U342 ( .A(G99GAT), .ZN(n291) );
  NAND2_X1 U343 ( .A1(n291), .A2(G85GAT), .ZN(n292) );
  NAND2_X1 U344 ( .A1(n293), .A2(n292), .ZN(n364) );
  XNOR2_X1 U345 ( .A(n364), .B(G92GAT), .ZN(n295) );
  XOR2_X1 U346 ( .A(G218GAT), .B(G162GAT), .Z(n294) );
  XNOR2_X1 U347 ( .A(n295), .B(n294), .ZN(n299) );
  INV_X1 U348 ( .A(n299), .ZN(n296) );
  NAND2_X1 U349 ( .A1(n297), .A2(n296), .ZN(n301) );
  NAND2_X1 U350 ( .A1(n299), .A2(n298), .ZN(n300) );
  NAND2_X1 U351 ( .A1(n301), .A2(n300), .ZN(n303) );
  NAND2_X1 U352 ( .A1(G232GAT), .A2(G233GAT), .ZN(n302) );
  XNOR2_X1 U353 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U354 ( .A(n305), .B(n304), .ZN(n313) );
  XOR2_X1 U355 ( .A(KEYINPUT8), .B(G50GAT), .Z(n307) );
  XNOR2_X1 U356 ( .A(G43GAT), .B(G29GAT), .ZN(n306) );
  XNOR2_X1 U357 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U358 ( .A(KEYINPUT7), .B(n308), .Z(n360) );
  XOR2_X1 U359 ( .A(KEYINPUT64), .B(KEYINPUT67), .Z(n310) );
  XNOR2_X1 U360 ( .A(KEYINPUT9), .B(KEYINPUT77), .ZN(n309) );
  XNOR2_X1 U361 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U362 ( .A(n360), .B(n311), .ZN(n312) );
  XNOR2_X1 U363 ( .A(n313), .B(n312), .ZN(n556) );
  INV_X1 U364 ( .A(n556), .ZN(n543) );
  XNOR2_X1 U365 ( .A(G120GAT), .B(G148GAT), .ZN(n314) );
  XNOR2_X1 U366 ( .A(n314), .B(G57GAT), .ZN(n377) );
  XOR2_X1 U367 ( .A(n377), .B(G85GAT), .Z(n316) );
  XOR2_X1 U368 ( .A(G113GAT), .B(G1GAT), .Z(n348) );
  XNOR2_X1 U369 ( .A(G29GAT), .B(n348), .ZN(n315) );
  XNOR2_X1 U370 ( .A(n316), .B(n315), .ZN(n321) );
  XNOR2_X1 U371 ( .A(G134GAT), .B(G127GAT), .ZN(n317) );
  XNOR2_X1 U372 ( .A(n317), .B(KEYINPUT0), .ZN(n443) );
  XOR2_X1 U373 ( .A(n443), .B(KEYINPUT1), .Z(n319) );
  NAND2_X1 U374 ( .A1(G225GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U375 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U376 ( .A(n321), .B(n320), .Z(n329) );
  XOR2_X1 U377 ( .A(KEYINPUT2), .B(G162GAT), .Z(n323) );
  XNOR2_X1 U378 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n322) );
  XNOR2_X1 U379 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U380 ( .A(G141GAT), .B(n324), .Z(n425) );
  XOR2_X1 U381 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n326) );
  XNOR2_X1 U382 ( .A(KEYINPUT88), .B(KEYINPUT6), .ZN(n325) );
  XNOR2_X1 U383 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U384 ( .A(n425), .B(n327), .ZN(n328) );
  XNOR2_X1 U385 ( .A(n329), .B(n328), .ZN(n468) );
  XNOR2_X1 U386 ( .A(KEYINPUT89), .B(n468), .ZN(n520) );
  INV_X1 U387 ( .A(KEYINPUT106), .ZN(n390) );
  XOR2_X1 U388 ( .A(G78GAT), .B(G211GAT), .Z(n331) );
  XNOR2_X1 U389 ( .A(G183GAT), .B(G127GAT), .ZN(n330) );
  XNOR2_X1 U390 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U391 ( .A(G71GAT), .B(KEYINPUT13), .Z(n373) );
  XOR2_X1 U392 ( .A(n332), .B(n373), .Z(n334) );
  XNOR2_X1 U393 ( .A(G1GAT), .B(G155GAT), .ZN(n333) );
  XNOR2_X1 U394 ( .A(n334), .B(n333), .ZN(n339) );
  XNOR2_X1 U395 ( .A(G15GAT), .B(G22GAT), .ZN(n335) );
  XNOR2_X1 U396 ( .A(n335), .B(KEYINPUT70), .ZN(n349) );
  XOR2_X1 U397 ( .A(n349), .B(KEYINPUT12), .Z(n337) );
  NAND2_X1 U398 ( .A1(G231GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U399 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U400 ( .A(n339), .B(n338), .Z(n347) );
  XOR2_X1 U401 ( .A(KEYINPUT80), .B(G64GAT), .Z(n341) );
  XNOR2_X1 U402 ( .A(G8GAT), .B(G57GAT), .ZN(n340) );
  XNOR2_X1 U403 ( .A(n341), .B(n340), .ZN(n345) );
  XOR2_X1 U404 ( .A(KEYINPUT79), .B(KEYINPUT15), .Z(n343) );
  XNOR2_X1 U405 ( .A(KEYINPUT78), .B(KEYINPUT14), .ZN(n342) );
  XNOR2_X1 U406 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U407 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U408 ( .A(n347), .B(n346), .Z(n583) );
  INV_X1 U409 ( .A(n583), .ZN(n570) );
  NAND2_X1 U410 ( .A1(n543), .A2(n570), .ZN(n387) );
  XOR2_X1 U411 ( .A(n349), .B(n348), .Z(n351) );
  XNOR2_X1 U412 ( .A(G197GAT), .B(G141GAT), .ZN(n350) );
  XNOR2_X1 U413 ( .A(n351), .B(n350), .ZN(n356) );
  XNOR2_X1 U414 ( .A(G169GAT), .B(G36GAT), .ZN(n352) );
  XNOR2_X1 U415 ( .A(n352), .B(G8GAT), .ZN(n415) );
  XOR2_X1 U416 ( .A(n415), .B(KEYINPUT68), .Z(n354) );
  NAND2_X1 U417 ( .A1(G229GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U418 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U419 ( .A(n356), .B(n355), .Z(n362) );
  XOR2_X1 U420 ( .A(KEYINPUT30), .B(KEYINPUT71), .Z(n358) );
  XNOR2_X1 U421 ( .A(KEYINPUT69), .B(KEYINPUT29), .ZN(n357) );
  XNOR2_X1 U422 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U423 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U424 ( .A(n362), .B(n361), .ZN(n575) );
  XNOR2_X1 U425 ( .A(G176GAT), .B(G92GAT), .ZN(n363) );
  XNOR2_X1 U426 ( .A(n363), .B(G64GAT), .ZN(n410) );
  NAND2_X1 U427 ( .A1(n410), .A2(n364), .ZN(n368) );
  INV_X1 U428 ( .A(n410), .ZN(n366) );
  INV_X1 U429 ( .A(n364), .ZN(n365) );
  NAND2_X1 U430 ( .A1(n366), .A2(n365), .ZN(n367) );
  NAND2_X1 U431 ( .A1(n368), .A2(n367), .ZN(n372) );
  AND2_X1 U432 ( .A1(G230GAT), .A2(G233GAT), .ZN(n370) );
  INV_X1 U433 ( .A(KEYINPUT73), .ZN(n369) );
  XNOR2_X1 U434 ( .A(G204GAT), .B(n373), .ZN(n374) );
  XNOR2_X1 U435 ( .A(n375), .B(n374), .ZN(n383) );
  XNOR2_X1 U436 ( .A(G106GAT), .B(G78GAT), .ZN(n376) );
  XNOR2_X1 U437 ( .A(n376), .B(KEYINPUT75), .ZN(n433) );
  XNOR2_X1 U438 ( .A(n433), .B(n377), .ZN(n381) );
  XOR2_X1 U439 ( .A(KEYINPUT32), .B(KEYINPUT31), .Z(n379) );
  XNOR2_X1 U440 ( .A(KEYINPUT74), .B(KEYINPUT33), .ZN(n378) );
  XOR2_X1 U441 ( .A(n379), .B(n378), .Z(n380) );
  XNOR2_X1 U442 ( .A(n391), .B(KEYINPUT41), .ZN(n563) );
  INV_X1 U443 ( .A(n563), .ZN(n552) );
  NAND2_X1 U444 ( .A1(n575), .A2(n552), .ZN(n385) );
  INV_X1 U445 ( .A(KEYINPUT46), .ZN(n384) );
  XNOR2_X1 U446 ( .A(n385), .B(n384), .ZN(n386) );
  NOR2_X1 U447 ( .A1(n387), .A2(n386), .ZN(n388) );
  XNOR2_X1 U448 ( .A(KEYINPUT47), .B(n388), .ZN(n389) );
  XNOR2_X1 U449 ( .A(n390), .B(n389), .ZN(n399) );
  XOR2_X1 U450 ( .A(KEYINPUT72), .B(n575), .Z(n560) );
  XOR2_X1 U451 ( .A(KEYINPUT107), .B(KEYINPUT45), .Z(n392) );
  XNOR2_X1 U452 ( .A(KEYINPUT65), .B(n392), .ZN(n394) );
  XOR2_X1 U453 ( .A(n556), .B(KEYINPUT36), .Z(n586) );
  NOR2_X1 U454 ( .A1(n586), .A2(n570), .ZN(n393) );
  XOR2_X1 U455 ( .A(n394), .B(n393), .Z(n395) );
  NAND2_X1 U456 ( .A1(n560), .A2(n395), .ZN(n396) );
  NOR2_X1 U457 ( .A1(n391), .A2(n396), .ZN(n397) );
  XNOR2_X1 U458 ( .A(KEYINPUT108), .B(n397), .ZN(n398) );
  NOR2_X1 U459 ( .A1(n399), .A2(n398), .ZN(n402) );
  INV_X1 U460 ( .A(n530), .ZN(n420) );
  XOR2_X1 U461 ( .A(G183GAT), .B(KEYINPUT82), .Z(n404) );
  XNOR2_X1 U462 ( .A(KEYINPUT19), .B(KEYINPUT17), .ZN(n403) );
  XNOR2_X1 U463 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U464 ( .A(n405), .B(KEYINPUT18), .Z(n407) );
  XNOR2_X1 U465 ( .A(KEYINPUT83), .B(G190GAT), .ZN(n406) );
  XNOR2_X1 U466 ( .A(n407), .B(n406), .ZN(n456) );
  XOR2_X1 U467 ( .A(KEYINPUT90), .B(KEYINPUT91), .Z(n409) );
  NAND2_X1 U468 ( .A1(G226GAT), .A2(G233GAT), .ZN(n408) );
  XNOR2_X1 U469 ( .A(n409), .B(n408), .ZN(n411) );
  XOR2_X1 U470 ( .A(n411), .B(n410), .Z(n417) );
  XOR2_X1 U471 ( .A(G211GAT), .B(G218GAT), .Z(n413) );
  XNOR2_X1 U472 ( .A(KEYINPUT21), .B(G204GAT), .ZN(n412) );
  XNOR2_X1 U473 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U474 ( .A(G197GAT), .B(n414), .Z(n426) );
  XNOR2_X1 U475 ( .A(n415), .B(n426), .ZN(n416) );
  XNOR2_X1 U476 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U477 ( .A(n456), .B(n418), .ZN(n523) );
  XOR2_X1 U478 ( .A(KEYINPUT117), .B(n523), .Z(n419) );
  NAND2_X1 U479 ( .A1(n420), .A2(n419), .ZN(n423) );
  XOR2_X1 U480 ( .A(KEYINPUT54), .B(KEYINPUT118), .Z(n421) );
  NOR2_X1 U481 ( .A1(n520), .A2(n424), .ZN(n572) );
  XNOR2_X1 U482 ( .A(n426), .B(n425), .ZN(n440) );
  XOR2_X1 U483 ( .A(KEYINPUT85), .B(G148GAT), .Z(n428) );
  XNOR2_X1 U484 ( .A(KEYINPUT84), .B(KEYINPUT86), .ZN(n427) );
  XNOR2_X1 U485 ( .A(n428), .B(n427), .ZN(n432) );
  XOR2_X1 U486 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n430) );
  XNOR2_X1 U487 ( .A(G22GAT), .B(KEYINPUT87), .ZN(n429) );
  XNOR2_X1 U488 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U489 ( .A(n432), .B(n431), .Z(n438) );
  XOR2_X1 U490 ( .A(KEYINPUT23), .B(n433), .Z(n435) );
  NAND2_X1 U491 ( .A1(G228GAT), .A2(G233GAT), .ZN(n434) );
  XNOR2_X1 U492 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U493 ( .A(G50GAT), .B(n436), .ZN(n437) );
  XNOR2_X1 U494 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U495 ( .A(n440), .B(n439), .ZN(n472) );
  NAND2_X1 U496 ( .A1(n572), .A2(n472), .ZN(n442) );
  XOR2_X1 U497 ( .A(n443), .B(G99GAT), .Z(n445) );
  NAND2_X1 U498 ( .A1(G227GAT), .A2(G233GAT), .ZN(n444) );
  XNOR2_X1 U499 ( .A(n445), .B(n444), .ZN(n449) );
  XOR2_X1 U500 ( .A(G120GAT), .B(G71GAT), .Z(n447) );
  XNOR2_X1 U501 ( .A(G113GAT), .B(G15GAT), .ZN(n446) );
  XNOR2_X1 U502 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U503 ( .A(n449), .B(n448), .Z(n454) );
  XOR2_X1 U504 ( .A(G176GAT), .B(KEYINPUT81), .Z(n451) );
  XNOR2_X1 U505 ( .A(G169GAT), .B(KEYINPUT20), .ZN(n450) );
  XNOR2_X1 U506 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U507 ( .A(G43GAT), .B(n452), .ZN(n453) );
  XNOR2_X1 U508 ( .A(n454), .B(n453), .ZN(n455) );
  NAND2_X1 U509 ( .A1(n457), .A2(n532), .ZN(n569) );
  NOR2_X1 U510 ( .A1(n543), .A2(n569), .ZN(n460) );
  INV_X1 U511 ( .A(G190GAT), .ZN(n458) );
  NOR2_X1 U512 ( .A1(n560), .A2(n391), .ZN(n493) );
  INV_X1 U513 ( .A(n493), .ZN(n478) );
  NOR2_X1 U514 ( .A1(n570), .A2(n556), .ZN(n461) );
  XNOR2_X1 U515 ( .A(n461), .B(KEYINPUT16), .ZN(n477) );
  NOR2_X1 U516 ( .A1(n472), .A2(n532), .ZN(n462) );
  XNOR2_X1 U517 ( .A(n462), .B(KEYINPUT26), .ZN(n573) );
  XNOR2_X1 U518 ( .A(n523), .B(KEYINPUT92), .ZN(n463) );
  XNOR2_X1 U519 ( .A(KEYINPUT27), .B(n463), .ZN(n471) );
  NAND2_X1 U520 ( .A1(n573), .A2(n471), .ZN(n467) );
  NAND2_X1 U521 ( .A1(n532), .A2(n523), .ZN(n464) );
  NAND2_X1 U522 ( .A1(n472), .A2(n464), .ZN(n465) );
  XOR2_X1 U523 ( .A(KEYINPUT25), .B(n465), .Z(n466) );
  NAND2_X1 U524 ( .A1(n467), .A2(n466), .ZN(n469) );
  NAND2_X1 U525 ( .A1(n469), .A2(n468), .ZN(n470) );
  XOR2_X1 U526 ( .A(KEYINPUT93), .B(n470), .Z(n476) );
  NAND2_X1 U527 ( .A1(n520), .A2(n471), .ZN(n529) );
  NOR2_X1 U528 ( .A1(n532), .A2(n529), .ZN(n474) );
  INV_X1 U529 ( .A(n534), .ZN(n473) );
  NAND2_X1 U530 ( .A1(n474), .A2(n473), .ZN(n475) );
  NAND2_X1 U531 ( .A1(n476), .A2(n475), .ZN(n488) );
  NAND2_X1 U532 ( .A1(n477), .A2(n488), .ZN(n505) );
  NOR2_X1 U533 ( .A1(n478), .A2(n505), .ZN(n486) );
  NAND2_X1 U534 ( .A1(n520), .A2(n486), .ZN(n479) );
  XNOR2_X1 U535 ( .A(n479), .B(KEYINPUT34), .ZN(n480) );
  XNOR2_X1 U536 ( .A(G1GAT), .B(n480), .ZN(G1324GAT) );
  NAND2_X1 U537 ( .A1(n523), .A2(n486), .ZN(n481) );
  XNOR2_X1 U538 ( .A(n481), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U539 ( .A(KEYINPUT35), .B(KEYINPUT95), .Z(n483) );
  NAND2_X1 U540 ( .A1(n486), .A2(n532), .ZN(n482) );
  XNOR2_X1 U541 ( .A(n483), .B(n482), .ZN(n485) );
  XOR2_X1 U542 ( .A(G15GAT), .B(KEYINPUT94), .Z(n484) );
  XNOR2_X1 U543 ( .A(n485), .B(n484), .ZN(G1326GAT) );
  NAND2_X1 U544 ( .A1(n486), .A2(n534), .ZN(n487) );
  XNOR2_X1 U545 ( .A(n487), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U546 ( .A(KEYINPUT39), .B(KEYINPUT98), .Z(n496) );
  NAND2_X1 U547 ( .A1(n570), .A2(n488), .ZN(n489) );
  XNOR2_X1 U548 ( .A(KEYINPUT96), .B(n489), .ZN(n490) );
  NOR2_X1 U549 ( .A1(n586), .A2(n490), .ZN(n492) );
  XNOR2_X1 U550 ( .A(KEYINPUT97), .B(KEYINPUT37), .ZN(n491) );
  XNOR2_X1 U551 ( .A(n492), .B(n491), .ZN(n517) );
  NAND2_X1 U552 ( .A1(n517), .A2(n493), .ZN(n494) );
  XOR2_X1 U553 ( .A(KEYINPUT38), .B(n494), .Z(n501) );
  NAND2_X1 U554 ( .A1(n501), .A2(n520), .ZN(n495) );
  XNOR2_X1 U555 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U556 ( .A(G29GAT), .B(n497), .ZN(G1328GAT) );
  NAND2_X1 U557 ( .A1(n501), .A2(n523), .ZN(n498) );
  XNOR2_X1 U558 ( .A(n498), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U559 ( .A1(n501), .A2(n532), .ZN(n499) );
  XNOR2_X1 U560 ( .A(n499), .B(KEYINPUT40), .ZN(n500) );
  XNOR2_X1 U561 ( .A(G43GAT), .B(n500), .ZN(G1330GAT) );
  XOR2_X1 U562 ( .A(G50GAT), .B(KEYINPUT99), .Z(n503) );
  NAND2_X1 U563 ( .A1(n534), .A2(n501), .ZN(n502) );
  XNOR2_X1 U564 ( .A(n503), .B(n502), .ZN(G1331GAT) );
  NOR2_X1 U565 ( .A1(n563), .A2(n575), .ZN(n504) );
  XOR2_X1 U566 ( .A(n504), .B(KEYINPUT100), .Z(n516) );
  NOR2_X1 U567 ( .A1(n516), .A2(n505), .ZN(n513) );
  NAND2_X1 U568 ( .A1(n520), .A2(n513), .ZN(n509) );
  XOR2_X1 U569 ( .A(KEYINPUT102), .B(KEYINPUT42), .Z(n507) );
  XNOR2_X1 U570 ( .A(G57GAT), .B(KEYINPUT101), .ZN(n506) );
  XNOR2_X1 U571 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U572 ( .A(n509), .B(n508), .ZN(G1332GAT) );
  XOR2_X1 U573 ( .A(G64GAT), .B(KEYINPUT103), .Z(n511) );
  NAND2_X1 U574 ( .A1(n513), .A2(n523), .ZN(n510) );
  XNOR2_X1 U575 ( .A(n511), .B(n510), .ZN(G1333GAT) );
  NAND2_X1 U576 ( .A1(n513), .A2(n532), .ZN(n512) );
  XNOR2_X1 U577 ( .A(n512), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U578 ( .A(G78GAT), .B(KEYINPUT43), .Z(n515) );
  NAND2_X1 U579 ( .A1(n513), .A2(n534), .ZN(n514) );
  XNOR2_X1 U580 ( .A(n515), .B(n514), .ZN(G1335GAT) );
  INV_X1 U581 ( .A(n516), .ZN(n518) );
  NAND2_X1 U582 ( .A1(n518), .A2(n517), .ZN(n519) );
  XOR2_X1 U583 ( .A(KEYINPUT104), .B(n519), .Z(n526) );
  NAND2_X1 U584 ( .A1(n526), .A2(n520), .ZN(n521) );
  XOR2_X1 U585 ( .A(KEYINPUT105), .B(n521), .Z(n522) );
  XNOR2_X1 U586 ( .A(G85GAT), .B(n522), .ZN(G1336GAT) );
  NAND2_X1 U587 ( .A1(n526), .A2(n523), .ZN(n524) );
  XNOR2_X1 U588 ( .A(n524), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U589 ( .A1(n526), .A2(n532), .ZN(n525) );
  XNOR2_X1 U590 ( .A(n525), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U591 ( .A1(n526), .A2(n534), .ZN(n527) );
  XNOR2_X1 U592 ( .A(n527), .B(KEYINPUT44), .ZN(n528) );
  XNOR2_X1 U593 ( .A(G106GAT), .B(n528), .ZN(G1339GAT) );
  NOR2_X1 U594 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U595 ( .A(KEYINPUT110), .B(n531), .ZN(n546) );
  NAND2_X1 U596 ( .A1(n532), .A2(n546), .ZN(n533) );
  NOR2_X1 U597 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U598 ( .A(KEYINPUT111), .B(n535), .ZN(n542) );
  NOR2_X1 U599 ( .A1(n560), .A2(n542), .ZN(n536) );
  XOR2_X1 U600 ( .A(KEYINPUT112), .B(n536), .Z(n537) );
  XNOR2_X1 U601 ( .A(G113GAT), .B(n537), .ZN(G1340GAT) );
  NOR2_X1 U602 ( .A1(n563), .A2(n542), .ZN(n539) );
  XNOR2_X1 U603 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n538) );
  XNOR2_X1 U604 ( .A(n539), .B(n538), .ZN(G1341GAT) );
  NOR2_X1 U605 ( .A1(n570), .A2(n542), .ZN(n540) );
  XOR2_X1 U606 ( .A(KEYINPUT50), .B(n540), .Z(n541) );
  XNOR2_X1 U607 ( .A(G127GAT), .B(n541), .ZN(G1342GAT) );
  NOR2_X1 U608 ( .A1(n543), .A2(n542), .ZN(n545) );
  XNOR2_X1 U609 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n544) );
  XNOR2_X1 U610 ( .A(n545), .B(n544), .ZN(G1343GAT) );
  XOR2_X1 U611 ( .A(G141GAT), .B(KEYINPUT113), .Z(n548) );
  AND2_X1 U612 ( .A1(n573), .A2(n546), .ZN(n557) );
  NAND2_X1 U613 ( .A1(n557), .A2(n575), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n548), .B(n547), .ZN(G1344GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT115), .B(KEYINPUT53), .Z(n550) );
  XNOR2_X1 U616 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n550), .B(n549), .ZN(n551) );
  XOR2_X1 U618 ( .A(KEYINPUT114), .B(n551), .Z(n554) );
  NAND2_X1 U619 ( .A1(n557), .A2(n552), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n554), .B(n553), .ZN(G1345GAT) );
  NAND2_X1 U621 ( .A1(n583), .A2(n557), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n555), .B(G155GAT), .ZN(G1346GAT) );
  XNOR2_X1 U623 ( .A(G162GAT), .B(KEYINPUT116), .ZN(n559) );
  NAND2_X1 U624 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n559), .B(n558), .ZN(G1347GAT) );
  NOR2_X1 U626 ( .A1(n560), .A2(n569), .ZN(n562) );
  XNOR2_X1 U627 ( .A(G169GAT), .B(KEYINPUT121), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(G1348GAT) );
  NOR2_X1 U629 ( .A1(n563), .A2(n569), .ZN(n568) );
  XOR2_X1 U630 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n565) );
  XNOR2_X1 U631 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U633 ( .A(KEYINPUT122), .B(n566), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(G1349GAT) );
  NOR2_X1 U635 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U636 ( .A(G183GAT), .B(n571), .Z(G1350GAT) );
  XOR2_X1 U637 ( .A(G197GAT), .B(KEYINPUT60), .Z(n577) );
  NAND2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U639 ( .A(KEYINPUT124), .B(n574), .ZN(n587) );
  INV_X1 U640 ( .A(n587), .ZN(n584) );
  NAND2_X1 U641 ( .A1(n575), .A2(n584), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n579) );
  XOR2_X1 U643 ( .A(KEYINPUT59), .B(KEYINPUT125), .Z(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1352GAT) );
  XOR2_X1 U645 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n581) );
  NAND2_X1 U646 ( .A1(n391), .A2(n584), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U648 ( .A(G204GAT), .B(n582), .ZN(G1353GAT) );
  NAND2_X1 U649 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n585), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U651 ( .A1(n587), .A2(n586), .ZN(n589) );
  XNOR2_X1 U652 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n589), .B(n588), .ZN(n590) );
  XNOR2_X1 U654 ( .A(G218GAT), .B(n590), .ZN(G1355GAT) );
endmodule

