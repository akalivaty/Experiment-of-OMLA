

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U550 ( .A(KEYINPUT31), .ZN(n721) );
  XNOR2_X1 U551 ( .A(n721), .B(KEYINPUT102), .ZN(n722) );
  XNOR2_X1 U552 ( .A(n723), .B(n722), .ZN(n724) );
  OR2_X1 U553 ( .A1(n681), .A2(n680), .ZN(n727) );
  NOR2_X1 U554 ( .A1(G1384), .A2(G164), .ZN(n678) );
  NOR2_X1 U555 ( .A1(G651), .A2(n626), .ZN(n637) );
  XNOR2_X1 U556 ( .A(KEYINPUT65), .B(n526), .ZN(G160) );
  AND2_X1 U557 ( .A1(G2104), .A2(G2105), .ZN(n877) );
  NAND2_X1 U558 ( .A1(G113), .A2(n877), .ZN(n516) );
  XNOR2_X1 U559 ( .A(n516), .B(KEYINPUT66), .ZN(n525) );
  INV_X1 U560 ( .A(G2104), .ZN(n520) );
  AND2_X1 U561 ( .A1(n520), .A2(G2105), .ZN(n876) );
  NAND2_X1 U562 ( .A1(G125), .A2(n876), .ZN(n519) );
  NOR2_X1 U563 ( .A1(G2104), .A2(G2105), .ZN(n517) );
  XOR2_X2 U564 ( .A(KEYINPUT17), .B(n517), .Z(n883) );
  NAND2_X1 U565 ( .A1(G137), .A2(n883), .ZN(n518) );
  NAND2_X1 U566 ( .A1(n519), .A2(n518), .ZN(n523) );
  NOR2_X2 U567 ( .A1(G2105), .A2(n520), .ZN(n881) );
  NAND2_X1 U568 ( .A1(G101), .A2(n881), .ZN(n521) );
  XNOR2_X1 U569 ( .A(KEYINPUT23), .B(n521), .ZN(n522) );
  NOR2_X1 U570 ( .A1(n523), .A2(n522), .ZN(n524) );
  NAND2_X1 U571 ( .A1(n525), .A2(n524), .ZN(n526) );
  NAND2_X1 U572 ( .A1(G138), .A2(n883), .ZN(n527) );
  XNOR2_X1 U573 ( .A(n527), .B(KEYINPUT90), .ZN(n533) );
  AND2_X1 U574 ( .A1(n876), .A2(G126), .ZN(n531) );
  NAND2_X1 U575 ( .A1(G114), .A2(n877), .ZN(n529) );
  NAND2_X1 U576 ( .A1(G102), .A2(n881), .ZN(n528) );
  NAND2_X1 U577 ( .A1(n529), .A2(n528), .ZN(n530) );
  NOR2_X1 U578 ( .A1(n531), .A2(n530), .ZN(n532) );
  AND2_X1 U579 ( .A1(n533), .A2(n532), .ZN(G164) );
  NOR2_X1 U580 ( .A1(G651), .A2(G543), .ZN(n644) );
  NAND2_X1 U581 ( .A1(G85), .A2(n644), .ZN(n536) );
  INV_X1 U582 ( .A(G651), .ZN(n537) );
  NOR2_X1 U583 ( .A1(G543), .A2(n537), .ZN(n534) );
  XOR2_X2 U584 ( .A(KEYINPUT1), .B(n534), .Z(n641) );
  NAND2_X1 U585 ( .A1(G60), .A2(n641), .ZN(n535) );
  NAND2_X1 U586 ( .A1(n536), .A2(n535), .ZN(n541) );
  XOR2_X1 U587 ( .A(KEYINPUT0), .B(G543), .Z(n626) );
  NOR2_X1 U588 ( .A1(n626), .A2(n537), .ZN(n639) );
  NAND2_X1 U589 ( .A1(G72), .A2(n639), .ZN(n539) );
  NAND2_X1 U590 ( .A1(G47), .A2(n637), .ZN(n538) );
  NAND2_X1 U591 ( .A1(n539), .A2(n538), .ZN(n540) );
  OR2_X1 U592 ( .A1(n541), .A2(n540), .ZN(G290) );
  AND2_X1 U593 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U594 ( .A1(G123), .A2(n876), .ZN(n542) );
  XNOR2_X1 U595 ( .A(n542), .B(KEYINPUT18), .ZN(n549) );
  NAND2_X1 U596 ( .A1(G111), .A2(n877), .ZN(n544) );
  NAND2_X1 U597 ( .A1(G135), .A2(n883), .ZN(n543) );
  NAND2_X1 U598 ( .A1(n544), .A2(n543), .ZN(n547) );
  NAND2_X1 U599 ( .A1(G99), .A2(n881), .ZN(n545) );
  XNOR2_X1 U600 ( .A(KEYINPUT79), .B(n545), .ZN(n546) );
  NOR2_X1 U601 ( .A1(n547), .A2(n546), .ZN(n548) );
  NAND2_X1 U602 ( .A1(n549), .A2(n548), .ZN(n997) );
  XNOR2_X1 U603 ( .A(G2096), .B(n997), .ZN(n550) );
  OR2_X1 U604 ( .A1(G2100), .A2(n550), .ZN(G156) );
  INV_X1 U605 ( .A(G57), .ZN(G237) );
  INV_X1 U606 ( .A(G132), .ZN(G219) );
  INV_X1 U607 ( .A(G82), .ZN(G220) );
  NAND2_X1 U608 ( .A1(n644), .A2(G89), .ZN(n551) );
  XNOR2_X1 U609 ( .A(KEYINPUT4), .B(n551), .ZN(n554) );
  NAND2_X1 U610 ( .A1(n639), .A2(G76), .ZN(n552) );
  XOR2_X1 U611 ( .A(KEYINPUT77), .B(n552), .Z(n553) );
  NAND2_X1 U612 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U613 ( .A(n555), .B(KEYINPUT5), .ZN(n560) );
  NAND2_X1 U614 ( .A1(G63), .A2(n641), .ZN(n557) );
  NAND2_X1 U615 ( .A1(G51), .A2(n637), .ZN(n556) );
  NAND2_X1 U616 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U617 ( .A(KEYINPUT6), .B(n558), .Z(n559) );
  NAND2_X1 U618 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U619 ( .A(n561), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U620 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U621 ( .A1(G7), .A2(G661), .ZN(n562) );
  XNOR2_X1 U622 ( .A(n562), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U623 ( .A(G223), .ZN(n821) );
  NAND2_X1 U624 ( .A1(n821), .A2(G567), .ZN(n563) );
  XOR2_X1 U625 ( .A(KEYINPUT11), .B(n563), .Z(G234) );
  NAND2_X1 U626 ( .A1(G56), .A2(n641), .ZN(n564) );
  XOR2_X1 U627 ( .A(KEYINPUT14), .B(n564), .Z(n570) );
  NAND2_X1 U628 ( .A1(n644), .A2(G81), .ZN(n565) );
  XNOR2_X1 U629 ( .A(n565), .B(KEYINPUT12), .ZN(n567) );
  NAND2_X1 U630 ( .A1(G68), .A2(n639), .ZN(n566) );
  NAND2_X1 U631 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U632 ( .A(KEYINPUT13), .B(n568), .Z(n569) );
  NOR2_X1 U633 ( .A1(n570), .A2(n569), .ZN(n572) );
  NAND2_X1 U634 ( .A1(n637), .A2(G43), .ZN(n571) );
  NAND2_X1 U635 ( .A1(n572), .A2(n571), .ZN(n978) );
  XOR2_X1 U636 ( .A(G860), .B(KEYINPUT72), .Z(n605) );
  NOR2_X1 U637 ( .A1(n978), .A2(n605), .ZN(n573) );
  XNOR2_X1 U638 ( .A(n573), .B(KEYINPUT73), .ZN(G153) );
  NAND2_X1 U639 ( .A1(n637), .A2(G52), .ZN(n574) );
  XNOR2_X1 U640 ( .A(KEYINPUT67), .B(n574), .ZN(n580) );
  NAND2_X1 U641 ( .A1(G90), .A2(n644), .ZN(n576) );
  NAND2_X1 U642 ( .A1(G77), .A2(n639), .ZN(n575) );
  NAND2_X1 U643 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U644 ( .A(KEYINPUT9), .B(n577), .Z(n578) );
  XNOR2_X1 U645 ( .A(KEYINPUT68), .B(n578), .ZN(n579) );
  NOR2_X1 U646 ( .A1(n580), .A2(n579), .ZN(n582) );
  NAND2_X1 U647 ( .A1(n641), .A2(G64), .ZN(n581) );
  NAND2_X1 U648 ( .A1(n582), .A2(n581), .ZN(G301) );
  NAND2_X1 U649 ( .A1(G54), .A2(n637), .ZN(n589) );
  NAND2_X1 U650 ( .A1(G92), .A2(n644), .ZN(n584) );
  NAND2_X1 U651 ( .A1(G79), .A2(n639), .ZN(n583) );
  NAND2_X1 U652 ( .A1(n584), .A2(n583), .ZN(n587) );
  NAND2_X1 U653 ( .A1(n641), .A2(G66), .ZN(n585) );
  XOR2_X1 U654 ( .A(KEYINPUT74), .B(n585), .Z(n586) );
  NOR2_X1 U655 ( .A1(n587), .A2(n586), .ZN(n588) );
  NAND2_X1 U656 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U657 ( .A(n590), .B(KEYINPUT15), .ZN(n591) );
  XOR2_X1 U658 ( .A(KEYINPUT75), .B(n591), .Z(n963) );
  INV_X1 U659 ( .A(n963), .ZN(n696) );
  INV_X1 U660 ( .A(G868), .ZN(n659) );
  NAND2_X1 U661 ( .A1(n696), .A2(n659), .ZN(n592) );
  XNOR2_X1 U662 ( .A(n592), .B(KEYINPUT76), .ZN(n594) );
  NAND2_X1 U663 ( .A1(G868), .A2(G301), .ZN(n593) );
  NAND2_X1 U664 ( .A1(n594), .A2(n593), .ZN(G284) );
  NAND2_X1 U665 ( .A1(G53), .A2(n637), .ZN(n595) );
  XNOR2_X1 U666 ( .A(n595), .B(KEYINPUT70), .ZN(n598) );
  NAND2_X1 U667 ( .A1(G78), .A2(n639), .ZN(n596) );
  XOR2_X1 U668 ( .A(KEYINPUT69), .B(n596), .Z(n597) );
  NAND2_X1 U669 ( .A1(n598), .A2(n597), .ZN(n602) );
  NAND2_X1 U670 ( .A1(G91), .A2(n644), .ZN(n600) );
  NAND2_X1 U671 ( .A1(G65), .A2(n641), .ZN(n599) );
  NAND2_X1 U672 ( .A1(n600), .A2(n599), .ZN(n601) );
  NOR2_X1 U673 ( .A1(n602), .A2(n601), .ZN(n975) );
  XNOR2_X1 U674 ( .A(n975), .B(KEYINPUT71), .ZN(G299) );
  NAND2_X1 U675 ( .A1(G286), .A2(G868), .ZN(n604) );
  NAND2_X1 U676 ( .A1(G299), .A2(n659), .ZN(n603) );
  NAND2_X1 U677 ( .A1(n604), .A2(n603), .ZN(G297) );
  NAND2_X1 U678 ( .A1(n605), .A2(G559), .ZN(n606) );
  NAND2_X1 U679 ( .A1(n606), .A2(n963), .ZN(n607) );
  XNOR2_X1 U680 ( .A(n607), .B(KEYINPUT16), .ZN(n608) );
  XNOR2_X1 U681 ( .A(KEYINPUT78), .B(n608), .ZN(G148) );
  NOR2_X1 U682 ( .A1(G868), .A2(n978), .ZN(n611) );
  NAND2_X1 U683 ( .A1(G868), .A2(n963), .ZN(n609) );
  NOR2_X1 U684 ( .A1(G559), .A2(n609), .ZN(n610) );
  NOR2_X1 U685 ( .A1(n611), .A2(n610), .ZN(G282) );
  NAND2_X1 U686 ( .A1(n963), .A2(G559), .ZN(n657) );
  XNOR2_X1 U687 ( .A(n978), .B(n657), .ZN(n612) );
  NOR2_X1 U688 ( .A1(G860), .A2(n612), .ZN(n622) );
  NAND2_X1 U689 ( .A1(n644), .A2(G93), .ZN(n613) );
  XOR2_X1 U690 ( .A(KEYINPUT81), .B(n613), .Z(n615) );
  NAND2_X1 U691 ( .A1(n639), .A2(G80), .ZN(n614) );
  NAND2_X1 U692 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U693 ( .A(KEYINPUT82), .B(n616), .ZN(n620) );
  NAND2_X1 U694 ( .A1(G67), .A2(n641), .ZN(n618) );
  NAND2_X1 U695 ( .A1(G55), .A2(n637), .ZN(n617) );
  NAND2_X1 U696 ( .A1(n618), .A2(n617), .ZN(n619) );
  OR2_X1 U697 ( .A1(n620), .A2(n619), .ZN(n660) );
  XOR2_X1 U698 ( .A(n660), .B(KEYINPUT80), .Z(n621) );
  XNOR2_X1 U699 ( .A(n622), .B(n621), .ZN(G145) );
  NAND2_X1 U700 ( .A1(G49), .A2(n637), .ZN(n624) );
  NAND2_X1 U701 ( .A1(G74), .A2(G651), .ZN(n623) );
  NAND2_X1 U702 ( .A1(n624), .A2(n623), .ZN(n625) );
  XNOR2_X1 U703 ( .A(KEYINPUT83), .B(n625), .ZN(n630) );
  NAND2_X1 U704 ( .A1(G87), .A2(n626), .ZN(n627) );
  XOR2_X1 U705 ( .A(KEYINPUT84), .B(n627), .Z(n628) );
  NOR2_X1 U706 ( .A1(n641), .A2(n628), .ZN(n629) );
  NAND2_X1 U707 ( .A1(n630), .A2(n629), .ZN(G288) );
  NAND2_X1 U708 ( .A1(G88), .A2(n644), .ZN(n632) );
  NAND2_X1 U709 ( .A1(G75), .A2(n639), .ZN(n631) );
  NAND2_X1 U710 ( .A1(n632), .A2(n631), .ZN(n636) );
  NAND2_X1 U711 ( .A1(G62), .A2(n641), .ZN(n634) );
  NAND2_X1 U712 ( .A1(G50), .A2(n637), .ZN(n633) );
  NAND2_X1 U713 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U714 ( .A1(n636), .A2(n635), .ZN(G166) );
  NAND2_X1 U715 ( .A1(G48), .A2(n637), .ZN(n638) );
  XNOR2_X1 U716 ( .A(n638), .B(KEYINPUT86), .ZN(n649) );
  NAND2_X1 U717 ( .A1(n639), .A2(G73), .ZN(n640) );
  XNOR2_X1 U718 ( .A(n640), .B(KEYINPUT2), .ZN(n643) );
  NAND2_X1 U719 ( .A1(G61), .A2(n641), .ZN(n642) );
  NAND2_X1 U720 ( .A1(n643), .A2(n642), .ZN(n647) );
  NAND2_X1 U721 ( .A1(G86), .A2(n644), .ZN(n645) );
  XNOR2_X1 U722 ( .A(KEYINPUT85), .B(n645), .ZN(n646) );
  NOR2_X1 U723 ( .A1(n647), .A2(n646), .ZN(n648) );
  NAND2_X1 U724 ( .A1(n649), .A2(n648), .ZN(G305) );
  XOR2_X1 U725 ( .A(KEYINPUT87), .B(KEYINPUT19), .Z(n650) );
  XNOR2_X1 U726 ( .A(G288), .B(n650), .ZN(n651) );
  XOR2_X1 U727 ( .A(n660), .B(n651), .Z(n653) );
  XNOR2_X1 U728 ( .A(n978), .B(G166), .ZN(n652) );
  XNOR2_X1 U729 ( .A(n653), .B(n652), .ZN(n654) );
  XNOR2_X1 U730 ( .A(n654), .B(G305), .ZN(n655) );
  XNOR2_X1 U731 ( .A(n655), .B(G290), .ZN(n656) );
  XNOR2_X1 U732 ( .A(n656), .B(G299), .ZN(n894) );
  XOR2_X1 U733 ( .A(n894), .B(n657), .Z(n658) );
  NAND2_X1 U734 ( .A1(G868), .A2(n658), .ZN(n662) );
  NAND2_X1 U735 ( .A1(n660), .A2(n659), .ZN(n661) );
  NAND2_X1 U736 ( .A1(n662), .A2(n661), .ZN(G295) );
  XOR2_X1 U737 ( .A(KEYINPUT88), .B(KEYINPUT20), .Z(n664) );
  NAND2_X1 U738 ( .A1(G2078), .A2(G2084), .ZN(n663) );
  XNOR2_X1 U739 ( .A(n664), .B(n663), .ZN(n665) );
  NAND2_X1 U740 ( .A1(G2090), .A2(n665), .ZN(n666) );
  XNOR2_X1 U741 ( .A(KEYINPUT21), .B(n666), .ZN(n667) );
  NAND2_X1 U742 ( .A1(n667), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U743 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U744 ( .A1(G220), .A2(G219), .ZN(n668) );
  XOR2_X1 U745 ( .A(KEYINPUT22), .B(n668), .Z(n669) );
  NOR2_X1 U746 ( .A1(G218), .A2(n669), .ZN(n670) );
  NAND2_X1 U747 ( .A1(G96), .A2(n670), .ZN(n826) );
  NAND2_X1 U748 ( .A1(G2106), .A2(n826), .ZN(n674) );
  NAND2_X1 U749 ( .A1(G120), .A2(G108), .ZN(n671) );
  NOR2_X1 U750 ( .A1(G237), .A2(n671), .ZN(n672) );
  NAND2_X1 U751 ( .A1(G69), .A2(n672), .ZN(n827) );
  NAND2_X1 U752 ( .A1(G567), .A2(n827), .ZN(n673) );
  NAND2_X1 U753 ( .A1(n674), .A2(n673), .ZN(n675) );
  XNOR2_X1 U754 ( .A(KEYINPUT89), .B(n675), .ZN(G319) );
  INV_X1 U755 ( .A(G319), .ZN(n677) );
  NAND2_X1 U756 ( .A1(G661), .A2(G483), .ZN(n676) );
  NOR2_X1 U757 ( .A1(n677), .A2(n676), .ZN(n825) );
  NAND2_X1 U758 ( .A1(n825), .A2(G36), .ZN(G176) );
  INV_X1 U759 ( .A(G166), .ZN(G303) );
  XNOR2_X1 U760 ( .A(KEYINPUT106), .B(KEYINPUT40), .ZN(n820) );
  XNOR2_X1 U761 ( .A(G1986), .B(G290), .ZN(n967) );
  NAND2_X1 U762 ( .A1(G160), .A2(G40), .ZN(n680) );
  XNOR2_X1 U763 ( .A(n678), .B(KEYINPUT64), .ZN(n679) );
  NOR2_X1 U764 ( .A1(n680), .A2(n679), .ZN(n814) );
  NAND2_X1 U765 ( .A1(n967), .A2(n814), .ZN(n802) );
  INV_X1 U766 ( .A(n679), .ZN(n681) );
  NAND2_X1 U767 ( .A1(G8), .A2(n727), .ZN(n762) );
  NOR2_X1 U768 ( .A1(G1981), .A2(G305), .ZN(n682) );
  XOR2_X1 U769 ( .A(n682), .B(KEYINPUT24), .Z(n683) );
  NOR2_X1 U770 ( .A1(n762), .A2(n683), .ZN(n767) );
  INV_X1 U771 ( .A(n727), .ZN(n708) );
  NAND2_X1 U772 ( .A1(n708), .A2(G2072), .ZN(n684) );
  XNOR2_X1 U773 ( .A(n684), .B(KEYINPUT27), .ZN(n686) );
  INV_X1 U774 ( .A(G1956), .ZN(n916) );
  NOR2_X1 U775 ( .A1(n916), .A2(n708), .ZN(n685) );
  NOR2_X1 U776 ( .A1(n686), .A2(n685), .ZN(n702) );
  NOR2_X1 U777 ( .A1(n702), .A2(n975), .ZN(n687) );
  XOR2_X1 U778 ( .A(n687), .B(KEYINPUT28), .Z(n706) );
  INV_X1 U779 ( .A(G1996), .ZN(n939) );
  OR2_X1 U780 ( .A1(n727), .A2(n939), .ZN(n688) );
  XNOR2_X1 U781 ( .A(n688), .B(KEYINPUT26), .ZN(n690) );
  NAND2_X1 U782 ( .A1(n727), .A2(G1341), .ZN(n689) );
  NAND2_X1 U783 ( .A1(n690), .A2(n689), .ZN(n691) );
  NOR2_X1 U784 ( .A1(n691), .A2(n978), .ZN(n695) );
  NOR2_X1 U785 ( .A1(n708), .A2(G1348), .ZN(n693) );
  NOR2_X1 U786 ( .A1(G2067), .A2(n727), .ZN(n692) );
  NOR2_X1 U787 ( .A1(n693), .A2(n692), .ZN(n697) );
  NAND2_X1 U788 ( .A1(n696), .A2(n697), .ZN(n694) );
  NAND2_X1 U789 ( .A1(n695), .A2(n694), .ZN(n699) );
  OR2_X1 U790 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U791 ( .A1(n699), .A2(n698), .ZN(n701) );
  INV_X1 U792 ( .A(KEYINPUT100), .ZN(n700) );
  XNOR2_X1 U793 ( .A(n701), .B(n700), .ZN(n704) );
  NAND2_X1 U794 ( .A1(n702), .A2(n975), .ZN(n703) );
  NAND2_X1 U795 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U796 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U797 ( .A(n707), .B(KEYINPUT29), .ZN(n712) );
  XOR2_X1 U798 ( .A(G2078), .B(KEYINPUT25), .Z(n944) );
  NOR2_X1 U799 ( .A1(n944), .A2(n727), .ZN(n710) );
  NOR2_X1 U800 ( .A1(n708), .A2(G1961), .ZN(n709) );
  NOR2_X1 U801 ( .A1(n710), .A2(n709), .ZN(n718) );
  NOR2_X1 U802 ( .A1(G301), .A2(n718), .ZN(n711) );
  NOR2_X1 U803 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U804 ( .A(n713), .B(KEYINPUT101), .ZN(n725) );
  NOR2_X1 U805 ( .A1(G1966), .A2(n762), .ZN(n740) );
  NOR2_X1 U806 ( .A1(G2084), .A2(n727), .ZN(n714) );
  XOR2_X1 U807 ( .A(KEYINPUT98), .B(n714), .Z(n736) );
  NAND2_X1 U808 ( .A1(G8), .A2(n736), .ZN(n715) );
  NOR2_X1 U809 ( .A1(n740), .A2(n715), .ZN(n716) );
  XOR2_X1 U810 ( .A(KEYINPUT30), .B(n716), .Z(n717) );
  NOR2_X1 U811 ( .A1(G168), .A2(n717), .ZN(n720) );
  AND2_X1 U812 ( .A1(G301), .A2(n718), .ZN(n719) );
  NOR2_X1 U813 ( .A1(n720), .A2(n719), .ZN(n723) );
  NAND2_X1 U814 ( .A1(n725), .A2(n724), .ZN(n741) );
  AND2_X1 U815 ( .A1(G286), .A2(G8), .ZN(n726) );
  NAND2_X1 U816 ( .A1(n741), .A2(n726), .ZN(n734) );
  INV_X1 U817 ( .A(G8), .ZN(n732) );
  NOR2_X1 U818 ( .A1(G1971), .A2(n762), .ZN(n729) );
  NOR2_X1 U819 ( .A1(G2090), .A2(n727), .ZN(n728) );
  NOR2_X1 U820 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U821 ( .A1(n730), .A2(G303), .ZN(n731) );
  OR2_X1 U822 ( .A1(n732), .A2(n731), .ZN(n733) );
  AND2_X1 U823 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U824 ( .A(n735), .B(KEYINPUT32), .ZN(n758) );
  INV_X1 U825 ( .A(n736), .ZN(n737) );
  NAND2_X1 U826 ( .A1(G8), .A2(n737), .ZN(n738) );
  XNOR2_X1 U827 ( .A(KEYINPUT99), .B(n738), .ZN(n739) );
  NOR2_X1 U828 ( .A1(n740), .A2(n739), .ZN(n742) );
  NAND2_X1 U829 ( .A1(n742), .A2(n741), .ZN(n757) );
  NAND2_X1 U830 ( .A1(G1976), .A2(G288), .ZN(n968) );
  AND2_X1 U831 ( .A1(n757), .A2(n968), .ZN(n743) );
  NAND2_X1 U832 ( .A1(n758), .A2(n743), .ZN(n750) );
  INV_X1 U833 ( .A(n968), .ZN(n745) );
  NOR2_X1 U834 ( .A1(G1976), .A2(G288), .ZN(n751) );
  NOR2_X1 U835 ( .A1(G1971), .A2(G303), .ZN(n744) );
  NOR2_X1 U836 ( .A1(n751), .A2(n744), .ZN(n980) );
  OR2_X1 U837 ( .A1(n745), .A2(n980), .ZN(n746) );
  OR2_X1 U838 ( .A1(n762), .A2(n746), .ZN(n748) );
  INV_X1 U839 ( .A(KEYINPUT33), .ZN(n747) );
  AND2_X1 U840 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U841 ( .A1(n750), .A2(n749), .ZN(n756) );
  NAND2_X1 U842 ( .A1(n751), .A2(KEYINPUT33), .ZN(n752) );
  NOR2_X1 U843 ( .A1(n762), .A2(n752), .ZN(n754) );
  XOR2_X1 U844 ( .A(G1981), .B(G305), .Z(n970) );
  INV_X1 U845 ( .A(n970), .ZN(n753) );
  NOR2_X1 U846 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U847 ( .A1(n756), .A2(n755), .ZN(n765) );
  NAND2_X1 U848 ( .A1(n758), .A2(n757), .ZN(n761) );
  NOR2_X1 U849 ( .A1(G2090), .A2(G303), .ZN(n759) );
  NAND2_X1 U850 ( .A1(G8), .A2(n759), .ZN(n760) );
  NAND2_X1 U851 ( .A1(n761), .A2(n760), .ZN(n763) );
  NAND2_X1 U852 ( .A1(n763), .A2(n762), .ZN(n764) );
  NAND2_X1 U853 ( .A1(n765), .A2(n764), .ZN(n766) );
  NOR2_X1 U854 ( .A1(n767), .A2(n766), .ZN(n800) );
  XOR2_X1 U855 ( .A(KEYINPUT95), .B(G1991), .Z(n943) );
  NAND2_X1 U856 ( .A1(G119), .A2(n876), .ZN(n769) );
  NAND2_X1 U857 ( .A1(G131), .A2(n883), .ZN(n768) );
  NAND2_X1 U858 ( .A1(n769), .A2(n768), .ZN(n772) );
  NAND2_X1 U859 ( .A1(n881), .A2(G95), .ZN(n770) );
  XOR2_X1 U860 ( .A(KEYINPUT94), .B(n770), .Z(n771) );
  NOR2_X1 U861 ( .A1(n772), .A2(n771), .ZN(n774) );
  NAND2_X1 U862 ( .A1(n877), .A2(G107), .ZN(n773) );
  NAND2_X1 U863 ( .A1(n774), .A2(n773), .ZN(n856) );
  NAND2_X1 U864 ( .A1(n943), .A2(n856), .ZN(n784) );
  NAND2_X1 U865 ( .A1(n881), .A2(G105), .ZN(n775) );
  XNOR2_X1 U866 ( .A(n775), .B(KEYINPUT38), .ZN(n782) );
  NAND2_X1 U867 ( .A1(G129), .A2(n876), .ZN(n777) );
  NAND2_X1 U868 ( .A1(G117), .A2(n877), .ZN(n776) );
  NAND2_X1 U869 ( .A1(n777), .A2(n776), .ZN(n780) );
  NAND2_X1 U870 ( .A1(G141), .A2(n883), .ZN(n778) );
  XOR2_X1 U871 ( .A(KEYINPUT96), .B(n778), .Z(n779) );
  NOR2_X1 U872 ( .A1(n780), .A2(n779), .ZN(n781) );
  NAND2_X1 U873 ( .A1(n782), .A2(n781), .ZN(n872) );
  NAND2_X1 U874 ( .A1(G1996), .A2(n872), .ZN(n783) );
  NAND2_X1 U875 ( .A1(n784), .A2(n783), .ZN(n1000) );
  NAND2_X1 U876 ( .A1(n1000), .A2(n814), .ZN(n785) );
  XNOR2_X1 U877 ( .A(n785), .B(KEYINPUT97), .ZN(n805) );
  INV_X1 U878 ( .A(n805), .ZN(n798) );
  XNOR2_X1 U879 ( .A(KEYINPUT37), .B(G2067), .ZN(n811) );
  XNOR2_X1 U880 ( .A(KEYINPUT93), .B(KEYINPUT35), .ZN(n790) );
  NAND2_X1 U881 ( .A1(n876), .A2(G128), .ZN(n786) );
  XNOR2_X1 U882 ( .A(n786), .B(KEYINPUT92), .ZN(n788) );
  NAND2_X1 U883 ( .A1(G116), .A2(n877), .ZN(n787) );
  NAND2_X1 U884 ( .A1(n788), .A2(n787), .ZN(n789) );
  XNOR2_X1 U885 ( .A(n790), .B(n789), .ZN(n796) );
  NAND2_X1 U886 ( .A1(G104), .A2(n881), .ZN(n792) );
  NAND2_X1 U887 ( .A1(G140), .A2(n883), .ZN(n791) );
  NAND2_X1 U888 ( .A1(n792), .A2(n791), .ZN(n793) );
  XOR2_X1 U889 ( .A(KEYINPUT34), .B(n793), .Z(n794) );
  XNOR2_X1 U890 ( .A(KEYINPUT91), .B(n794), .ZN(n795) );
  NOR2_X1 U891 ( .A1(n796), .A2(n795), .ZN(n797) );
  XNOR2_X1 U892 ( .A(KEYINPUT36), .B(n797), .ZN(n875) );
  NOR2_X1 U893 ( .A1(n811), .A2(n875), .ZN(n994) );
  NAND2_X1 U894 ( .A1(n814), .A2(n994), .ZN(n809) );
  NAND2_X1 U895 ( .A1(n798), .A2(n809), .ZN(n799) );
  NOR2_X1 U896 ( .A1(n800), .A2(n799), .ZN(n801) );
  NAND2_X1 U897 ( .A1(n802), .A2(n801), .ZN(n818) );
  NOR2_X1 U898 ( .A1(G1996), .A2(n872), .ZN(n991) );
  NOR2_X1 U899 ( .A1(G1986), .A2(G290), .ZN(n803) );
  NOR2_X1 U900 ( .A1(n943), .A2(n856), .ZN(n996) );
  NOR2_X1 U901 ( .A1(n803), .A2(n996), .ZN(n804) );
  NOR2_X1 U902 ( .A1(n805), .A2(n804), .ZN(n806) );
  NOR2_X1 U903 ( .A1(n991), .A2(n806), .ZN(n807) );
  XOR2_X1 U904 ( .A(n807), .B(KEYINPUT39), .Z(n808) );
  XNOR2_X1 U905 ( .A(KEYINPUT103), .B(n808), .ZN(n810) );
  NAND2_X1 U906 ( .A1(n810), .A2(n809), .ZN(n813) );
  NAND2_X1 U907 ( .A1(n875), .A2(n811), .ZN(n812) );
  XNOR2_X1 U908 ( .A(n812), .B(KEYINPUT104), .ZN(n1009) );
  NAND2_X1 U909 ( .A1(n813), .A2(n1009), .ZN(n815) );
  NAND2_X1 U910 ( .A1(n815), .A2(n814), .ZN(n816) );
  XOR2_X1 U911 ( .A(KEYINPUT105), .B(n816), .Z(n817) );
  NAND2_X1 U912 ( .A1(n818), .A2(n817), .ZN(n819) );
  XNOR2_X1 U913 ( .A(n820), .B(n819), .ZN(G329) );
  NAND2_X1 U914 ( .A1(G2106), .A2(n821), .ZN(G217) );
  NAND2_X1 U915 ( .A1(G15), .A2(G2), .ZN(n822) );
  XNOR2_X1 U916 ( .A(KEYINPUT109), .B(n822), .ZN(n823) );
  NAND2_X1 U917 ( .A1(n823), .A2(G661), .ZN(G259) );
  NAND2_X1 U918 ( .A1(G3), .A2(G1), .ZN(n824) );
  NAND2_X1 U919 ( .A1(n825), .A2(n824), .ZN(G188) );
  XNOR2_X1 U920 ( .A(G108), .B(KEYINPUT121), .ZN(G238) );
  INV_X1 U922 ( .A(G120), .ZN(G236) );
  INV_X1 U923 ( .A(G96), .ZN(G221) );
  NOR2_X1 U924 ( .A1(n827), .A2(n826), .ZN(G325) );
  INV_X1 U925 ( .A(G325), .ZN(G261) );
  XOR2_X1 U926 ( .A(KEYINPUT112), .B(G2678), .Z(n829) );
  XNOR2_X1 U927 ( .A(KEYINPUT43), .B(G2096), .ZN(n828) );
  XNOR2_X1 U928 ( .A(n829), .B(n828), .ZN(n830) );
  XOR2_X1 U929 ( .A(n830), .B(KEYINPUT42), .Z(n832) );
  XNOR2_X1 U930 ( .A(G2067), .B(G2078), .ZN(n831) );
  XNOR2_X1 U931 ( .A(n832), .B(n831), .ZN(n836) );
  XOR2_X1 U932 ( .A(G2100), .B(G2090), .Z(n834) );
  XNOR2_X1 U933 ( .A(G2084), .B(G2072), .ZN(n833) );
  XNOR2_X1 U934 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U935 ( .A(n836), .B(n835), .Z(n838) );
  XNOR2_X1 U936 ( .A(KEYINPUT110), .B(KEYINPUT111), .ZN(n837) );
  XNOR2_X1 U937 ( .A(n838), .B(n837), .ZN(G227) );
  XOR2_X1 U938 ( .A(G1986), .B(G1976), .Z(n840) );
  XNOR2_X1 U939 ( .A(G1956), .B(G1971), .ZN(n839) );
  XNOR2_X1 U940 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U941 ( .A(G1981), .B(G1966), .Z(n842) );
  XNOR2_X1 U942 ( .A(G1996), .B(G1991), .ZN(n841) );
  XNOR2_X1 U943 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U944 ( .A(n844), .B(n843), .Z(n846) );
  XNOR2_X1 U945 ( .A(KEYINPUT113), .B(G2474), .ZN(n845) );
  XNOR2_X1 U946 ( .A(n846), .B(n845), .ZN(n848) );
  XOR2_X1 U947 ( .A(G1961), .B(KEYINPUT41), .Z(n847) );
  XNOR2_X1 U948 ( .A(n848), .B(n847), .ZN(G229) );
  NAND2_X1 U949 ( .A1(n876), .A2(G124), .ZN(n849) );
  XNOR2_X1 U950 ( .A(n849), .B(KEYINPUT44), .ZN(n851) );
  NAND2_X1 U951 ( .A1(G112), .A2(n877), .ZN(n850) );
  NAND2_X1 U952 ( .A1(n851), .A2(n850), .ZN(n855) );
  NAND2_X1 U953 ( .A1(G100), .A2(n881), .ZN(n853) );
  NAND2_X1 U954 ( .A1(G136), .A2(n883), .ZN(n852) );
  NAND2_X1 U955 ( .A1(n853), .A2(n852), .ZN(n854) );
  NOR2_X1 U956 ( .A1(n855), .A2(n854), .ZN(G162) );
  XNOR2_X1 U957 ( .A(G162), .B(n856), .ZN(n857) );
  XNOR2_X1 U958 ( .A(n857), .B(n997), .ZN(n858) );
  XOR2_X1 U959 ( .A(n858), .B(KEYINPUT118), .Z(n860) );
  XNOR2_X1 U960 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n859) );
  XNOR2_X1 U961 ( .A(n860), .B(n859), .ZN(n871) );
  NAND2_X1 U962 ( .A1(n881), .A2(G106), .ZN(n861) );
  XOR2_X1 U963 ( .A(KEYINPUT115), .B(n861), .Z(n863) );
  NAND2_X1 U964 ( .A1(n883), .A2(G142), .ZN(n862) );
  NAND2_X1 U965 ( .A1(n863), .A2(n862), .ZN(n864) );
  XNOR2_X1 U966 ( .A(n864), .B(KEYINPUT45), .ZN(n866) );
  NAND2_X1 U967 ( .A1(G118), .A2(n877), .ZN(n865) );
  NAND2_X1 U968 ( .A1(n866), .A2(n865), .ZN(n869) );
  NAND2_X1 U969 ( .A1(n876), .A2(G130), .ZN(n867) );
  XOR2_X1 U970 ( .A(KEYINPUT114), .B(n867), .Z(n868) );
  NOR2_X1 U971 ( .A1(n869), .A2(n868), .ZN(n870) );
  XNOR2_X1 U972 ( .A(n871), .B(n870), .ZN(n874) );
  XNOR2_X1 U973 ( .A(n872), .B(G164), .ZN(n873) );
  XNOR2_X1 U974 ( .A(n874), .B(n873), .ZN(n891) );
  XNOR2_X1 U975 ( .A(G160), .B(n875), .ZN(n889) );
  NAND2_X1 U976 ( .A1(G127), .A2(n876), .ZN(n879) );
  NAND2_X1 U977 ( .A1(G115), .A2(n877), .ZN(n878) );
  NAND2_X1 U978 ( .A1(n879), .A2(n878), .ZN(n880) );
  XNOR2_X1 U979 ( .A(KEYINPUT47), .B(n880), .ZN(n888) );
  NAND2_X1 U980 ( .A1(G103), .A2(n881), .ZN(n882) );
  XOR2_X1 U981 ( .A(KEYINPUT116), .B(n882), .Z(n886) );
  NAND2_X1 U982 ( .A1(G139), .A2(n883), .ZN(n884) );
  XNOR2_X1 U983 ( .A(KEYINPUT117), .B(n884), .ZN(n885) );
  NOR2_X1 U984 ( .A1(n886), .A2(n885), .ZN(n887) );
  NAND2_X1 U985 ( .A1(n888), .A2(n887), .ZN(n1003) );
  XNOR2_X1 U986 ( .A(n889), .B(n1003), .ZN(n890) );
  XOR2_X1 U987 ( .A(n891), .B(n890), .Z(n892) );
  NOR2_X1 U988 ( .A1(G37), .A2(n892), .ZN(n893) );
  XOR2_X1 U989 ( .A(KEYINPUT119), .B(n893), .Z(G395) );
  INV_X1 U990 ( .A(G301), .ZN(G171) );
  XNOR2_X1 U991 ( .A(n963), .B(G286), .ZN(n895) );
  XNOR2_X1 U992 ( .A(n895), .B(n894), .ZN(n896) );
  XNOR2_X1 U993 ( .A(n896), .B(G171), .ZN(n897) );
  NOR2_X1 U994 ( .A1(G37), .A2(n897), .ZN(n898) );
  XNOR2_X1 U995 ( .A(KEYINPUT120), .B(n898), .ZN(G397) );
  XNOR2_X1 U996 ( .A(G2443), .B(G2427), .ZN(n908) );
  XOR2_X1 U997 ( .A(G2430), .B(KEYINPUT108), .Z(n900) );
  XNOR2_X1 U998 ( .A(G2454), .B(G2435), .ZN(n899) );
  XNOR2_X1 U999 ( .A(n900), .B(n899), .ZN(n904) );
  XOR2_X1 U1000 ( .A(G2438), .B(KEYINPUT107), .Z(n902) );
  XNOR2_X1 U1001 ( .A(G1348), .B(G1341), .ZN(n901) );
  XNOR2_X1 U1002 ( .A(n902), .B(n901), .ZN(n903) );
  XOR2_X1 U1003 ( .A(n904), .B(n903), .Z(n906) );
  XNOR2_X1 U1004 ( .A(G2451), .B(G2446), .ZN(n905) );
  XNOR2_X1 U1005 ( .A(n906), .B(n905), .ZN(n907) );
  XNOR2_X1 U1006 ( .A(n908), .B(n907), .ZN(n909) );
  NAND2_X1 U1007 ( .A1(n909), .A2(G14), .ZN(n915) );
  NAND2_X1 U1008 ( .A1(G319), .A2(n915), .ZN(n912) );
  NOR2_X1 U1009 ( .A1(G227), .A2(G229), .ZN(n910) );
  XNOR2_X1 U1010 ( .A(KEYINPUT49), .B(n910), .ZN(n911) );
  NOR2_X1 U1011 ( .A1(n912), .A2(n911), .ZN(n914) );
  NOR2_X1 U1012 ( .A1(G395), .A2(G397), .ZN(n913) );
  NAND2_X1 U1013 ( .A1(n914), .A2(n913), .ZN(G225) );
  INV_X1 U1014 ( .A(G225), .ZN(G308) );
  INV_X1 U1015 ( .A(G69), .ZN(G235) );
  INV_X1 U1016 ( .A(n915), .ZN(G401) );
  XNOR2_X1 U1017 ( .A(G20), .B(n916), .ZN(n920) );
  XNOR2_X1 U1018 ( .A(G1341), .B(G19), .ZN(n918) );
  XNOR2_X1 U1019 ( .A(G1981), .B(G6), .ZN(n917) );
  NOR2_X1 U1020 ( .A1(n918), .A2(n917), .ZN(n919) );
  NAND2_X1 U1021 ( .A1(n920), .A2(n919), .ZN(n923) );
  XOR2_X1 U1022 ( .A(KEYINPUT59), .B(G1348), .Z(n921) );
  XNOR2_X1 U1023 ( .A(G4), .B(n921), .ZN(n922) );
  NOR2_X1 U1024 ( .A1(n923), .A2(n922), .ZN(n924) );
  XNOR2_X1 U1025 ( .A(KEYINPUT60), .B(n924), .ZN(n925) );
  XNOR2_X1 U1026 ( .A(n925), .B(KEYINPUT126), .ZN(n929) );
  XNOR2_X1 U1027 ( .A(G1966), .B(G21), .ZN(n927) );
  XNOR2_X1 U1028 ( .A(G1961), .B(G5), .ZN(n926) );
  NOR2_X1 U1029 ( .A1(n927), .A2(n926), .ZN(n928) );
  NAND2_X1 U1030 ( .A1(n929), .A2(n928), .ZN(n936) );
  XNOR2_X1 U1031 ( .A(G1971), .B(G22), .ZN(n931) );
  XNOR2_X1 U1032 ( .A(G23), .B(G1976), .ZN(n930) );
  NOR2_X1 U1033 ( .A1(n931), .A2(n930), .ZN(n933) );
  XOR2_X1 U1034 ( .A(G1986), .B(G24), .Z(n932) );
  NAND2_X1 U1035 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1036 ( .A(KEYINPUT58), .B(n934), .ZN(n935) );
  NOR2_X1 U1037 ( .A1(n936), .A2(n935), .ZN(n937) );
  XOR2_X1 U1038 ( .A(KEYINPUT61), .B(n937), .Z(n938) );
  NOR2_X1 U1039 ( .A1(G16), .A2(n938), .ZN(n962) );
  XNOR2_X1 U1040 ( .A(KEYINPUT125), .B(G29), .ZN(n959) );
  XOR2_X1 U1041 ( .A(KEYINPUT55), .B(KEYINPUT124), .Z(n1014) );
  XNOR2_X1 U1042 ( .A(G32), .B(n939), .ZN(n940) );
  NAND2_X1 U1043 ( .A1(n940), .A2(G28), .ZN(n950) );
  XNOR2_X1 U1044 ( .A(G2067), .B(G26), .ZN(n942) );
  XNOR2_X1 U1045 ( .A(G33), .B(G2072), .ZN(n941) );
  NOR2_X1 U1046 ( .A1(n942), .A2(n941), .ZN(n948) );
  XNOR2_X1 U1047 ( .A(n943), .B(G25), .ZN(n946) );
  XNOR2_X1 U1048 ( .A(G27), .B(n944), .ZN(n945) );
  NOR2_X1 U1049 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1050 ( .A1(n948), .A2(n947), .ZN(n949) );
  NOR2_X1 U1051 ( .A1(n950), .A2(n949), .ZN(n951) );
  XOR2_X1 U1052 ( .A(KEYINPUT53), .B(n951), .Z(n954) );
  XOR2_X1 U1053 ( .A(KEYINPUT54), .B(G34), .Z(n952) );
  XNOR2_X1 U1054 ( .A(G2084), .B(n952), .ZN(n953) );
  NAND2_X1 U1055 ( .A1(n954), .A2(n953), .ZN(n956) );
  XNOR2_X1 U1056 ( .A(G35), .B(G2090), .ZN(n955) );
  NOR2_X1 U1057 ( .A1(n956), .A2(n955), .ZN(n957) );
  XOR2_X1 U1058 ( .A(n1014), .B(n957), .Z(n958) );
  NAND2_X1 U1059 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1060 ( .A1(G11), .A2(n960), .ZN(n961) );
  NOR2_X1 U1061 ( .A1(n962), .A2(n961), .ZN(n988) );
  XNOR2_X1 U1062 ( .A(KEYINPUT56), .B(G16), .ZN(n986) );
  XNOR2_X1 U1063 ( .A(G1348), .B(n963), .ZN(n965) );
  NAND2_X1 U1064 ( .A1(G1971), .A2(G303), .ZN(n964) );
  NAND2_X1 U1065 ( .A1(n965), .A2(n964), .ZN(n966) );
  NOR2_X1 U1066 ( .A1(n967), .A2(n966), .ZN(n969) );
  NAND2_X1 U1067 ( .A1(n969), .A2(n968), .ZN(n974) );
  XNOR2_X1 U1068 ( .A(G1966), .B(G168), .ZN(n971) );
  NAND2_X1 U1069 ( .A1(n971), .A2(n970), .ZN(n972) );
  XOR2_X1 U1070 ( .A(KEYINPUT57), .B(n972), .Z(n973) );
  NOR2_X1 U1071 ( .A1(n974), .A2(n973), .ZN(n984) );
  XNOR2_X1 U1072 ( .A(n975), .B(G1956), .ZN(n977) );
  XNOR2_X1 U1073 ( .A(G171), .B(G1961), .ZN(n976) );
  NAND2_X1 U1074 ( .A1(n977), .A2(n976), .ZN(n982) );
  XOR2_X1 U1075 ( .A(G1341), .B(n978), .Z(n979) );
  NAND2_X1 U1076 ( .A1(n980), .A2(n979), .ZN(n981) );
  NOR2_X1 U1077 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1078 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1079 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1080 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1081 ( .A(n989), .B(KEYINPUT127), .ZN(n1018) );
  XOR2_X1 U1082 ( .A(G2090), .B(G162), .Z(n990) );
  NOR2_X1 U1083 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1084 ( .A(n992), .B(KEYINPUT51), .ZN(n993) );
  NOR2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n1002) );
  XOR2_X1 U1086 ( .A(G2084), .B(G160), .Z(n995) );
  NOR2_X1 U1087 ( .A1(n996), .A2(n995), .ZN(n998) );
  NAND2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n999) );
  NOR2_X1 U1089 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1090 ( .A1(n1002), .A2(n1001), .ZN(n1012) );
  XNOR2_X1 U1091 ( .A(KEYINPUT122), .B(n1003), .ZN(n1004) );
  XOR2_X1 U1092 ( .A(G2072), .B(n1004), .Z(n1006) );
  XNOR2_X1 U1093 ( .A(G164), .B(G2078), .ZN(n1005) );
  NAND2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1095 ( .A(n1007), .B(KEYINPUT50), .ZN(n1008) );
  XNOR2_X1 U1096 ( .A(n1008), .B(KEYINPUT123), .ZN(n1010) );
  NAND2_X1 U1097 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NOR2_X1 U1098 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1099 ( .A(KEYINPUT52), .B(n1013), .ZN(n1015) );
  NAND2_X1 U1100 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1101 ( .A1(n1016), .A2(G29), .ZN(n1017) );
  NAND2_X1 U1102 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XOR2_X1 U1103 ( .A(KEYINPUT62), .B(n1019), .Z(G311) );
  INV_X1 U1104 ( .A(G311), .ZN(G150) );
endmodule

