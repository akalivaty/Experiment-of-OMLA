//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 1 1 0 1 0 1 1 1 1 0 0 1 0 0 1 1 0 0 1 0 1 0 0 1 1 1 0 0 0 1 0 1 0 1 0 1 0 0 0 1 0 0 1 1 0 1 0 0 1 0 0 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n724, new_n725, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n808, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n882, new_n883, new_n885,
    new_n886, new_n887, new_n888, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n943, new_n944, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n999, new_n1000;
  XOR2_X1   g000(.A(G134gat), .B(G162gat), .Z(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  AOI21_X1  g002(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT100), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT101), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT7), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(KEYINPUT101), .A2(KEYINPUT7), .ZN(new_n210));
  NAND4_X1  g009(.A1(new_n209), .A2(G85gat), .A3(G92gat), .A4(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G85gat), .ZN(new_n212));
  INV_X1    g011(.A(G92gat), .ZN(new_n213));
  OAI211_X1 g012(.A(new_n207), .B(new_n208), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(G99gat), .A2(G106gat), .ZN(new_n215));
  AOI22_X1  g014(.A1(KEYINPUT8), .A2(new_n215), .B1(new_n212), .B2(new_n213), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n211), .A2(new_n214), .A3(new_n216), .ZN(new_n217));
  XOR2_X1   g016(.A(G99gat), .B(G106gat), .Z(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT103), .ZN(new_n221));
  OAI21_X1  g020(.A(KEYINPUT102), .B1(new_n217), .B2(new_n218), .ZN(new_n222));
  INV_X1    g021(.A(new_n222), .ZN(new_n223));
  NOR3_X1   g022(.A1(new_n217), .A2(KEYINPUT102), .A3(new_n218), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n221), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  OR3_X1    g024(.A1(new_n217), .A2(KEYINPUT102), .A3(new_n218), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n226), .A2(KEYINPUT103), .A3(new_n222), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n220), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT104), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NOR3_X1   g029(.A1(new_n223), .A2(new_n221), .A3(new_n224), .ZN(new_n231));
  AOI21_X1  g030(.A(KEYINPUT103), .B1(new_n226), .B2(new_n222), .ZN(new_n232));
  OAI211_X1 g031(.A(new_n229), .B(new_n219), .C1(new_n231), .C2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  OAI21_X1  g033(.A(KEYINPUT105), .B1(new_n230), .B2(new_n234), .ZN(new_n235));
  XOR2_X1   g034(.A(G43gat), .B(G50gat), .Z(new_n236));
  INV_X1    g035(.A(KEYINPUT15), .ZN(new_n237));
  AOI22_X1  g036(.A1(new_n236), .A2(new_n237), .B1(G29gat), .B2(G36gat), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT95), .ZN(new_n239));
  OR3_X1    g038(.A1(new_n239), .A2(G29gat), .A3(G36gat), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n239), .B1(G29gat), .B2(G36gat), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n240), .A2(new_n241), .A3(KEYINPUT14), .ZN(new_n242));
  OR2_X1    g041(.A1(new_n241), .A2(KEYINPUT14), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n238), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n236), .A2(new_n237), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n245), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n247), .A2(new_n238), .A3(new_n242), .A4(new_n243), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT17), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n246), .A2(KEYINPUT17), .A3(new_n248), .ZN(new_n252));
  AND2_X1   g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n219), .B1(new_n231), .B2(new_n232), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(KEYINPUT104), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT105), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n255), .A2(new_n256), .A3(new_n233), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n235), .A2(new_n253), .A3(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n255), .A2(new_n249), .A3(new_n233), .ZN(new_n259));
  NAND3_X1  g058(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n260));
  AND2_X1   g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(G190gat), .ZN(new_n263));
  INV_X1    g062(.A(G190gat), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n258), .A2(new_n261), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(G218gat), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n206), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n263), .A2(G218gat), .A3(new_n265), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n205), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  AND3_X1   g069(.A1(new_n258), .A2(new_n261), .A3(new_n264), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n264), .B1(new_n258), .B2(new_n261), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n267), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n273), .A2(new_n269), .A3(KEYINPUT100), .A4(new_n205), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n203), .B1(new_n270), .B2(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(G57gat), .B(G64gat), .ZN(new_n277));
  AOI21_X1  g076(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n278));
  OR2_X1    g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(G71gat), .B(G78gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n279), .B(new_n280), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n281), .A2(KEYINPUT21), .ZN(new_n282));
  XNOR2_X1  g081(.A(G127gat), .B(G155gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n282), .B(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(G15gat), .B(G22gat), .ZN(new_n285));
  INV_X1    g084(.A(G1gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(KEYINPUT16), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n288), .B1(G1gat), .B2(new_n285), .ZN(new_n289));
  OR2_X1    g088(.A1(new_n289), .A2(G8gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(G8gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n292), .B1(KEYINPUT21), .B2(new_n281), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n284), .B(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(G231gat), .A2(G233gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n295), .B(KEYINPUT99), .ZN(new_n296));
  XOR2_X1   g095(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n297));
  XNOR2_X1  g096(.A(new_n296), .B(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(G183gat), .B(G211gat), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n298), .B(new_n299), .ZN(new_n300));
  XOR2_X1   g099(.A(new_n294), .B(new_n300), .Z(new_n301));
  NAND3_X1  g100(.A1(new_n273), .A2(new_n269), .A3(KEYINPUT100), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(new_n204), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n303), .A2(new_n202), .A3(new_n274), .ZN(new_n304));
  NAND2_X1  g103(.A1(G230gat), .A2(G233gat), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n255), .A2(KEYINPUT10), .A3(new_n281), .A4(new_n233), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT10), .ZN(new_n308));
  OR2_X1    g107(.A1(new_n217), .A2(KEYINPUT106), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n217), .A2(KEYINPUT106), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n309), .A2(new_n218), .A3(new_n310), .ZN(new_n311));
  OAI211_X1 g110(.A(new_n311), .B(new_n281), .C1(new_n223), .C2(new_n224), .ZN(new_n312));
  OAI211_X1 g111(.A(new_n308), .B(new_n312), .C1(new_n228), .C2(new_n281), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n306), .B1(new_n307), .B2(new_n313), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n312), .B1(new_n228), .B2(new_n281), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n314), .B1(new_n306), .B2(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(G120gat), .B(G148gat), .ZN(new_n317));
  XNOR2_X1  g116(.A(G176gat), .B(G204gat), .ZN(new_n318));
  XOR2_X1   g117(.A(new_n317), .B(new_n318), .Z(new_n319));
  OR2_X1    g118(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n316), .A2(new_n319), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  NAND4_X1  g122(.A1(new_n276), .A2(new_n301), .A3(new_n304), .A4(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT96), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n292), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n290), .A2(KEYINPUT96), .A3(new_n291), .ZN(new_n327));
  NAND4_X1  g126(.A1(new_n251), .A2(new_n252), .A3(new_n326), .A4(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n249), .A2(new_n292), .ZN(new_n329));
  NAND2_X1  g128(.A1(G229gat), .A2(G233gat), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n328), .A2(KEYINPUT18), .A3(new_n329), .A4(new_n330), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n249), .B(new_n292), .ZN(new_n332));
  XOR2_X1   g131(.A(new_n330), .B(KEYINPUT13), .Z(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(G113gat), .B(G141gat), .ZN(new_n335));
  XNOR2_X1  g134(.A(KEYINPUT93), .B(KEYINPUT11), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n335), .B(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(G169gat), .B(G197gat), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n337), .B(new_n338), .ZN(new_n339));
  XOR2_X1   g138(.A(new_n339), .B(KEYINPUT12), .Z(new_n340));
  AND3_X1   g139(.A1(new_n331), .A2(new_n334), .A3(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT18), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT98), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n342), .A2(KEYINPUT98), .A3(new_n343), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n341), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n344), .A2(KEYINPUT97), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n331), .A2(new_n334), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT97), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n351), .B1(new_n342), .B2(new_n343), .ZN(new_n352));
  NOR3_X1   g151(.A1(new_n349), .A2(new_n350), .A3(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n340), .B(KEYINPUT94), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n348), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  OR2_X1    g155(.A1(new_n324), .A2(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(KEYINPUT89), .B(KEYINPUT38), .ZN(new_n358));
  XNOR2_X1  g157(.A(G8gat), .B(G36gat), .ZN(new_n359));
  XNOR2_X1  g158(.A(G64gat), .B(G92gat), .ZN(new_n360));
  XOR2_X1   g159(.A(new_n359), .B(new_n360), .Z(new_n361));
  NAND2_X1  g160(.A1(G197gat), .A2(G204gat), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  NOR2_X1   g162(.A1(G197gat), .A2(G204gat), .ZN(new_n364));
  AND2_X1   g163(.A1(G211gat), .A2(G218gat), .ZN(new_n365));
  OAI22_X1  g164(.A1(new_n363), .A2(new_n364), .B1(new_n365), .B2(KEYINPUT22), .ZN(new_n366));
  NOR2_X1   g165(.A1(G211gat), .A2(G218gat), .ZN(new_n367));
  NOR3_X1   g166(.A1(new_n365), .A2(new_n367), .A3(KEYINPUT74), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT74), .ZN(new_n369));
  INV_X1    g168(.A(G211gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(new_n267), .ZN(new_n371));
  NAND2_X1  g170(.A1(G211gat), .A2(G218gat), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n369), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n366), .B1(new_n368), .B2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(G197gat), .ZN(new_n375));
  INV_X1    g174(.A(G204gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT22), .ZN(new_n378));
  AOI22_X1  g177(.A1(new_n377), .A2(new_n362), .B1(new_n378), .B2(new_n372), .ZN(new_n379));
  OAI21_X1  g178(.A(KEYINPUT74), .B1(new_n365), .B2(new_n367), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n371), .A2(new_n369), .A3(new_n372), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n374), .A2(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(new_n383), .B(KEYINPUT75), .ZN(new_n384));
  NAND2_X1  g183(.A1(G183gat), .A2(G190gat), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT68), .ZN(new_n386));
  NOR2_X1   g185(.A1(G169gat), .A2(G176gat), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n386), .B1(new_n387), .B2(KEYINPUT66), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT26), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT66), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n390), .B1(new_n389), .B2(KEYINPUT68), .ZN(new_n391));
  AOI22_X1  g190(.A1(new_n388), .A2(new_n389), .B1(new_n387), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(G169gat), .A2(G176gat), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT64), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(KEYINPUT64), .A2(G169gat), .A3(G176gat), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n385), .B1(new_n392), .B2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT69), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  OAI211_X1 g200(.A(KEYINPUT69), .B(new_n385), .C1(new_n392), .C2(new_n398), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(KEYINPUT27), .B(G183gat), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(new_n264), .ZN(new_n405));
  XNOR2_X1  g204(.A(new_n405), .B(KEYINPUT28), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n403), .A2(new_n407), .ZN(new_n408));
  AND2_X1   g207(.A1(G226gat), .A2(G233gat), .ZN(new_n409));
  INV_X1    g208(.A(G169gat), .ZN(new_n410));
  INV_X1    g209(.A(G176gat), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n410), .A2(new_n411), .A3(KEYINPUT23), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT23), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n413), .B1(G169gat), .B2(G176gat), .ZN(new_n414));
  AND3_X1   g213(.A1(KEYINPUT64), .A2(G169gat), .A3(G176gat), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT64), .B1(G169gat), .B2(G176gat), .ZN(new_n416));
  OAI211_X1 g215(.A(new_n412), .B(new_n414), .C1(new_n415), .C2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT65), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT24), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n420), .A2(G183gat), .A3(G190gat), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  XOR2_X1   g221(.A(G183gat), .B(G190gat), .Z(new_n423));
  AOI21_X1  g222(.A(new_n422), .B1(new_n423), .B2(KEYINPUT24), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n397), .A2(KEYINPUT65), .A3(new_n414), .A4(new_n412), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n419), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT25), .ZN(new_n427));
  INV_X1    g226(.A(new_n387), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n413), .B1(new_n428), .B2(new_n390), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n429), .B1(new_n390), .B2(new_n428), .ZN(new_n430));
  XNOR2_X1  g229(.A(G183gat), .B(G190gat), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n421), .B1(new_n431), .B2(new_n420), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n414), .B(KEYINPUT25), .C1(new_n415), .C2(new_n416), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  AOI22_X1  g233(.A1(new_n426), .A2(new_n427), .B1(new_n430), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n408), .A2(new_n409), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n406), .B1(new_n401), .B2(new_n402), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n432), .B1(new_n418), .B2(new_n417), .ZN(new_n439));
  AOI21_X1  g238(.A(KEYINPUT25), .B1(new_n439), .B2(new_n425), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n434), .A2(new_n430), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  OAI21_X1  g241(.A(KEYINPUT67), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT67), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n435), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n438), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n409), .A2(KEYINPUT29), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n384), .B(new_n437), .C1(new_n446), .C2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT76), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n426), .A2(new_n427), .ZN(new_n452));
  AND3_X1   g251(.A1(new_n452), .A2(new_n444), .A3(new_n441), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n444), .B1(new_n452), .B2(new_n441), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n409), .B(new_n408), .C1(new_n453), .C2(new_n454), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n447), .B1(new_n438), .B2(new_n435), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n383), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n408), .B1(new_n453), .B2(new_n454), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(new_n447), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n461), .A2(KEYINPUT76), .A3(new_n384), .A4(new_n437), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n451), .A2(new_n459), .A3(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n361), .B1(new_n463), .B2(KEYINPUT37), .ZN(new_n464));
  XOR2_X1   g263(.A(KEYINPUT90), .B(KEYINPUT37), .Z(new_n465));
  OAI22_X1  g264(.A1(new_n464), .A2(KEYINPUT91), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT91), .ZN(new_n467));
  AOI211_X1 g266(.A(new_n467), .B(new_n361), .C1(new_n463), .C2(KEYINPUT37), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n358), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  XNOR2_X1  g268(.A(G1gat), .B(G29gat), .ZN(new_n470));
  XNOR2_X1  g269(.A(new_n470), .B(KEYINPUT0), .ZN(new_n471));
  XNOR2_X1  g270(.A(G57gat), .B(G85gat), .ZN(new_n472));
  XOR2_X1   g271(.A(new_n471), .B(new_n472), .Z(new_n473));
  XOR2_X1   g272(.A(KEYINPUT71), .B(G113gat), .Z(new_n474));
  INV_X1    g273(.A(G120gat), .ZN(new_n475));
  XNOR2_X1  g274(.A(KEYINPUT70), .B(G120gat), .ZN(new_n476));
  INV_X1    g275(.A(G113gat), .ZN(new_n477));
  OAI22_X1  g276(.A1(new_n474), .A2(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  XOR2_X1   g277(.A(G127gat), .B(G134gat), .Z(new_n479));
  NOR2_X1   g278(.A1(new_n479), .A2(KEYINPUT1), .ZN(new_n480));
  AOI21_X1  g279(.A(KEYINPUT1), .B1(new_n477), .B2(new_n475), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n481), .B1(new_n477), .B2(new_n475), .ZN(new_n482));
  AOI22_X1  g281(.A1(new_n478), .A2(new_n480), .B1(new_n479), .B2(new_n482), .ZN(new_n483));
  XNOR2_X1  g282(.A(KEYINPUT79), .B(G155gat), .ZN(new_n484));
  INV_X1    g283(.A(G162gat), .ZN(new_n485));
  OAI21_X1  g284(.A(KEYINPUT2), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(G141gat), .ZN(new_n487));
  INV_X1    g286(.A(G148gat), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n485), .A2(G155gat), .ZN(new_n490));
  INV_X1    g289(.A(G155gat), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(G162gat), .ZN(new_n492));
  NAND2_X1  g291(.A1(G141gat), .A2(G148gat), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n489), .A2(new_n490), .A3(new_n492), .A4(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT2), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n489), .A2(new_n496), .A3(new_n493), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n490), .A2(new_n492), .ZN(new_n498));
  AOI22_X1  g297(.A1(new_n486), .A2(new_n495), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT4), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n483), .A2(KEYINPUT4), .A3(new_n499), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n478), .A2(new_n480), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n482), .A2(new_n479), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n497), .A2(new_n498), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n491), .A2(KEYINPUT79), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT79), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(G155gat), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n496), .B1(new_n513), .B2(G162gat), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n509), .B1(new_n514), .B2(new_n494), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(KEYINPUT3), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT3), .ZN(new_n517));
  OAI211_X1 g316(.A(new_n517), .B(new_n509), .C1(new_n514), .C2(new_n494), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n508), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(KEYINPUT80), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT80), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n508), .A2(new_n516), .A3(new_n521), .A4(new_n518), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n505), .A2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT5), .ZN(new_n525));
  NAND2_X1  g324(.A1(G225gat), .A2(G233gat), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  NOR3_X1   g326(.A1(new_n524), .A2(new_n525), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n508), .A2(new_n515), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(new_n500), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n525), .B1(new_n530), .B2(new_n527), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n504), .B1(new_n520), .B2(new_n522), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n531), .B1(new_n532), .B2(new_n526), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n473), .B1(new_n528), .B2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT6), .ZN(new_n535));
  INV_X1    g334(.A(new_n531), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n536), .B1(new_n524), .B2(new_n527), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n532), .A2(KEYINPUT5), .A3(new_n526), .ZN(new_n538));
  INV_X1    g337(.A(new_n473), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n534), .A2(new_n535), .A3(new_n540), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n537), .A2(new_n538), .A3(KEYINPUT6), .A4(new_n539), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n451), .A2(new_n462), .A3(new_n361), .A4(new_n459), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n463), .A2(new_n465), .ZN(new_n545));
  NOR3_X1   g344(.A1(new_n545), .A2(new_n358), .A3(new_n361), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n438), .A2(new_n435), .ZN(new_n547));
  AOI22_X1  g346(.A1(new_n460), .A2(new_n447), .B1(new_n409), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g347(.A(KEYINPUT88), .B1(new_n548), .B2(new_n384), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n549), .B1(new_n458), .B2(new_n457), .ZN(new_n550));
  NOR3_X1   g349(.A1(new_n548), .A2(KEYINPUT88), .A3(new_n384), .ZN(new_n551));
  OAI21_X1  g350(.A(KEYINPUT37), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n544), .B1(new_n546), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n469), .A2(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(G78gat), .B(G106gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(KEYINPUT31), .B(G50gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n555), .B(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT75), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n383), .B(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT29), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n518), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  OAI21_X1  g362(.A(KEYINPUT83), .B1(new_n560), .B2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT83), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n384), .A2(new_n565), .A3(new_n562), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n374), .A2(new_n561), .A3(new_n382), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n499), .B1(new_n568), .B2(new_n517), .ZN(new_n569));
  NAND2_X1  g368(.A1(G228gat), .A2(G233gat), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  XOR2_X1   g371(.A(KEYINPUT84), .B(G22gat), .Z(new_n573));
  NAND2_X1  g372(.A1(new_n568), .A2(new_n517), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(new_n515), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(KEYINPUT81), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT81), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n569), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n383), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n576), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(KEYINPUT82), .B1(new_n580), .B2(new_n570), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n579), .B1(new_n569), .B2(new_n577), .ZN(new_n582));
  AOI211_X1 g381(.A(KEYINPUT81), .B(new_n499), .C1(new_n568), .C2(new_n517), .ZN(new_n583));
  OAI211_X1 g382(.A(KEYINPUT82), .B(new_n570), .C1(new_n582), .C2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  OAI211_X1 g384(.A(new_n572), .B(new_n573), .C1(new_n581), .C2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n586), .A2(KEYINPUT86), .ZN(new_n587));
  INV_X1    g386(.A(new_n571), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n588), .B1(new_n564), .B2(new_n566), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n570), .B1(new_n582), .B2(new_n583), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT82), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n589), .B1(new_n592), .B2(new_n584), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT86), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n593), .A2(new_n594), .A3(new_n573), .ZN(new_n595));
  AND2_X1   g394(.A1(new_n587), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT85), .ZN(new_n597));
  OR2_X1    g396(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n593), .A2(new_n597), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n598), .A2(G22gat), .A3(new_n599), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n558), .B1(new_n596), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n586), .A2(new_n558), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n593), .A2(new_n573), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g403(.A(KEYINPUT87), .B1(new_n601), .B2(new_n604), .ZN(new_n605));
  OAI21_X1  g404(.A(G22gat), .B1(new_n593), .B2(new_n597), .ZN(new_n606));
  AOI211_X1 g405(.A(KEYINPUT85), .B(new_n589), .C1(new_n592), .C2(new_n584), .ZN(new_n607));
  OAI211_X1 g406(.A(new_n595), .B(new_n587), .C1(new_n606), .C2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(new_n557), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT87), .ZN(new_n610));
  INV_X1    g409(.A(new_n604), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n361), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n463), .A2(new_n613), .ZN(new_n614));
  AND2_X1   g413(.A1(new_n462), .A2(new_n459), .ZN(new_n615));
  NAND4_X1  g414(.A1(new_n615), .A2(KEYINPUT30), .A3(new_n361), .A4(new_n451), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT30), .ZN(new_n617));
  AND3_X1   g416(.A1(new_n543), .A2(KEYINPUT78), .A3(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(KEYINPUT78), .B1(new_n543), .B2(new_n617), .ZN(new_n619));
  OAI211_X1 g418(.A(new_n614), .B(new_n616), .C1(new_n618), .C2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n524), .A2(new_n527), .ZN(new_n621));
  OR2_X1    g420(.A1(new_n621), .A2(KEYINPUT39), .ZN(new_n622));
  OAI211_X1 g421(.A(new_n621), .B(KEYINPUT39), .C1(new_n527), .C2(new_n530), .ZN(new_n623));
  NAND4_X1  g422(.A1(new_n622), .A2(new_n623), .A3(KEYINPUT40), .A4(new_n473), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n622), .A2(new_n623), .A3(new_n473), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT40), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AND2_X1   g426(.A1(new_n627), .A2(new_n540), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n620), .A2(new_n624), .A3(new_n628), .ZN(new_n629));
  NAND4_X1  g428(.A1(new_n554), .A2(new_n605), .A3(new_n612), .A4(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT77), .ZN(new_n631));
  AND3_X1   g430(.A1(new_n616), .A2(new_n631), .A3(new_n614), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n631), .B1(new_n616), .B2(new_n614), .ZN(new_n633));
  OR2_X1    g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n541), .A2(new_n542), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n635), .B1(new_n618), .B2(new_n619), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n610), .B1(new_n609), .B2(new_n611), .ZN(new_n637));
  AOI211_X1 g436(.A(KEYINPUT87), .B(new_n604), .C1(new_n608), .C2(new_n557), .ZN(new_n638));
  OAI22_X1  g437(.A1(new_n634), .A2(new_n636), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT36), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT34), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n460), .A2(new_n483), .ZN(new_n642));
  OAI211_X1 g441(.A(new_n508), .B(new_n408), .C1(new_n453), .C2(new_n454), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(G227gat), .ZN(new_n645));
  INV_X1    g444(.A(G233gat), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n641), .B1(new_n644), .B2(new_n648), .ZN(new_n649));
  AOI211_X1 g448(.A(KEYINPUT34), .B(new_n647), .C1(new_n642), .C2(new_n643), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n642), .A2(new_n647), .A3(new_n643), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(KEYINPUT32), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT33), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g454(.A(G15gat), .B(G43gat), .Z(new_n656));
  XNOR2_X1  g455(.A(G71gat), .B(G99gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n653), .A2(new_n655), .A3(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n658), .ZN(new_n660));
  OAI211_X1 g459(.A(new_n652), .B(KEYINPUT32), .C1(new_n654), .C2(new_n660), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n651), .A2(new_n659), .A3(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT73), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND4_X1  g463(.A1(new_n651), .A2(new_n659), .A3(KEYINPUT73), .A4(new_n661), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n659), .A2(new_n661), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT72), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n651), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n659), .A2(KEYINPUT72), .A3(new_n661), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n640), .B1(new_n666), .B2(new_n672), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n651), .B1(new_n659), .B2(new_n661), .ZN(new_n674));
  AOI211_X1 g473(.A(KEYINPUT36), .B(new_n674), .C1(new_n664), .C2(new_n665), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  AND3_X1   g475(.A1(new_n630), .A2(new_n639), .A3(new_n676), .ZN(new_n677));
  NOR3_X1   g476(.A1(new_n636), .A2(new_n632), .A3(new_n633), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n651), .B1(new_n667), .B2(new_n668), .ZN(new_n679));
  AOI22_X1  g478(.A1(new_n671), .A2(new_n679), .B1(new_n664), .B2(new_n665), .ZN(new_n680));
  NAND4_X1  g479(.A1(new_n678), .A2(new_n680), .A3(new_n605), .A4(new_n612), .ZN(new_n681));
  NOR3_X1   g480(.A1(new_n637), .A2(new_n638), .A3(new_n620), .ZN(new_n682));
  INV_X1    g481(.A(new_n674), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n666), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n635), .ZN(new_n685));
  OR2_X1    g484(.A1(new_n685), .A2(KEYINPUT35), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  AOI22_X1  g486(.A1(KEYINPUT35), .A2(new_n681), .B1(new_n682), .B2(new_n687), .ZN(new_n688));
  OAI21_X1  g487(.A(KEYINPUT92), .B1(new_n677), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n681), .A2(KEYINPUT35), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n682), .A2(new_n687), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n630), .A2(new_n676), .A3(new_n639), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT92), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n692), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n357), .B1(new_n689), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(new_n685), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g497(.A(KEYINPUT16), .B(G8gat), .Z(new_n699));
  NAND4_X1  g498(.A1(new_n696), .A2(KEYINPUT42), .A3(new_n620), .A4(new_n699), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(KEYINPUT110), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n696), .A2(new_n620), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT108), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n696), .A2(KEYINPUT108), .A3(new_n620), .ZN(new_n705));
  AND3_X1   g504(.A1(new_n704), .A2(G8gat), .A3(new_n705), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n701), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n704), .A2(new_n705), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(new_n699), .ZN(new_n709));
  XOR2_X1   g508(.A(KEYINPUT107), .B(KEYINPUT42), .Z(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  AOI21_X1  g510(.A(KEYINPUT109), .B1(new_n709), .B2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n699), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n713), .B1(new_n704), .B2(new_n705), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT109), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n714), .A2(new_n715), .A3(new_n710), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n707), .B1(new_n712), .B2(new_n716), .ZN(G1325gat));
  INV_X1    g516(.A(new_n696), .ZN(new_n718));
  OR3_X1    g517(.A1(new_n718), .A2(G15gat), .A3(new_n684), .ZN(new_n719));
  OAI21_X1  g518(.A(G15gat), .B1(new_n718), .B2(new_n676), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(G1326gat));
  NOR2_X1   g520(.A1(new_n637), .A2(new_n638), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n696), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g523(.A(KEYINPUT43), .B(G22gat), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n724), .B(new_n725), .ZN(G1327gat));
  NOR3_X1   g525(.A1(new_n322), .A2(new_n356), .A3(new_n301), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT44), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n689), .A2(new_n695), .ZN(new_n729));
  AND3_X1   g528(.A1(new_n303), .A2(new_n202), .A3(new_n274), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n202), .B1(new_n303), .B2(new_n274), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n728), .B1(new_n729), .B2(new_n733), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n732), .B1(new_n692), .B2(new_n693), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(new_n728), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  OAI211_X1 g536(.A(new_n685), .B(new_n727), .C1(new_n734), .C2(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(G29gat), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT45), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n729), .A2(new_n733), .A3(new_n727), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n635), .A2(G29gat), .ZN(new_n742));
  INV_X1    g541(.A(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n740), .B1(new_n741), .B2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(new_n741), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n745), .A2(KEYINPUT45), .A3(new_n742), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n739), .A2(new_n744), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(KEYINPUT111), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT111), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n739), .A2(new_n749), .A3(new_n744), .A4(new_n746), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n748), .A2(new_n750), .ZN(G1328gat));
  NAND2_X1  g550(.A1(new_n729), .A2(new_n733), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(KEYINPUT44), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(new_n736), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(new_n727), .ZN(new_n755));
  INV_X1    g554(.A(new_n620), .ZN(new_n756));
  OAI21_X1  g555(.A(G36gat), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n756), .A2(G36gat), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  OAI21_X1  g558(.A(KEYINPUT46), .B1(new_n741), .B2(new_n759), .ZN(new_n760));
  OR3_X1    g559(.A1(new_n741), .A2(KEYINPUT46), .A3(new_n759), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n757), .A2(new_n760), .A3(new_n761), .ZN(G1329gat));
  NOR2_X1   g561(.A1(new_n684), .A2(G43gat), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  OR3_X1    g563(.A1(new_n741), .A2(KEYINPUT112), .A3(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(KEYINPUT112), .B1(new_n741), .B2(new_n764), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(new_n676), .ZN(new_n768));
  OAI211_X1 g567(.A(new_n768), .B(new_n727), .C1(new_n734), .C2(new_n737), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(G43gat), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n767), .A2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT47), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n767), .A2(new_n770), .A3(KEYINPUT47), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(G1330gat));
  INV_X1    g574(.A(G50gat), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n776), .B1(new_n741), .B2(new_n722), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n722), .A2(new_n776), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n777), .B1(new_n755), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(KEYINPUT48), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT48), .ZN(new_n782));
  OAI211_X1 g581(.A(new_n782), .B(new_n777), .C1(new_n755), .C2(new_n779), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n781), .A2(new_n783), .ZN(G1331gat));
  NOR2_X1   g583(.A1(new_n677), .A2(new_n688), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n732), .A2(new_n356), .A3(new_n301), .A4(new_n322), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  OR2_X1    g586(.A1(new_n787), .A2(KEYINPUT113), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(KEYINPUT113), .ZN(new_n789));
  AND2_X1   g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  XOR2_X1   g589(.A(new_n635), .B(KEYINPUT114), .Z(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n792), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g592(.A1(new_n788), .A2(new_n789), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n794), .A2(new_n756), .ZN(new_n795));
  NOR2_X1   g594(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n796));
  AND2_X1   g595(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n795), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n798), .B1(new_n795), .B2(new_n796), .ZN(G1333gat));
  NOR2_X1   g598(.A1(new_n684), .A2(G71gat), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n790), .A2(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(G71gat), .B1(new_n794), .B2(new_n676), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT50), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n801), .A2(new_n802), .A3(KEYINPUT50), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(G1334gat));
  NAND2_X1  g606(.A1(new_n790), .A2(new_n723), .ZN(new_n808));
  XNOR2_X1  g607(.A(new_n808), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g608(.A1(new_n355), .A2(new_n301), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n810), .A2(new_n322), .ZN(new_n811));
  OAI211_X1 g610(.A(new_n685), .B(new_n811), .C1(new_n734), .C2(new_n737), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n212), .B1(new_n812), .B2(KEYINPUT115), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n813), .B1(KEYINPUT115), .B2(new_n812), .ZN(new_n814));
  AND3_X1   g613(.A1(new_n735), .A2(KEYINPUT51), .A3(new_n810), .ZN(new_n815));
  AOI21_X1  g614(.A(KEYINPUT51), .B1(new_n735), .B2(new_n810), .ZN(new_n816));
  OR2_X1    g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(new_n322), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n685), .A2(new_n212), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n814), .B1(new_n818), .B2(new_n819), .ZN(G1336gat));
  NOR2_X1   g619(.A1(new_n756), .A2(new_n213), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n754), .A2(new_n811), .A3(new_n821), .ZN(new_n822));
  OAI211_X1 g621(.A(new_n620), .B(new_n322), .C1(new_n815), .C2(new_n816), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT52), .ZN(new_n824));
  AOI22_X1  g623(.A1(new_n823), .A2(new_n213), .B1(KEYINPUT116), .B2(new_n824), .ZN(new_n825));
  OR2_X1    g624(.A1(new_n824), .A2(KEYINPUT116), .ZN(new_n826));
  AND3_X1   g625(.A1(new_n822), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n826), .B1(new_n822), .B2(new_n825), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n827), .A2(new_n828), .ZN(G1337gat));
  NAND3_X1  g628(.A1(new_n754), .A2(new_n768), .A3(new_n811), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(G99gat), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n684), .A2(new_n323), .A3(G99gat), .ZN(new_n832));
  XNOR2_X1  g631(.A(new_n832), .B(KEYINPUT117), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n831), .A2(new_n834), .ZN(G1338gat));
  OAI211_X1 g634(.A(new_n723), .B(new_n811), .C1(new_n734), .C2(new_n737), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(G106gat), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(KEYINPUT118), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n722), .A2(G106gat), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n817), .A2(new_n322), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n838), .A2(new_n841), .A3(KEYINPUT53), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT53), .ZN(new_n843));
  OAI211_X1 g642(.A(new_n837), .B(new_n840), .C1(KEYINPUT118), .C2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n842), .A2(new_n844), .ZN(G1339gat));
  INV_X1    g644(.A(new_n301), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n307), .A2(new_n313), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n305), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n307), .A2(new_n306), .A3(new_n313), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n848), .A2(new_n849), .A3(KEYINPUT54), .ZN(new_n850));
  XNOR2_X1  g649(.A(KEYINPUT119), .B(KEYINPUT54), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n319), .B1(new_n314), .B2(new_n851), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n850), .A2(KEYINPUT55), .A3(new_n852), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n355), .A2(new_n853), .A3(new_n321), .ZN(new_n854));
  AOI21_X1  g653(.A(KEYINPUT55), .B1(new_n850), .B2(new_n852), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(new_n339), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n330), .B1(new_n328), .B2(new_n329), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n332), .A2(new_n333), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n857), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n348), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n861), .B1(new_n320), .B2(new_n321), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n856), .A2(new_n862), .ZN(new_n863));
  NOR3_X1   g662(.A1(new_n730), .A2(new_n731), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n853), .A2(new_n321), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n865), .A2(new_n861), .A3(new_n855), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n867), .B1(new_n276), .B2(new_n304), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n846), .B1(new_n864), .B2(new_n868), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n732), .A2(new_n356), .A3(new_n301), .A4(new_n323), .ZN(new_n870));
  AOI211_X1 g669(.A(new_n723), .B(new_n684), .C1(new_n869), .C2(new_n870), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n620), .A2(new_n635), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g672(.A(G113gat), .B1(new_n873), .B2(new_n356), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n869), .A2(new_n870), .ZN(new_n875));
  NAND4_X1  g674(.A1(new_n875), .A2(new_n680), .A3(new_n682), .A4(new_n791), .ZN(new_n876));
  OR2_X1    g675(.A1(new_n356), .A2(new_n474), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n874), .B1(new_n876), .B2(new_n877), .ZN(G1340gat));
  OAI21_X1  g677(.A(G120gat), .B1(new_n873), .B2(new_n323), .ZN(new_n879));
  OR2_X1    g678(.A1(new_n323), .A2(new_n476), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n879), .B1(new_n876), .B2(new_n880), .ZN(G1341gat));
  OAI21_X1  g680(.A(G127gat), .B1(new_n873), .B2(new_n846), .ZN(new_n882));
  OR2_X1    g681(.A1(new_n846), .A2(G127gat), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n882), .B1(new_n876), .B2(new_n883), .ZN(G1342gat));
  OR3_X1    g683(.A1(new_n876), .A2(G134gat), .A3(new_n732), .ZN(new_n885));
  OR2_X1    g684(.A1(new_n885), .A2(KEYINPUT56), .ZN(new_n886));
  OAI21_X1  g685(.A(G134gat), .B1(new_n873), .B2(new_n732), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n885), .A2(KEYINPUT56), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(G1343gat));
  NOR3_X1   g688(.A1(new_n768), .A2(new_n722), .A3(new_n620), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n875), .A2(new_n791), .A3(new_n890), .ZN(new_n891));
  NOR3_X1   g690(.A1(new_n891), .A2(G141gat), .A3(new_n356), .ZN(new_n892));
  INV_X1    g691(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(KEYINPUT121), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n676), .A2(new_n872), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n875), .A2(new_n723), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT57), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n722), .A2(new_n897), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n866), .B1(new_n730), .B2(new_n731), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n855), .B(KEYINPUT120), .ZN(new_n901));
  OAI22_X1  g700(.A1(new_n901), .A2(new_n854), .B1(new_n323), .B2(new_n861), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n276), .A2(new_n902), .A3(new_n304), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n301), .B1(new_n900), .B2(new_n903), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n324), .A2(new_n355), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n899), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n895), .B1(new_n898), .B2(new_n906), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n487), .B1(new_n907), .B2(new_n355), .ZN(new_n908));
  OAI211_X1 g707(.A(KEYINPUT58), .B(new_n894), .C1(new_n908), .C2(new_n892), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT58), .ZN(new_n910));
  AOI211_X1 g709(.A(new_n356), .B(new_n895), .C1(new_n898), .C2(new_n906), .ZN(new_n911));
  OAI221_X1 g710(.A(new_n893), .B1(KEYINPUT121), .B2(new_n910), .C1(new_n911), .C2(new_n487), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n909), .A2(new_n912), .ZN(G1344gat));
  NAND2_X1  g712(.A1(new_n898), .A2(new_n906), .ZN(new_n914));
  INV_X1    g713(.A(new_n895), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n914), .A2(new_n322), .A3(new_n915), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n488), .A2(KEYINPUT59), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI211_X1 g717(.A(new_n276), .B(new_n304), .C1(new_n862), .C2(new_n856), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n301), .B1(new_n919), .B2(new_n900), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n899), .B1(new_n920), .B2(new_n905), .ZN(new_n921));
  AND3_X1   g720(.A1(new_n276), .A2(new_n902), .A3(new_n304), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n846), .B1(new_n922), .B2(new_n868), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n722), .B1(new_n923), .B2(new_n870), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n921), .B1(new_n924), .B2(KEYINPUT57), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n895), .A2(new_n323), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n488), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT122), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT59), .ZN(new_n929));
  NOR3_X1   g728(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n723), .B1(new_n904), .B2(new_n905), .ZN(new_n931));
  AOI22_X1  g730(.A1(new_n931), .A2(new_n897), .B1(new_n875), .B2(new_n899), .ZN(new_n932));
  INV_X1    g731(.A(new_n926), .ZN(new_n933));
  OAI21_X1  g732(.A(G148gat), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  AOI21_X1  g733(.A(KEYINPUT122), .B1(new_n934), .B2(KEYINPUT59), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n918), .B1(new_n930), .B2(new_n935), .ZN(new_n936));
  INV_X1    g735(.A(new_n891), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n937), .A2(new_n488), .A3(new_n322), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n936), .A2(new_n938), .ZN(G1345gat));
  NAND3_X1  g738(.A1(new_n937), .A2(new_n484), .A3(new_n301), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n907), .A2(new_n301), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n940), .B1(new_n941), .B2(new_n484), .ZN(G1346gat));
  AOI21_X1  g741(.A(G162gat), .B1(new_n937), .B2(new_n733), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n732), .A2(new_n485), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n943), .B1(new_n907), .B2(new_n944), .ZN(G1347gat));
  NOR2_X1   g744(.A1(new_n791), .A2(new_n756), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n871), .A2(new_n946), .ZN(new_n947));
  NOR3_X1   g746(.A1(new_n947), .A2(new_n410), .A3(new_n356), .ZN(new_n948));
  AOI211_X1 g747(.A(new_n685), .B(new_n756), .C1(new_n869), .C2(new_n870), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n949), .A2(new_n722), .A3(new_n680), .ZN(new_n950));
  INV_X1    g749(.A(new_n950), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(new_n355), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n948), .B1(new_n952), .B2(new_n410), .ZN(G1348gat));
  INV_X1    g752(.A(new_n947), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n954), .A2(G176gat), .A3(new_n322), .ZN(new_n955));
  AND2_X1   g754(.A1(new_n955), .A2(KEYINPUT123), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n955), .A2(KEYINPUT123), .ZN(new_n957));
  AOI21_X1  g756(.A(G176gat), .B1(new_n951), .B2(new_n322), .ZN(new_n958));
  NOR3_X1   g757(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(G1349gat));
  NAND3_X1  g758(.A1(new_n951), .A2(new_n404), .A3(new_n301), .ZN(new_n960));
  OAI21_X1  g759(.A(G183gat), .B1(new_n947), .B2(new_n846), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n962), .A2(KEYINPUT60), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT60), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n960), .A2(new_n964), .A3(new_n961), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n963), .A2(new_n965), .ZN(G1350gat));
  NAND3_X1  g765(.A1(new_n951), .A2(new_n264), .A3(new_n733), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT124), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n968), .A2(KEYINPUT61), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n733), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n264), .B1(new_n968), .B2(KEYINPUT61), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n969), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  OAI211_X1 g771(.A(new_n969), .B(new_n971), .C1(new_n947), .C2(new_n732), .ZN(new_n973));
  INV_X1    g772(.A(new_n973), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n967), .B1(new_n972), .B2(new_n974), .ZN(G1351gat));
  NOR2_X1   g774(.A1(new_n768), .A2(new_n722), .ZN(new_n976));
  AND4_X1   g775(.A1(new_n375), .A2(new_n949), .A3(new_n355), .A4(new_n976), .ZN(new_n977));
  XNOR2_X1  g776(.A(new_n977), .B(KEYINPUT125), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n676), .A2(new_n946), .ZN(new_n979));
  NOR3_X1   g778(.A1(new_n932), .A2(new_n356), .A3(new_n979), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n978), .B1(new_n375), .B2(new_n980), .ZN(G1352gat));
  NAND2_X1  g780(.A1(new_n949), .A2(new_n976), .ZN(new_n982));
  NOR2_X1   g781(.A1(new_n323), .A2(G204gat), .ZN(new_n983));
  INV_X1    g782(.A(new_n983), .ZN(new_n984));
  OR3_X1    g783(.A1(new_n982), .A2(KEYINPUT62), .A3(new_n984), .ZN(new_n985));
  OAI21_X1  g784(.A(KEYINPUT62), .B1(new_n982), .B2(new_n984), .ZN(new_n986));
  NOR3_X1   g785(.A1(new_n932), .A2(new_n323), .A3(new_n979), .ZN(new_n987));
  OAI211_X1 g786(.A(new_n985), .B(new_n986), .C1(new_n376), .C2(new_n987), .ZN(G1353gat));
  INV_X1    g787(.A(new_n982), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n989), .A2(new_n370), .A3(new_n301), .ZN(new_n990));
  NAND2_X1  g789(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n991));
  NOR2_X1   g790(.A1(new_n932), .A2(new_n979), .ZN(new_n992));
  AOI21_X1  g791(.A(new_n370), .B1(new_n992), .B2(new_n301), .ZN(new_n993));
  NOR2_X1   g792(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n994));
  INV_X1    g793(.A(new_n994), .ZN(new_n995));
  OAI21_X1  g794(.A(new_n991), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  AOI211_X1 g795(.A(new_n370), .B(new_n994), .C1(new_n992), .C2(new_n301), .ZN(new_n997));
  OAI21_X1  g796(.A(new_n990), .B1(new_n996), .B2(new_n997), .ZN(G1354gat));
  NAND3_X1  g797(.A1(new_n989), .A2(new_n267), .A3(new_n733), .ZN(new_n999));
  NOR3_X1   g798(.A1(new_n932), .A2(new_n732), .A3(new_n979), .ZN(new_n1000));
  OAI21_X1  g799(.A(new_n999), .B1(new_n1000), .B2(new_n267), .ZN(G1355gat));
endmodule


