//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 0 1 1 0 1 1 0 1 1 0 1 0 0 1 0 0 1 1 1 1 0 0 1 0 0 0 0 1 1 1 1 0 0 1 0 0 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:51 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1271, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G77), .ZN(new_n203));
  INV_X1    g0003(.A(G244), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  AOI22_X1  g0005(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n206));
  INV_X1    g0006(.A(G68), .ZN(new_n207));
  INV_X1    g0007(.A(G238), .ZN(new_n208));
  INV_X1    g0008(.A(G107), .ZN(new_n209));
  INV_X1    g0009(.A(G264), .ZN(new_n210));
  OAI221_X1 g0010(.A(new_n206), .B1(new_n207), .B2(new_n208), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  AOI211_X1 g0011(.A(new_n205), .B(new_n211), .C1(G116), .C2(G270), .ZN(new_n212));
  INV_X1    g0012(.A(G50), .ZN(new_n213));
  INV_X1    g0013(.A(G226), .ZN(new_n214));
  INV_X1    g0014(.A(G58), .ZN(new_n215));
  INV_X1    g0015(.A(G232), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n212), .B1(new_n213), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G20), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT1), .Z(new_n220));
  NOR2_X1   g0020(.A1(new_n218), .A2(G13), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n221), .B(G250), .C1(G257), .C2(G264), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT0), .ZN(new_n223));
  AND2_X1   g0023(.A1(KEYINPUT64), .A2(G20), .ZN(new_n224));
  NOR2_X1   g0024(.A1(KEYINPUT64), .A2(G20), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n215), .A2(new_n207), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(G50), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n220), .B(new_n223), .C1(new_n229), .C2(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT65), .ZN(G361));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(new_n216), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(new_n210), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G270), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n237), .B(new_n240), .Z(G358));
  XNOR2_X1  g0041(.A(KEYINPUT66), .B(G107), .ZN(new_n242));
  INV_X1    g0042(.A(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G68), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G50), .B(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n246), .B(new_n249), .Z(G351));
  NAND2_X1  g0050(.A1(G33), .A2(G41), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n228), .A2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT3), .ZN(new_n254));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G222), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n258), .B1(new_n259), .B2(G1698), .ZN(new_n260));
  INV_X1    g0060(.A(G1698), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT68), .ZN(new_n262));
  OR2_X1    g0062(.A1(new_n262), .A2(G223), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(G223), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n261), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  OAI221_X1 g0065(.A(new_n253), .B1(G77), .B2(new_n258), .C1(new_n260), .C2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G1), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n267), .B1(G41), .B2(G45), .ZN(new_n268));
  INV_X1    g0068(.A(G274), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT67), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n227), .B1(new_n272), .B2(new_n251), .ZN(new_n273));
  NAND3_X1  g0073(.A1(KEYINPUT67), .A2(G33), .A3(G41), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(new_n268), .ZN(new_n276));
  OAI211_X1 g0076(.A(new_n266), .B(new_n271), .C1(new_n214), .C2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G200), .ZN(new_n278));
  INV_X1    g0078(.A(new_n277), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G190), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n267), .A2(G13), .A3(G20), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(new_n213), .ZN(new_n283));
  NAND3_X1  g0083(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n284));
  AND3_X1   g0084(.A1(new_n284), .A2(KEYINPUT69), .A3(new_n227), .ZN(new_n285));
  AOI21_X1  g0085(.A(KEYINPUT69), .B1(new_n284), .B2(new_n227), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n287), .A2(new_n282), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n267), .A2(G20), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n288), .A2(G50), .A3(new_n289), .ZN(new_n290));
  XNOR2_X1  g0090(.A(KEYINPUT8), .B(G58), .ZN(new_n291));
  OAI21_X1  g0091(.A(G33), .B1(new_n224), .B2(new_n225), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(KEYINPUT70), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT70), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n294), .B(G33), .C1(new_n224), .C2(new_n225), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n291), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(G20), .A2(G33), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G150), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT71), .ZN(new_n301));
  NOR3_X1   g0101(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n302));
  INV_X1    g0102(.A(G20), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  OAI211_X1 g0104(.A(KEYINPUT71), .B(G20), .C1(new_n230), .C2(G50), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NOR3_X1   g0106(.A1(new_n296), .A2(new_n300), .A3(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n287), .ZN(new_n308));
  NOR3_X1   g0108(.A1(new_n307), .A2(KEYINPUT72), .A3(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT72), .ZN(new_n310));
  INV_X1    g0110(.A(new_n291), .ZN(new_n311));
  XNOR2_X1  g0111(.A(KEYINPUT64), .B(G20), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n294), .B1(new_n312), .B2(G33), .ZN(new_n313));
  INV_X1    g0113(.A(new_n295), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n311), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n300), .ZN(new_n316));
  INV_X1    g0116(.A(new_n306), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n310), .B1(new_n318), .B2(new_n287), .ZN(new_n319));
  OAI211_X1 g0119(.A(new_n283), .B(new_n290), .C1(new_n309), .C2(new_n319), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n320), .A2(KEYINPUT9), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT9), .ZN(new_n322));
  INV_X1    g0122(.A(new_n290), .ZN(new_n323));
  OAI21_X1  g0123(.A(KEYINPUT72), .B1(new_n307), .B2(new_n308), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n318), .A2(new_n310), .A3(new_n287), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n323), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n322), .B1(new_n326), .B2(new_n283), .ZN(new_n327));
  OAI211_X1 g0127(.A(new_n278), .B(new_n280), .C1(new_n321), .C2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(KEYINPUT75), .A2(KEYINPUT10), .ZN(new_n329));
  OR2_X1    g0129(.A1(KEYINPUT75), .A2(KEYINPUT10), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n214), .A2(G1698), .ZN(new_n332));
  AND2_X1   g0132(.A1(KEYINPUT3), .A2(G33), .ZN(new_n333));
  NOR2_X1   g0133(.A1(KEYINPUT3), .A2(G33), .ZN(new_n334));
  OAI221_X1 g0134(.A(new_n332), .B1(G223), .B2(G1698), .C1(new_n333), .C2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(G33), .A2(G87), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n252), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n275), .A2(G232), .A3(new_n268), .ZN(new_n339));
  NAND4_X1  g0139(.A1(new_n338), .A2(G179), .A3(new_n339), .A4(new_n271), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n271), .ZN(new_n341));
  OAI21_X1  g0141(.A(G169), .B1(new_n341), .B2(new_n337), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT16), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n333), .A2(new_n334), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n346), .A2(new_n312), .A3(KEYINPUT7), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n256), .A2(new_n303), .A3(new_n257), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT7), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n207), .B1(new_n347), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(G58), .A2(G68), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(KEYINPUT81), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT81), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n354), .A2(G58), .A3(G68), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n353), .A2(new_n355), .A3(new_n230), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(G20), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n297), .A2(G159), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n345), .B1(new_n351), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(KEYINPUT82), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n284), .A2(new_n227), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT82), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n363), .B(new_n345), .C1(new_n351), .C2(new_n359), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n346), .A2(new_n312), .A3(new_n349), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n348), .A2(KEYINPUT7), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n365), .A2(new_n366), .A3(G68), .ZN(new_n367));
  AOI22_X1  g0167(.A1(new_n356), .A2(G20), .B1(G159), .B2(new_n297), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n367), .A2(KEYINPUT16), .A3(new_n368), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n361), .A2(new_n362), .A3(new_n364), .A4(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n291), .B1(new_n267), .B2(G20), .ZN(new_n371));
  AOI22_X1  g0171(.A1(new_n288), .A2(new_n371), .B1(new_n282), .B2(new_n291), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n344), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n373), .A2(KEYINPUT18), .ZN(new_n374));
  INV_X1    g0174(.A(new_n372), .ZN(new_n375));
  AND2_X1   g0175(.A1(new_n364), .A2(new_n369), .ZN(new_n376));
  INV_X1    g0176(.A(new_n362), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n377), .B1(new_n360), .B2(KEYINPUT82), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n375), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT18), .ZN(new_n380));
  NOR3_X1   g0180(.A1(new_n379), .A2(new_n380), .A3(new_n344), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n374), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(G190), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n338), .A2(new_n383), .A3(new_n339), .A4(new_n271), .ZN(new_n384));
  OR2_X1    g0184(.A1(new_n384), .A2(KEYINPUT83), .ZN(new_n385));
  INV_X1    g0185(.A(G200), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n386), .B1(new_n341), .B2(new_n337), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n384), .A2(new_n387), .A3(KEYINPUT83), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n370), .A2(new_n385), .A3(new_n372), .A4(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT17), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n379), .A2(KEYINPUT17), .A3(new_n385), .A4(new_n388), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n382), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n320), .A2(KEYINPUT9), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n326), .A2(new_n322), .A3(new_n283), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n395), .A2(new_n396), .B1(G190), .B2(new_n279), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n397), .A2(KEYINPUT75), .A3(KEYINPUT10), .A4(new_n278), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n277), .A2(G179), .ZN(new_n399));
  INV_X1    g0199(.A(G169), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n399), .B1(new_n400), .B2(new_n277), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(new_n320), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n331), .A2(new_n394), .A3(new_n398), .A4(new_n402), .ZN(new_n403));
  XNOR2_X1  g0203(.A(KEYINPUT15), .B(G87), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n292), .A2(new_n404), .ZN(new_n405));
  XNOR2_X1  g0205(.A(new_n405), .B(KEYINPUT73), .ZN(new_n406));
  OAI221_X1 g0206(.A(new_n406), .B1(new_n203), .B2(new_n312), .C1(new_n298), .C2(new_n291), .ZN(new_n407));
  AOI22_X1  g0207(.A1(new_n407), .A2(new_n362), .B1(new_n203), .B2(new_n282), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n377), .A2(new_n289), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n409), .A2(new_n203), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  AND2_X1   g0211(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  AND2_X1   g0212(.A1(new_n275), .A2(new_n268), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(G244), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n261), .A2(G232), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n258), .B(new_n415), .C1(new_n208), .C2(new_n261), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n416), .B(new_n253), .C1(G107), .C2(new_n258), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n414), .A2(new_n271), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(new_n400), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(KEYINPUT74), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n418), .A2(G179), .ZN(new_n421));
  MUX2_X1   g0221(.A(new_n420), .B(KEYINPUT74), .S(new_n421), .Z(new_n422));
  NOR2_X1   g0222(.A1(new_n412), .A2(new_n422), .ZN(new_n423));
  XNOR2_X1  g0223(.A(KEYINPUT77), .B(KEYINPUT13), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n214), .A2(new_n261), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n216), .A2(G1698), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n425), .B(new_n426), .C1(new_n333), .C2(new_n334), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT76), .ZN(new_n428));
  NAND2_X1  g0228(.A1(G33), .A2(G97), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n427), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n428), .B1(new_n427), .B2(new_n429), .ZN(new_n432));
  NOR3_X1   g0232(.A1(new_n431), .A2(new_n432), .A3(new_n252), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n271), .B1(new_n276), .B2(new_n208), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n424), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n434), .ZN(new_n436));
  INV_X1    g0236(.A(new_n432), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n437), .A2(new_n253), .A3(new_n430), .ZN(new_n438));
  INV_X1    g0238(.A(new_n424), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n436), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n435), .A2(new_n440), .A3(KEYINPUT78), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n433), .A2(new_n434), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT78), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n442), .A2(new_n443), .A3(new_n439), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n441), .A2(G169), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(KEYINPUT14), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT13), .ZN(new_n447));
  OAI211_X1 g0247(.A(G179), .B(new_n440), .C1(new_n442), .C2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT14), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n441), .A2(new_n444), .A3(new_n449), .A4(G169), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n446), .A2(new_n448), .A3(new_n450), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n298), .A2(new_n213), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n303), .A2(G68), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n293), .A2(new_n295), .ZN(new_n454));
  AOI211_X1 g0254(.A(new_n452), .B(new_n453), .C1(new_n454), .C2(G77), .ZN(new_n455));
  OAI21_X1  g0255(.A(KEYINPUT11), .B1(new_n455), .B2(new_n308), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n454), .A2(G77), .ZN(new_n457));
  INV_X1    g0257(.A(new_n452), .ZN(new_n458));
  INV_X1    g0258(.A(new_n453), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT11), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n460), .A2(new_n461), .A3(new_n287), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n456), .A2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT79), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n464), .B1(new_n281), .B2(G68), .ZN(new_n465));
  XNOR2_X1  g0265(.A(new_n465), .B(KEYINPUT12), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n409), .A2(new_n207), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(KEYINPUT80), .B1(new_n463), .B2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT80), .ZN(new_n470));
  INV_X1    g0270(.A(new_n468), .ZN(new_n471));
  AOI211_X1 g0271(.A(new_n470), .B(new_n471), .C1(new_n456), .C2(new_n462), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n451), .A2(new_n473), .ZN(new_n474));
  OAI211_X1 g0274(.A(G190), .B(new_n440), .C1(new_n442), .C2(new_n447), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n441), .A2(G200), .A3(new_n444), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n475), .B(new_n476), .C1(new_n469), .C2(new_n472), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n418), .A2(G200), .ZN(new_n478));
  OR2_X1    g0278(.A1(new_n418), .A2(new_n383), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n408), .A2(new_n411), .A3(new_n478), .A4(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n474), .A2(new_n477), .A3(new_n480), .ZN(new_n481));
  NOR3_X1   g0281(.A1(new_n403), .A2(new_n423), .A3(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT25), .ZN(new_n483));
  AOI211_X1 g0283(.A(KEYINPUT90), .B(new_n483), .C1(new_n282), .C2(new_n209), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n282), .B(new_n209), .C1(KEYINPUT90), .C2(new_n483), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n485), .B1(KEYINPUT90), .B2(new_n483), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n267), .A2(G33), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n281), .B(new_n487), .C1(new_n285), .C2(new_n286), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  AOI211_X1 g0289(.A(new_n484), .B(new_n486), .C1(new_n489), .C2(G107), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT89), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT22), .ZN(new_n492));
  OAI22_X1  g0292(.A1(new_n225), .A2(new_n224), .B1(new_n333), .B2(new_n334), .ZN(new_n493));
  INV_X1    g0293(.A(G87), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(KEYINPUT23), .A2(G107), .ZN(new_n496));
  AOI21_X1  g0296(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n496), .B1(new_n497), .B2(G20), .ZN(new_n498));
  NOR3_X1   g0298(.A1(new_n224), .A2(new_n225), .A3(KEYINPUT23), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n498), .B1(new_n499), .B2(new_n209), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n258), .A2(new_n312), .A3(KEYINPUT22), .A4(G87), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n495), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(KEYINPUT24), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT24), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n495), .A2(new_n500), .A3(new_n504), .A4(new_n501), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n491), .B1(new_n506), .B2(new_n362), .ZN(new_n507));
  AOI211_X1 g0307(.A(KEYINPUT89), .B(new_n377), .C1(new_n503), .C2(new_n505), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n490), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(G179), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n258), .B1(G257), .B2(new_n261), .ZN(new_n511));
  NOR2_X1   g0311(.A1(G250), .A2(G1698), .ZN(new_n512));
  INV_X1    g0312(.A(G294), .ZN(new_n513));
  OAI22_X1  g0313(.A1(new_n511), .A2(new_n512), .B1(new_n255), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n253), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT5), .ZN(new_n516));
  OAI21_X1  g0316(.A(KEYINPUT86), .B1(new_n516), .B2(G41), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT86), .ZN(new_n518));
  INV_X1    g0318(.A(G41), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n518), .A2(new_n519), .A3(KEYINPUT5), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n517), .A2(new_n520), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n267), .B(G45), .C1(new_n519), .C2(KEYINPUT5), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n521), .A2(new_n523), .B1(new_n273), .B2(new_n274), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(G264), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n269), .B1(new_n273), .B2(new_n274), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n522), .B1(new_n517), .B2(new_n520), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AND4_X1   g0328(.A1(new_n510), .A2(new_n515), .A3(new_n525), .A4(new_n528), .ZN(new_n529));
  AND2_X1   g0329(.A1(new_n515), .A2(new_n525), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n528), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n529), .B1(new_n531), .B2(new_n400), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n509), .A2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n530), .A2(G190), .A3(new_n528), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n490), .B(new_n535), .C1(new_n507), .C2(new_n508), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n531), .A2(G200), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  OAI21_X1  g0339(.A(KEYINPUT91), .B1(new_n534), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n506), .A2(new_n362), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(KEYINPUT89), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n506), .A2(new_n491), .A3(new_n362), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n544), .A2(new_n490), .A3(new_n537), .A4(new_n535), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT91), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n545), .A2(new_n546), .A3(new_n533), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n540), .A2(new_n547), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n303), .A2(G116), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n549), .A2(new_n267), .A3(G13), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n377), .A2(G116), .A3(new_n281), .A4(new_n487), .ZN(new_n551));
  NAND2_X1  g0351(.A1(G33), .A2(G283), .ZN(new_n552));
  INV_X1    g0352(.A(G97), .ZN(new_n553));
  OAI221_X1 g0353(.A(new_n552), .B1(G33), .B2(new_n553), .C1(new_n224), .C2(new_n225), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n549), .B1(new_n227), .B2(new_n284), .ZN(new_n555));
  AND3_X1   g0355(.A1(new_n554), .A2(KEYINPUT20), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(KEYINPUT20), .B1(new_n554), .B2(new_n555), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n550), .B(new_n551), .C1(new_n556), .C2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n524), .A2(G270), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n261), .A2(G257), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n258), .B(new_n560), .C1(new_n210), .C2(new_n261), .ZN(new_n561));
  INV_X1    g0361(.A(G303), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n346), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n561), .A2(new_n253), .A3(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n559), .A2(new_n528), .A3(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n558), .A2(new_n565), .A3(G169), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT21), .ZN(new_n567));
  AND3_X1   g0367(.A1(new_n566), .A2(KEYINPUT88), .A3(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n567), .B1(new_n566), .B2(KEYINPUT88), .ZN(new_n569));
  INV_X1    g0369(.A(new_n558), .ZN(new_n570));
  NOR3_X1   g0370(.A1(new_n570), .A2(new_n510), .A3(new_n565), .ZN(new_n571));
  NOR3_X1   g0371(.A1(new_n568), .A2(new_n569), .A3(new_n571), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n488), .A2(new_n553), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT6), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n553), .A2(new_n209), .ZN(new_n575));
  NOR2_X1   g0375(.A1(G97), .A2(G107), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n574), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n209), .A2(KEYINPUT6), .A3(G97), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n312), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n298), .A2(new_n203), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  AND2_X1   g0382(.A1(new_n347), .A2(new_n350), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n580), .B(new_n582), .C1(new_n583), .C2(new_n209), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n573), .B1(new_n584), .B2(new_n362), .ZN(new_n585));
  OAI211_X1 g0385(.A(G250), .B(G1698), .C1(new_n333), .C2(new_n334), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT4), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n587), .A2(KEYINPUT85), .B1(G33), .B2(G283), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT84), .ZN(new_n590));
  AOI21_X1  g0390(.A(KEYINPUT85), .B1(new_n590), .B2(new_n587), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n204), .A2(G1698), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n591), .B1(new_n258), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n589), .A2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT85), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n261), .A2(G244), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n596), .B1(new_n256), .B2(new_n257), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n595), .B(KEYINPUT4), .C1(new_n597), .C2(KEYINPUT84), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n252), .B1(new_n594), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n524), .A2(G257), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n528), .ZN(new_n601));
  OAI21_X1  g0401(.A(G200), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(new_n598), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n588), .B(new_n586), .C1(new_n597), .C2(new_n591), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n253), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n524), .A2(G257), .B1(new_n527), .B2(new_n526), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n605), .A2(new_n606), .A3(G190), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n282), .A2(new_n553), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n585), .A2(new_n602), .A3(new_n607), .A4(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n573), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n209), .B1(new_n347), .B2(new_n350), .ZN(new_n611));
  NOR3_X1   g0411(.A1(new_n611), .A2(new_n581), .A3(new_n579), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n610), .B(new_n608), .C1(new_n612), .C2(new_n377), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n605), .A2(new_n606), .A3(new_n510), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n400), .B1(new_n599), .B2(new_n601), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  AND2_X1   g0416(.A1(new_n609), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n565), .A2(G200), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n570), .B(new_n618), .C1(new_n383), .C2(new_n565), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n204), .A2(G1698), .ZN(new_n620));
  OAI221_X1 g0420(.A(new_n620), .B1(G238), .B2(G1698), .C1(new_n333), .C2(new_n334), .ZN(new_n621));
  NAND2_X1  g0421(.A1(G33), .A2(G116), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n252), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(G250), .ZN(new_n625));
  INV_X1    g0425(.A(G45), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n625), .B1(new_n626), .B2(G1), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n267), .A2(new_n269), .A3(G45), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n275), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n624), .A2(G190), .A3(new_n629), .ZN(new_n630));
  XNOR2_X1  g0430(.A(new_n630), .B(KEYINPUT87), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n624), .A2(new_n629), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(G200), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT19), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n634), .B1(new_n292), .B2(new_n553), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n494), .A2(new_n553), .A3(new_n209), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n429), .A2(new_n634), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n636), .B1(new_n226), .B2(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n258), .A2(new_n312), .A3(G68), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n635), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  AOI22_X1  g0440(.A1(new_n640), .A2(new_n362), .B1(new_n282), .B2(new_n404), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n489), .A2(G87), .ZN(new_n642));
  AND3_X1   g0442(.A1(new_n633), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n629), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n644), .A2(new_n623), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n510), .ZN(new_n646));
  INV_X1    g0446(.A(new_n404), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n489), .A2(new_n647), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n641), .A2(new_n648), .B1(new_n632), .B2(new_n400), .ZN(new_n649));
  AOI22_X1  g0449(.A1(new_n631), .A2(new_n643), .B1(new_n646), .B2(new_n649), .ZN(new_n650));
  AND4_X1   g0450(.A1(new_n572), .A2(new_n617), .A3(new_n619), .A4(new_n650), .ZN(new_n651));
  AND3_X1   g0451(.A1(new_n482), .A2(new_n548), .A3(new_n651), .ZN(G372));
  INV_X1    g0452(.A(KEYINPUT26), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n641), .A2(new_n648), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n632), .A2(new_n400), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n654), .A2(new_n655), .A3(new_n646), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n633), .A2(new_n641), .A3(new_n642), .A4(new_n630), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n653), .B1(new_n658), .B2(new_n616), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(KEYINPUT93), .ZN(new_n660));
  INV_X1    g0460(.A(new_n616), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n650), .A2(KEYINPUT26), .A3(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT93), .ZN(new_n663));
  OAI211_X1 g0463(.A(new_n663), .B(new_n653), .C1(new_n658), .C2(new_n616), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n660), .A2(new_n662), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(new_n656), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(KEYINPUT92), .B1(new_n533), .B2(new_n572), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n658), .ZN(new_n670));
  OAI211_X1 g0470(.A(new_n617), .B(new_n670), .C1(new_n536), .C2(new_n538), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n533), .A2(new_n572), .A3(KEYINPUT92), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n669), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n667), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n482), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g0476(.A(KEYINPUT94), .B(KEYINPUT95), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n678), .B1(new_n374), .B2(new_n381), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n373), .A2(KEYINPUT18), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n380), .B1(new_n379), .B2(new_n344), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n680), .A2(new_n681), .A3(new_n677), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  AOI22_X1  g0483(.A1(new_n423), .A2(new_n477), .B1(new_n451), .B2(new_n473), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n683), .B1(new_n684), .B2(new_n393), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n331), .A2(new_n398), .ZN(new_n686));
  AOI22_X1  g0486(.A1(new_n685), .A2(new_n686), .B1(new_n320), .B2(new_n401), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n676), .A2(new_n687), .ZN(G369));
  NAND2_X1  g0488(.A1(new_n312), .A2(G13), .ZN(new_n689));
  OR3_X1    g0489(.A1(new_n689), .A2(KEYINPUT27), .A3(G1), .ZN(new_n690));
  OAI21_X1  g0490(.A(KEYINPUT27), .B1(new_n689), .B2(G1), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n690), .A2(new_n691), .A3(G213), .ZN(new_n692));
  INV_X1    g0492(.A(G343), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n509), .A2(new_n694), .ZN(new_n695));
  AND3_X1   g0495(.A1(new_n545), .A2(new_n546), .A3(new_n533), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n546), .B1(new_n545), .B2(new_n533), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n695), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(KEYINPUT97), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT97), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n548), .A2(new_n700), .A3(new_n695), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n572), .A2(new_n694), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n699), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n694), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n534), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n699), .A2(new_n701), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n533), .A2(new_n704), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n694), .A2(new_n558), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n572), .A2(new_n619), .A3(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n713), .B1(new_n572), .B2(new_n712), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT96), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n714), .A2(new_n715), .A3(G330), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n715), .B1(new_n714), .B2(G330), .ZN(new_n718));
  OR2_X1    g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n711), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n707), .A2(new_n720), .ZN(G399));
  INV_X1    g0521(.A(new_n221), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(G41), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n636), .A2(G116), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n724), .A2(G1), .A3(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n726), .B1(new_n231), .B2(new_n724), .ZN(new_n727));
  XNOR2_X1  g0527(.A(new_n727), .B(KEYINPUT28), .ZN(new_n728));
  XNOR2_X1  g0528(.A(new_n656), .B(KEYINPUT98), .ZN(new_n729));
  OAI21_X1  g0529(.A(KEYINPUT26), .B1(new_n658), .B2(new_n616), .ZN(new_n730));
  AND2_X1   g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n650), .A2(new_n653), .A3(new_n661), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n533), .A2(new_n572), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  OAI211_X1 g0534(.A(new_n731), .B(new_n732), .C1(new_n734), .C2(new_n671), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n735), .A2(KEYINPUT29), .A3(new_n704), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n694), .B1(new_n667), .B2(new_n674), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n736), .B1(new_n737), .B2(KEYINPUT29), .ZN(new_n738));
  OAI211_X1 g0538(.A(new_n651), .B(new_n704), .C1(new_n696), .C2(new_n697), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n565), .A2(new_n510), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n599), .A2(new_n601), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n740), .A2(new_n741), .A3(new_n530), .A4(new_n645), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT30), .ZN(new_n743));
  OR2_X1    g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n742), .A2(new_n743), .ZN(new_n745));
  INV_X1    g0545(.A(new_n741), .ZN(new_n746));
  AND2_X1   g0546(.A1(new_n565), .A2(new_n510), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n531), .A2(new_n746), .A3(new_n747), .A4(new_n632), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n744), .A2(new_n745), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(new_n694), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(KEYINPUT31), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT31), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n749), .A2(new_n752), .A3(new_n694), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n739), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(G330), .ZN(new_n756));
  AND2_X1   g0556(.A1(new_n738), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n728), .B1(new_n757), .B2(G1), .ZN(G364));
  NAND3_X1  g0558(.A1(new_n312), .A2(G13), .A3(G45), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR3_X1   g0560(.A1(new_n760), .A2(new_n723), .A3(new_n267), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n312), .A2(new_n510), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n383), .A2(new_n386), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n258), .B1(new_n766), .B2(G326), .ZN(new_n767));
  INV_X1    g0567(.A(G283), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n386), .A2(G190), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n226), .A2(new_n510), .A3(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(G311), .ZN(new_n771));
  NOR2_X1   g0571(.A1(G190), .A2(G200), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n763), .A2(new_n772), .ZN(new_n773));
  OAI221_X1 g0573(.A(new_n767), .B1(new_n768), .B2(new_n770), .C1(new_n771), .C2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n383), .A2(G200), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n226), .B1(new_n776), .B2(G179), .ZN(new_n777));
  INV_X1    g0577(.A(KEYINPUT103), .ZN(new_n778));
  OR2_X1    g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n777), .A2(new_n778), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n774), .B1(G294), .B2(new_n782), .ZN(new_n783));
  XOR2_X1   g0583(.A(KEYINPUT104), .B(G317), .Z(new_n784));
  XNOR2_X1  g0584(.A(new_n784), .B(KEYINPUT33), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n763), .A2(new_n769), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n226), .A2(new_n510), .A3(new_n772), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n785), .A2(new_n787), .B1(G329), .B2(new_n789), .ZN(new_n790));
  AND2_X1   g0590(.A1(new_n783), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n764), .A2(G20), .A3(new_n510), .ZN(new_n792));
  INV_X1    g0592(.A(G322), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n763), .A2(new_n775), .ZN(new_n794));
  OAI221_X1 g0594(.A(new_n791), .B1(new_n562), .B2(new_n792), .C1(new_n793), .C2(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n782), .A2(G97), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n796), .B1(new_n207), .B2(new_n786), .ZN(new_n797));
  INV_X1    g0597(.A(G159), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n788), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(KEYINPUT32), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n801), .B1(new_n215), .B2(new_n794), .ZN(new_n802));
  INV_X1    g0602(.A(new_n792), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(G87), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n804), .B1(new_n773), .B2(new_n203), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n258), .B1(new_n799), .B2(new_n800), .ZN(new_n806));
  NOR4_X1   g0606(.A1(new_n797), .A2(new_n802), .A3(new_n805), .A4(new_n806), .ZN(new_n807));
  OAI221_X1 g0607(.A(new_n807), .B1(new_n213), .B2(new_n765), .C1(new_n209), .C2(new_n770), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n795), .A2(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n227), .B1(G20), .B2(new_n400), .ZN(new_n810));
  NOR2_X1   g0610(.A1(G13), .A2(G33), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n812), .A2(G20), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n813), .A2(new_n810), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n258), .A2(G355), .A3(new_n221), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n249), .A2(G45), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n816), .B(KEYINPUT101), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n722), .A2(new_n258), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n818), .B1(G45), .B2(new_n231), .ZN(new_n819));
  XOR2_X1   g0619(.A(new_n819), .B(KEYINPUT102), .Z(new_n820));
  OAI221_X1 g0620(.A(new_n815), .B1(G116), .B2(new_n221), .C1(new_n817), .C2(new_n820), .ZN(new_n821));
  AOI22_X1  g0621(.A1(new_n809), .A2(new_n810), .B1(new_n814), .B2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n813), .ZN(new_n823));
  OR2_X1    g0623(.A1(new_n714), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n762), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT100), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n719), .B(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n714), .A2(G330), .ZN(new_n829));
  XOR2_X1   g0629(.A(new_n829), .B(KEYINPUT99), .Z(new_n830));
  AND2_X1   g0630(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n826), .B1(new_n831), .B2(new_n761), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(KEYINPUT105), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT105), .ZN(new_n834));
  OAI211_X1 g0634(.A(new_n834), .B(new_n826), .C1(new_n831), .C2(new_n761), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n833), .A2(new_n835), .ZN(G396));
  NAND2_X1  g0636(.A1(new_n675), .A2(new_n704), .ZN(new_n837));
  OR2_X1    g0637(.A1(new_n412), .A2(new_n422), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n480), .B1(new_n412), .B2(new_n704), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NOR3_X1   g0640(.A1(new_n412), .A2(new_n422), .A3(new_n694), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n837), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n841), .B1(new_n838), .B2(new_n839), .ZN(new_n845));
  AND3_X1   g0645(.A1(new_n533), .A2(KEYINPUT92), .A3(new_n572), .ZN(new_n846));
  NOR3_X1   g0646(.A1(new_n846), .A2(new_n668), .A3(new_n671), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n704), .B(new_n845), .C1(new_n847), .C2(new_n666), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n844), .A2(new_n848), .ZN(new_n849));
  OR2_X1    g0649(.A1(new_n849), .A2(new_n756), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(new_n756), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n850), .A2(new_n762), .A3(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n794), .ZN(new_n853));
  XNOR2_X1  g0653(.A(KEYINPUT106), .B(G143), .ZN(new_n854));
  AOI22_X1  g0654(.A1(G150), .A2(new_n787), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(G137), .ZN(new_n856));
  OAI221_X1 g0656(.A(new_n855), .B1(new_n856), .B2(new_n765), .C1(new_n798), .C2(new_n773), .ZN(new_n857));
  XOR2_X1   g0657(.A(KEYINPUT107), .B(KEYINPUT34), .Z(new_n858));
  XNOR2_X1  g0658(.A(new_n857), .B(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n770), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(G68), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n346), .B1(new_n803), .B2(G50), .ZN(new_n862));
  INV_X1    g0662(.A(G132), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n861), .B(new_n862), .C1(new_n863), .C2(new_n788), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n864), .B1(new_n782), .B2(G58), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n859), .A2(new_n865), .ZN(new_n866));
  OAI22_X1  g0666(.A1(new_n768), .A2(new_n786), .B1(new_n765), .B2(new_n562), .ZN(new_n867));
  OAI221_X1 g0667(.A(new_n796), .B1(new_n243), .B2(new_n773), .C1(new_n513), .C2(new_n794), .ZN(new_n868));
  AOI211_X1 g0668(.A(new_n867), .B(new_n868), .C1(G107), .C2(new_n803), .ZN(new_n869));
  OAI221_X1 g0669(.A(new_n869), .B1(new_n494), .B2(new_n770), .C1(new_n771), .C2(new_n788), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n866), .B1(new_n870), .B2(new_n258), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(new_n810), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n810), .A2(new_n811), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(new_n203), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n843), .A2(new_n811), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n872), .A2(new_n761), .A3(new_n874), .A4(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n852), .A2(new_n876), .ZN(G384));
  NAND2_X1  g0677(.A1(new_n577), .A2(new_n578), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n228), .B(new_n226), .C1(new_n878), .C2(KEYINPUT35), .ZN(new_n879));
  AOI211_X1 g0679(.A(new_n243), .B(new_n879), .C1(KEYINPUT35), .C2(new_n878), .ZN(new_n880));
  XOR2_X1   g0680(.A(new_n880), .B(KEYINPUT36), .Z(new_n881));
  NAND2_X1  g0681(.A1(new_n353), .A2(new_n355), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n230), .A2(G50), .A3(G77), .ZN(new_n883));
  OAI22_X1  g0683(.A1(new_n882), .A2(new_n883), .B1(G50), .B2(new_n207), .ZN(new_n884));
  INV_X1    g0684(.A(G13), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n884), .A2(G1), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n881), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n887), .B(KEYINPUT108), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n843), .B1(new_n739), .B2(new_n754), .ZN(new_n889));
  INV_X1    g0689(.A(new_n477), .ZN(new_n890));
  OAI211_X1 g0690(.A(new_n473), .B(new_n694), .C1(new_n890), .C2(new_n451), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n473), .A2(new_n694), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n474), .A2(new_n477), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  AND2_X1   g0694(.A1(new_n889), .A2(new_n894), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n391), .A2(new_n392), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n679), .A2(new_n896), .A3(new_n682), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n692), .B1(new_n370), .B2(new_n372), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n373), .ZN(new_n900));
  AND3_X1   g0700(.A1(new_n370), .A2(new_n385), .A3(new_n372), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n898), .B1(new_n901), .B2(new_n388), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n389), .B(KEYINPUT94), .C1(new_n379), .C2(new_n692), .ZN(new_n903));
  AOI22_X1  g0703(.A1(new_n900), .A2(new_n902), .B1(new_n903), .B2(KEYINPUT37), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n389), .B1(new_n379), .B2(new_n692), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT37), .ZN(new_n906));
  NOR4_X1   g0706(.A1(new_n905), .A2(KEYINPUT94), .A3(new_n906), .A4(new_n373), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n899), .A2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT38), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n369), .A2(new_n287), .ZN(new_n912));
  AOI21_X1  g0712(.A(KEYINPUT16), .B1(new_n367), .B2(new_n368), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n372), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(KEYINPUT109), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT109), .ZN(new_n916));
  OAI211_X1 g0716(.A(new_n916), .B(new_n372), .C1(new_n912), .C2(new_n913), .ZN(new_n917));
  INV_X1    g0717(.A(new_n692), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n915), .B(new_n917), .C1(new_n343), .C2(new_n918), .ZN(new_n919));
  AND3_X1   g0719(.A1(new_n919), .A2(KEYINPUT37), .A3(new_n389), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n902), .A2(new_n900), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n920), .B1(new_n921), .B2(new_n906), .ZN(new_n922));
  AND2_X1   g0722(.A1(new_n915), .A2(new_n917), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n918), .B(new_n923), .C1(new_n382), .C2(new_n393), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n922), .A2(new_n924), .A3(KEYINPUT38), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n911), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n895), .A2(new_n926), .A3(KEYINPUT40), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT40), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n889), .A2(new_n894), .ZN(new_n929));
  AND3_X1   g0729(.A1(new_n922), .A2(new_n924), .A3(KEYINPUT38), .ZN(new_n930));
  AOI21_X1  g0730(.A(KEYINPUT38), .B1(new_n922), .B2(new_n924), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n928), .B1(new_n929), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n927), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n482), .A2(new_n755), .ZN(new_n935));
  XOR2_X1   g0735(.A(new_n934), .B(new_n935), .Z(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(G330), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n683), .A2(new_n918), .ZN(new_n938));
  AND2_X1   g0738(.A1(new_n891), .A2(new_n893), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n939), .B1(new_n848), .B2(new_n842), .ZN(new_n940));
  INV_X1    g0740(.A(new_n931), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(new_n925), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n938), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT39), .ZN(new_n944));
  AOI21_X1  g0744(.A(KEYINPUT38), .B1(new_n899), .B2(new_n908), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n944), .B1(new_n945), .B2(new_n930), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n941), .A2(KEYINPUT39), .A3(new_n925), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n474), .A2(new_n694), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n946), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n943), .A2(new_n949), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n937), .B(new_n950), .ZN(new_n951));
  OAI211_X1 g0751(.A(new_n482), .B(new_n736), .C1(KEYINPUT29), .C2(new_n737), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(new_n687), .ZN(new_n953));
  XOR2_X1   g0753(.A(new_n951), .B(new_n953), .Z(new_n954));
  NAND2_X1  g0754(.A1(new_n689), .A2(G1), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n888), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT110), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n956), .B(new_n957), .ZN(G367));
  NAND2_X1  g0758(.A1(new_n613), .A2(new_n694), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n617), .A2(new_n959), .ZN(new_n960));
  OR3_X1    g0760(.A1(new_n703), .A2(KEYINPUT42), .A3(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n616), .B1(new_n960), .B2(new_n533), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(new_n704), .ZN(new_n963));
  OAI21_X1  g0763(.A(KEYINPUT42), .B1(new_n703), .B2(new_n960), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n961), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n704), .B1(new_n641), .B2(new_n642), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT111), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(new_n670), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n656), .B2(new_n967), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(KEYINPUT43), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n965), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n661), .A2(new_n694), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n960), .A2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n720), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n971), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n969), .A2(KEYINPUT43), .ZN(new_n977));
  INV_X1    g0777(.A(new_n975), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n978), .A2(new_n970), .A3(new_n965), .ZN(new_n979));
  AND3_X1   g0779(.A1(new_n976), .A2(new_n977), .A3(new_n979), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n977), .B1(new_n976), .B2(new_n979), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n723), .B(KEYINPUT41), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT45), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n706), .B2(new_n974), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n703), .A2(KEYINPUT45), .A3(new_n705), .A4(new_n973), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n973), .B1(new_n703), .B2(new_n705), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT44), .ZN(new_n990));
  OR2_X1    g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n989), .A2(new_n990), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n988), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n720), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(new_n702), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n700), .B1(new_n548), .B2(new_n695), .ZN(new_n997));
  INV_X1    g0797(.A(new_n695), .ZN(new_n998));
  AOI211_X1 g0798(.A(KEYINPUT97), .B(new_n998), .C1(new_n540), .C2(new_n547), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n710), .B(new_n996), .C1(new_n997), .C2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(KEYINPUT112), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT112), .ZN(new_n1002));
  NAND4_X1  g0802(.A1(new_n708), .A2(new_n1002), .A3(new_n710), .A4(new_n996), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n1001), .A2(new_n703), .A3(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1004), .A2(new_n828), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n1001), .A2(new_n719), .A3(new_n703), .A4(new_n1003), .ZN(new_n1006));
  AND3_X1   g0806(.A1(new_n1005), .A2(new_n757), .A3(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n989), .B(KEYINPUT44), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1008), .A2(new_n720), .A3(new_n988), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n995), .A2(new_n1007), .A3(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n984), .B1(new_n1010), .B2(new_n757), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n760), .A2(new_n267), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n982), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n770), .A2(new_n553), .ZN(new_n1015));
  AOI211_X1 g0815(.A(new_n258), .B(new_n1015), .C1(G317), .C2(new_n789), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n1016), .A2(KEYINPUT114), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n792), .A2(new_n243), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT46), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n768), .A2(new_n773), .B1(new_n786), .B2(new_n513), .ZN(new_n1020));
  NOR3_X1   g0820(.A1(new_n1017), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n1016), .A2(KEYINPUT114), .B1(G311), .B2(new_n766), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n1021), .B(new_n1022), .C1(new_n562), .C2(new_n794), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(G107), .B2(new_n782), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n789), .A2(G137), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n792), .A2(new_n215), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n782), .A2(G68), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n773), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n346), .B1(new_n1028), .B2(G50), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n766), .A2(new_n854), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n853), .A2(G150), .B1(G77), .B2(new_n860), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1027), .A2(new_n1029), .A3(new_n1030), .A4(new_n1031), .ZN(new_n1032));
  AOI211_X1 g0832(.A(new_n1026), .B(new_n1032), .C1(G159), .C2(new_n787), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1024), .B1(new_n1025), .B2(new_n1033), .ZN(new_n1034));
  XOR2_X1   g0834(.A(new_n1034), .B(KEYINPUT47), .Z(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(new_n810), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n818), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n814), .B1(new_n221), .B2(new_n404), .C1(new_n240), .C2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1038), .A2(new_n761), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT113), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1036), .B(new_n1040), .C1(new_n823), .C2(new_n969), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1014), .A2(new_n1041), .ZN(G387));
  AOI21_X1  g0842(.A(new_n757), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1043));
  NOR3_X1   g0843(.A1(new_n1007), .A2(new_n1043), .A3(new_n724), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n792), .A2(new_n203), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n258), .B1(new_n299), .B2(new_n788), .C1(new_n765), .C2(new_n798), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n1046), .B(new_n1047), .C1(new_n311), .C2(new_n787), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1015), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n853), .A2(G50), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n782), .A2(new_n647), .B1(G68), .B2(new_n1028), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1048), .A2(new_n1049), .A3(new_n1050), .A4(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(G317), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n562), .A2(new_n773), .B1(new_n794), .B2(new_n1053), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n1054), .B(KEYINPUT116), .Z(new_n1055));
  OAI221_X1 g0855(.A(new_n1055), .B1(new_n771), .B2(new_n786), .C1(new_n793), .C2(new_n765), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT48), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n1057), .B1(new_n768), .B2(new_n781), .C1(new_n513), .C2(new_n792), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT49), .Z(new_n1059));
  AOI21_X1  g0859(.A(new_n258), .B1(new_n789), .B2(G326), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(new_n243), .B2(new_n770), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1052), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1062), .A2(new_n810), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n237), .A2(G45), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT115), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n291), .A2(G50), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT50), .ZN(new_n1067));
  AOI21_X1  g0867(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1067), .A2(new_n725), .A3(new_n1068), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1065), .A2(new_n818), .A3(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n258), .A2(new_n221), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n1070), .B1(G107), .B2(new_n221), .C1(new_n725), .C2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n762), .B1(new_n1072), .B2(new_n814), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n1063), .B(new_n1073), .C1(new_n711), .C2(new_n823), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1005), .A2(new_n1013), .A3(new_n1006), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1045), .A2(new_n1077), .ZN(G393));
  NAND3_X1  g0878(.A1(new_n1005), .A2(new_n757), .A3(new_n1006), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1009), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n720), .B1(new_n1008), .B2(new_n988), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1079), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1082), .A2(new_n723), .A3(new_n1010), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n771), .A2(new_n794), .B1(new_n765), .B2(new_n1053), .ZN(new_n1084));
  XOR2_X1   g0884(.A(new_n1084), .B(KEYINPUT52), .Z(new_n1085));
  AOI21_X1  g0885(.A(new_n1085), .B1(G303), .B2(new_n787), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n782), .A2(G116), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1028), .A2(G294), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n770), .A2(new_n209), .B1(new_n768), .B2(new_n792), .ZN(new_n1089));
  AOI211_X1 g0889(.A(new_n258), .B(new_n1089), .C1(G322), .C2(new_n789), .ZN(new_n1090));
  NAND4_X1  g0890(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .A4(new_n1090), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n299), .A2(new_n765), .B1(new_n794), .B2(new_n798), .ZN(new_n1092));
  XOR2_X1   g0892(.A(new_n1092), .B(KEYINPUT51), .Z(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(G50), .B2(new_n787), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n789), .A2(new_n854), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n782), .A2(G77), .B1(G87), .B2(new_n860), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n346), .B1(new_n803), .B2(G68), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n1094), .A2(new_n1095), .A3(new_n1096), .A4(new_n1097), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n773), .A2(new_n291), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1091), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n762), .B1(new_n1100), .B2(new_n810), .ZN(new_n1101));
  OAI221_X1 g0901(.A(new_n814), .B1(new_n553), .B2(new_n221), .C1(new_n246), .C2(new_n1037), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n1101), .B(new_n1102), .C1(new_n823), .C2(new_n973), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1103), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1104), .B1(new_n1105), .B2(new_n1013), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1083), .A2(new_n1106), .ZN(G390));
  AND3_X1   g0907(.A1(new_n889), .A2(G330), .A3(new_n894), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n848), .A2(new_n842), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(new_n894), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n948), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n1110), .A2(new_n1111), .B1(new_n946), .B2(new_n947), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n735), .A2(new_n704), .A3(new_n840), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n939), .B1(new_n842), .B2(new_n1113), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n945), .A2(new_n930), .ZN(new_n1115));
  NOR3_X1   g0915(.A1(new_n1114), .A2(new_n1115), .A3(new_n948), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1108), .B1(new_n1112), .B2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(KEYINPUT39), .B1(new_n911), .B2(new_n925), .ZN(new_n1118));
  NOR3_X1   g0918(.A1(new_n930), .A2(new_n931), .A3(new_n944), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n1118), .A2(new_n1119), .B1(new_n940), .B2(new_n948), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n889), .A2(G330), .A3(new_n894), .ZN(new_n1121));
  AND2_X1   g0921(.A1(new_n1113), .A2(new_n842), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n926), .B(new_n1111), .C1(new_n939), .C2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1120), .A2(new_n1121), .A3(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1117), .A2(new_n1124), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n403), .A2(new_n423), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n481), .ZN(new_n1127));
  NAND4_X1  g0927(.A1(new_n1126), .A2(G330), .A3(new_n755), .A4(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n482), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1128), .B(new_n687), .C1(new_n738), .C2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n894), .B1(new_n889), .B2(G330), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1109), .B1(new_n1108), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n889), .A2(G330), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(new_n939), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1134), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1130), .B1(new_n1132), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1125), .A2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1117), .A2(new_n1136), .A3(new_n1124), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1138), .A2(new_n723), .A3(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1117), .A2(new_n1124), .A3(new_n1013), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n811), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n873), .A2(new_n291), .ZN(new_n1143));
  INV_X1    g0943(.A(G128), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n1144), .A2(new_n765), .B1(new_n794), .B2(new_n863), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1145), .B(KEYINPUT117), .ZN(new_n1146));
  XOR2_X1   g0946(.A(KEYINPUT54), .B(G143), .Z(new_n1147));
  NAND2_X1  g0947(.A1(new_n1028), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n789), .A2(G125), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n860), .A2(G50), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n1146), .A2(new_n1148), .A3(new_n1149), .A4(new_n1150), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n786), .A2(new_n856), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n781), .A2(new_n798), .ZN(new_n1153));
  OR3_X1    g0953(.A1(new_n792), .A2(KEYINPUT53), .A3(new_n299), .ZN(new_n1154));
  OAI21_X1  g0954(.A(KEYINPUT53), .B1(new_n792), .B2(new_n299), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1154), .A2(new_n1155), .A3(new_n258), .ZN(new_n1156));
  NOR4_X1   g0956(.A1(new_n1151), .A2(new_n1152), .A3(new_n1153), .A4(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n782), .A2(G77), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n258), .B1(new_n787), .B2(G107), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1158), .A2(new_n804), .A3(new_n861), .A4(new_n1159), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n794), .A2(new_n243), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n773), .A2(new_n553), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n765), .A2(new_n768), .B1(new_n513), .B2(new_n788), .ZN(new_n1163));
  NOR4_X1   g0963(.A1(new_n1160), .A2(new_n1161), .A3(new_n1162), .A4(new_n1163), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n810), .B1(new_n1157), .B2(new_n1164), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1142), .A2(new_n761), .A3(new_n1143), .A4(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT118), .ZN(new_n1167));
  AND3_X1   g0967(.A1(new_n1141), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1167), .B1(new_n1141), .B2(new_n1166), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1140), .B1(new_n1168), .B2(new_n1169), .ZN(G378));
  OAI21_X1  g0970(.A(new_n213), .B1(new_n333), .B2(G41), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n803), .A2(new_n1147), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n782), .A2(G150), .B1(G125), .B2(new_n766), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT120), .ZN(new_n1174));
  AND2_X1   g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1176));
  OAI221_X1 g0976(.A(new_n1172), .B1(new_n1144), .B2(new_n794), .C1(new_n1175), .C2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(G137), .B2(new_n1028), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1178), .B1(new_n863), .B2(new_n786), .ZN(new_n1179));
  OR2_X1    g0979(.A1(new_n1179), .A2(KEYINPUT59), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n860), .A2(G159), .ZN(new_n1181));
  AOI21_X1  g0981(.A(G41), .B1(new_n789), .B2(G124), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1180), .A2(new_n255), .A3(new_n1181), .A4(new_n1182), .ZN(new_n1183));
  AND2_X1   g0983(.A1(new_n1179), .A2(KEYINPUT59), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1171), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n765), .A2(new_n243), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n258), .B(new_n1046), .C1(G58), .C2(new_n860), .ZN(new_n1187));
  OAI221_X1 g0987(.A(new_n1187), .B1(new_n768), .B2(new_n788), .C1(new_n404), .C2(new_n773), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n1186), .B(new_n1188), .C1(G97), .C2(new_n787), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n853), .A2(G107), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n1190), .B(KEYINPUT119), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1189), .A2(new_n519), .A3(new_n1027), .A4(new_n1191), .ZN(new_n1192));
  XOR2_X1   g0992(.A(new_n1192), .B(KEYINPUT58), .Z(new_n1193));
  OAI21_X1  g0993(.A(new_n810), .B1(new_n1185), .B2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n873), .A2(new_n213), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n331), .A2(new_n398), .A3(new_n402), .ZN(new_n1196));
  XOR2_X1   g0996(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n320), .A2(new_n918), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1197), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n331), .A2(new_n398), .A3(new_n402), .A4(new_n1201), .ZN(new_n1202));
  AND3_X1   g1002(.A1(new_n1198), .A2(new_n1200), .A3(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1200), .B1(new_n1198), .B2(new_n1202), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n811), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1194), .A2(new_n761), .A3(new_n1195), .A4(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n927), .A2(new_n933), .A3(G330), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT121), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1210));
  AND3_X1   g1010(.A1(new_n943), .A2(new_n1210), .A3(new_n949), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1210), .B1(new_n943), .B2(new_n949), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1208), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1210), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n950), .A2(new_n1214), .ZN(new_n1215));
  AND3_X1   g1015(.A1(new_n927), .A2(G330), .A3(new_n933), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n943), .A2(new_n1210), .A3(new_n949), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1215), .A2(new_n1216), .A3(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1213), .A2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1207), .B1(new_n1219), .B2(new_n1013), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1130), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1139), .A2(new_n1221), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1222), .A2(new_n1219), .A3(KEYINPUT57), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(new_n723), .ZN(new_n1224));
  AOI21_X1  g1024(.A(KEYINPUT57), .B1(new_n1222), .B2(new_n1219), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1220), .B1(new_n1224), .B2(new_n1225), .ZN(G375));
  NAND2_X1  g1026(.A1(new_n1132), .A2(new_n1135), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1227), .A2(new_n1013), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT122), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n939), .A2(new_n811), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n873), .A2(new_n207), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n794), .A2(new_n856), .B1(new_n215), .B2(new_n770), .ZN(new_n1233));
  AOI211_X1 g1033(.A(new_n346), .B(new_n1233), .C1(new_n787), .C2(new_n1147), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1028), .A2(G150), .ZN(new_n1235));
  OAI22_X1  g1035(.A1(new_n788), .A2(new_n1144), .B1(new_n798), .B2(new_n792), .ZN(new_n1236));
  XOR2_X1   g1036(.A(new_n1236), .B(KEYINPUT123), .Z(new_n1237));
  NAND2_X1  g1037(.A1(new_n782), .A2(G50), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1234), .A2(new_n1235), .A3(new_n1237), .A4(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1239), .B1(G132), .B2(new_n766), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n782), .A2(new_n647), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n860), .A2(G77), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n803), .A2(G97), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n258), .B1(new_n1028), .B2(G107), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1241), .A2(new_n1242), .A3(new_n1243), .A4(new_n1244), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n786), .A2(new_n243), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n788), .A2(new_n562), .ZN(new_n1247));
  OAI22_X1  g1047(.A1(new_n768), .A2(new_n794), .B1(new_n765), .B2(new_n513), .ZN(new_n1248));
  NOR4_X1   g1048(.A1(new_n1245), .A2(new_n1246), .A3(new_n1247), .A4(new_n1248), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n810), .B1(new_n1240), .B2(new_n1249), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1231), .A2(new_n761), .A3(new_n1232), .A4(new_n1250), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1227), .A2(KEYINPUT122), .A3(new_n1013), .ZN(new_n1252));
  AND3_X1   g1052(.A1(new_n1230), .A2(new_n1251), .A3(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1132), .A2(new_n1135), .A3(new_n1130), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1137), .A2(new_n983), .A3(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1253), .A2(new_n1255), .ZN(G381));
  NOR2_X1   g1056(.A1(G387), .A2(G390), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(G381), .A2(G384), .ZN(new_n1258));
  AND2_X1   g1058(.A1(new_n1141), .A2(new_n1166), .ZN(new_n1259));
  AND2_X1   g1059(.A1(new_n1140), .A2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(G375), .A2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(G396), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1263), .A2(new_n1045), .A3(new_n1077), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1257), .A2(new_n1258), .A3(new_n1262), .A4(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT124), .ZN(new_n1267));
  AND2_X1   g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1269));
  OR2_X1    g1069(.A1(new_n1268), .A2(new_n1269), .ZN(G407));
  NAND2_X1  g1070(.A1(new_n1262), .A2(new_n693), .ZN(new_n1271));
  OAI211_X1 g1071(.A(G213), .B(new_n1271), .C1(new_n1268), .C2(new_n1269), .ZN(G409));
  INV_X1    g1072(.A(G213), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1273), .A2(G343), .ZN(new_n1274));
  OAI211_X1 g1074(.A(G378), .B(new_n1220), .C1(new_n1224), .C2(new_n1225), .ZN(new_n1275));
  AND3_X1   g1075(.A1(new_n1222), .A2(new_n1219), .A3(new_n983), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1219), .A2(new_n1013), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(new_n1206), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1260), .B1(new_n1276), .B2(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1274), .B1(new_n1275), .B2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT62), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT60), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1254), .A2(new_n1282), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1132), .A2(new_n1135), .A3(new_n1130), .A4(KEYINPUT60), .ZN(new_n1284));
  AND4_X1   g1084(.A1(new_n723), .A2(new_n1283), .A3(new_n1137), .A4(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1230), .A2(new_n1251), .A3(new_n1252), .ZN(new_n1286));
  OAI211_X1 g1086(.A(new_n852), .B(new_n876), .C1(new_n1285), .C2(new_n1286), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1283), .A2(new_n1137), .A3(new_n723), .A4(new_n1284), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1253), .A2(G384), .A3(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1287), .A2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  AND3_X1   g1091(.A1(new_n1280), .A2(new_n1281), .A3(new_n1291), .ZN(new_n1292));
  XOR2_X1   g1092(.A(KEYINPUT127), .B(KEYINPUT61), .Z(new_n1293));
  NAND2_X1  g1093(.A1(new_n1274), .A2(G2897), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1290), .A2(new_n1295), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1287), .A2(new_n1289), .A3(new_n1294), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1293), .B1(new_n1280), .B2(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1281), .B1(new_n1280), .B2(new_n1291), .ZN(new_n1300));
  NOR3_X1   g1100(.A1(new_n1292), .A2(new_n1299), .A3(new_n1300), .ZN(new_n1301));
  AND3_X1   g1101(.A1(new_n1014), .A2(new_n1041), .A3(G390), .ZN(new_n1302));
  OAI21_X1  g1102(.A(G396), .B1(new_n1044), .B2(new_n1076), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1264), .A2(new_n1303), .ZN(new_n1304));
  AOI21_X1  g1104(.A(G390), .B1(new_n1014), .B2(new_n1041), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT126), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1264), .A2(new_n1306), .A3(new_n1303), .ZN(new_n1307));
  AOI22_X1  g1107(.A1(new_n1302), .A2(new_n1304), .B1(new_n1305), .B2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(G390), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(G387), .A2(new_n1309), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1014), .A2(G390), .A3(new_n1041), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1307), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1310), .A2(new_n1311), .A3(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1308), .A2(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1314), .ZN(new_n1315));
  AOI211_X1 g1115(.A(new_n1274), .B(new_n1290), .C1(new_n1275), .C2(new_n1279), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT125), .ZN(new_n1317));
  OAI21_X1  g1117(.A(KEYINPUT63), .B1(new_n1316), .B2(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1275), .A2(new_n1279), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1274), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1319), .A2(new_n1320), .A3(new_n1291), .ZN(new_n1321));
  INV_X1    g1121(.A(KEYINPUT63), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1321), .A2(KEYINPUT125), .A3(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1318), .A2(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1325));
  AND2_X1   g1125(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT61), .ZN(new_n1328));
  NAND4_X1  g1128(.A1(new_n1327), .A2(new_n1308), .A3(new_n1328), .A4(new_n1313), .ZN(new_n1329));
  OAI22_X1  g1129(.A1(new_n1301), .A2(new_n1315), .B1(new_n1324), .B2(new_n1329), .ZN(G405));
  NAND2_X1  g1130(.A1(G375), .A2(new_n1260), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1331), .A2(new_n1275), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1332), .A2(new_n1291), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1331), .A2(new_n1275), .A3(new_n1290), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1333), .A2(new_n1334), .ZN(new_n1335));
  XNOR2_X1  g1135(.A(new_n1314), .B(new_n1335), .ZN(G402));
endmodule


