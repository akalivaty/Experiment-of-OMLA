

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U559 ( .A(n694), .B(KEYINPUT26), .ZN(n695) );
  BUF_X1 U560 ( .A(n688), .Z(G160) );
  NOR2_X1 U561 ( .A1(n703), .A2(n702), .ZN(n697) );
  XOR2_X1 U562 ( .A(KEYINPUT70), .B(n578), .Z(n524) );
  OR2_X1 U563 ( .A1(n770), .A2(n769), .ZN(n525) );
  AND2_X1 U564 ( .A1(n979), .A2(n821), .ZN(n526) );
  NOR2_X1 U565 ( .A1(n807), .A2(n526), .ZN(n808) );
  NOR2_X1 U566 ( .A1(G651), .A2(G543), .ZN(n644) );
  XOR2_X1 U567 ( .A(n591), .B(KEYINPUT15), .Z(n984) );
  NAND2_X1 U568 ( .A1(G89), .A2(n644), .ZN(n527) );
  XOR2_X1 U569 ( .A(KEYINPUT4), .B(n527), .Z(n528) );
  XNOR2_X1 U570 ( .A(n528), .B(KEYINPUT73), .ZN(n530) );
  XOR2_X1 U571 ( .A(G543), .B(KEYINPUT0), .Z(n641) );
  INV_X1 U572 ( .A(G651), .ZN(n532) );
  NOR2_X4 U573 ( .A1(n641), .A2(n532), .ZN(n649) );
  NAND2_X1 U574 ( .A1(G76), .A2(n649), .ZN(n529) );
  NAND2_X1 U575 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U576 ( .A(KEYINPUT5), .B(n531), .ZN(n539) );
  NOR2_X1 U577 ( .A1(G543), .A2(n532), .ZN(n533) );
  XOR2_X2 U578 ( .A(KEYINPUT1), .B(n533), .Z(n646) );
  NAND2_X1 U579 ( .A1(G63), .A2(n646), .ZN(n535) );
  NOR2_X2 U580 ( .A1(G651), .A2(n641), .ZN(n655) );
  NAND2_X1 U581 ( .A1(G51), .A2(n655), .ZN(n534) );
  NAND2_X1 U582 ( .A1(n535), .A2(n534), .ZN(n537) );
  XOR2_X1 U583 ( .A(KEYINPUT6), .B(KEYINPUT74), .Z(n536) );
  XNOR2_X1 U584 ( .A(n537), .B(n536), .ZN(n538) );
  NAND2_X1 U585 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U586 ( .A(KEYINPUT7), .B(n540), .ZN(G168) );
  XOR2_X1 U587 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U588 ( .A1(G52), .A2(n655), .ZN(n541) );
  XOR2_X1 U589 ( .A(KEYINPUT68), .B(n541), .Z(n548) );
  NAND2_X1 U590 ( .A1(G77), .A2(n649), .ZN(n543) );
  NAND2_X1 U591 ( .A1(G90), .A2(n644), .ZN(n542) );
  NAND2_X1 U592 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U593 ( .A(n544), .B(KEYINPUT9), .ZN(n546) );
  NAND2_X1 U594 ( .A1(G64), .A2(n646), .ZN(n545) );
  NAND2_X1 U595 ( .A1(n546), .A2(n545), .ZN(n547) );
  NOR2_X1 U596 ( .A1(n548), .A2(n547), .ZN(G171) );
  NOR2_X1 U597 ( .A1(G2104), .A2(G2105), .ZN(n549) );
  XOR2_X2 U598 ( .A(KEYINPUT17), .B(n549), .Z(n885) );
  NAND2_X1 U599 ( .A1(G137), .A2(n885), .ZN(n560) );
  AND2_X1 U600 ( .A1(G2104), .A2(G2105), .ZN(n888) );
  NAND2_X1 U601 ( .A1(G113), .A2(n888), .ZN(n550) );
  XNOR2_X1 U602 ( .A(n550), .B(KEYINPUT66), .ZN(n554) );
  NAND2_X1 U603 ( .A1(G2104), .A2(G101), .ZN(n551) );
  OR2_X1 U604 ( .A1(G2105), .A2(n551), .ZN(n552) );
  XOR2_X1 U605 ( .A(KEYINPUT23), .B(n552), .Z(n553) );
  NAND2_X1 U606 ( .A1(n554), .A2(n553), .ZN(n558) );
  INV_X1 U607 ( .A(G2104), .ZN(n555) );
  NAND2_X1 U608 ( .A1(n555), .A2(G2105), .ZN(n556) );
  XNOR2_X2 U609 ( .A(n556), .B(KEYINPUT65), .ZN(n890) );
  AND2_X1 U610 ( .A1(G125), .A2(n890), .ZN(n557) );
  NOR2_X1 U611 ( .A1(n558), .A2(n557), .ZN(n559) );
  AND2_X1 U612 ( .A1(n560), .A2(n559), .ZN(n688) );
  AND2_X1 U613 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U614 ( .A1(G65), .A2(n646), .ZN(n563) );
  NAND2_X1 U615 ( .A1(G53), .A2(n655), .ZN(n562) );
  NAND2_X1 U616 ( .A1(n563), .A2(n562), .ZN(n567) );
  NAND2_X1 U617 ( .A1(G78), .A2(n649), .ZN(n565) );
  NAND2_X1 U618 ( .A1(G91), .A2(n644), .ZN(n564) );
  NAND2_X1 U619 ( .A1(n565), .A2(n564), .ZN(n566) );
  NOR2_X1 U620 ( .A1(n567), .A2(n566), .ZN(n973) );
  INV_X1 U621 ( .A(n973), .ZN(G299) );
  INV_X1 U622 ( .A(G132), .ZN(G219) );
  INV_X1 U623 ( .A(G82), .ZN(G220) );
  INV_X1 U624 ( .A(G120), .ZN(G236) );
  INV_X1 U625 ( .A(G69), .ZN(G235) );
  NOR2_X1 U626 ( .A1(G2105), .A2(n555), .ZN(n884) );
  NAND2_X1 U627 ( .A1(G102), .A2(n884), .ZN(n569) );
  NAND2_X1 U628 ( .A1(G138), .A2(n885), .ZN(n568) );
  NAND2_X1 U629 ( .A1(n569), .A2(n568), .ZN(n573) );
  NAND2_X1 U630 ( .A1(G126), .A2(n890), .ZN(n571) );
  NAND2_X1 U631 ( .A1(G114), .A2(n888), .ZN(n570) );
  NAND2_X1 U632 ( .A1(n571), .A2(n570), .ZN(n572) );
  NOR2_X1 U633 ( .A1(n573), .A2(n572), .ZN(G164) );
  NAND2_X1 U634 ( .A1(G7), .A2(G661), .ZN(n574) );
  XOR2_X1 U635 ( .A(n574), .B(KEYINPUT10), .Z(n921) );
  NAND2_X1 U636 ( .A1(n921), .A2(G567), .ZN(n575) );
  XOR2_X1 U637 ( .A(KEYINPUT11), .B(n575), .Z(G234) );
  NAND2_X1 U638 ( .A1(G56), .A2(n646), .ZN(n576) );
  XOR2_X1 U639 ( .A(KEYINPUT14), .B(n576), .Z(n582) );
  NAND2_X1 U640 ( .A1(n644), .A2(G81), .ZN(n577) );
  XOR2_X1 U641 ( .A(KEYINPUT12), .B(n577), .Z(n579) );
  NAND2_X1 U642 ( .A1(n649), .A2(G68), .ZN(n578) );
  NOR2_X1 U643 ( .A1(n579), .A2(n524), .ZN(n580) );
  XNOR2_X1 U644 ( .A(n580), .B(KEYINPUT13), .ZN(n581) );
  NOR2_X1 U645 ( .A1(n582), .A2(n581), .ZN(n584) );
  NAND2_X1 U646 ( .A1(n655), .A2(G43), .ZN(n583) );
  NAND2_X1 U647 ( .A1(n584), .A2(n583), .ZN(n989) );
  INV_X1 U648 ( .A(G860), .ZN(n598) );
  OR2_X1 U649 ( .A1(n989), .A2(n598), .ZN(G153) );
  NAND2_X1 U650 ( .A1(G54), .A2(n655), .ZN(n586) );
  NAND2_X1 U651 ( .A1(G92), .A2(n644), .ZN(n585) );
  NAND2_X1 U652 ( .A1(n586), .A2(n585), .ZN(n590) );
  NAND2_X1 U653 ( .A1(G66), .A2(n646), .ZN(n588) );
  NAND2_X1 U654 ( .A1(G79), .A2(n649), .ZN(n587) );
  NAND2_X1 U655 ( .A1(n588), .A2(n587), .ZN(n589) );
  NOR2_X1 U656 ( .A1(n590), .A2(n589), .ZN(n591) );
  NOR2_X1 U657 ( .A1(n984), .A2(G868), .ZN(n592) );
  XOR2_X1 U658 ( .A(KEYINPUT72), .B(n592), .Z(n595) );
  INV_X1 U659 ( .A(G868), .ZN(n668) );
  NOR2_X1 U660 ( .A1(G171), .A2(n668), .ZN(n593) );
  XNOR2_X1 U661 ( .A(KEYINPUT71), .B(n593), .ZN(n594) );
  NAND2_X1 U662 ( .A1(n595), .A2(n594), .ZN(G284) );
  NOR2_X1 U663 ( .A1(G286), .A2(n668), .ZN(n597) );
  NOR2_X1 U664 ( .A1(G868), .A2(G299), .ZN(n596) );
  NOR2_X1 U665 ( .A1(n597), .A2(n596), .ZN(G297) );
  NAND2_X1 U666 ( .A1(n598), .A2(G559), .ZN(n599) );
  NAND2_X1 U667 ( .A1(n599), .A2(n984), .ZN(n600) );
  XNOR2_X1 U668 ( .A(n600), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U669 ( .A1(G868), .A2(n989), .ZN(n603) );
  NAND2_X1 U670 ( .A1(G868), .A2(n984), .ZN(n601) );
  NOR2_X1 U671 ( .A1(G559), .A2(n601), .ZN(n602) );
  NOR2_X1 U672 ( .A1(n603), .A2(n602), .ZN(G282) );
  XOR2_X1 U673 ( .A(KEYINPUT75), .B(KEYINPUT18), .Z(n605) );
  NAND2_X1 U674 ( .A1(G123), .A2(n890), .ZN(n604) );
  XNOR2_X1 U675 ( .A(n605), .B(n604), .ZN(n612) );
  NAND2_X1 U676 ( .A1(G99), .A2(n884), .ZN(n607) );
  NAND2_X1 U677 ( .A1(G111), .A2(n888), .ZN(n606) );
  NAND2_X1 U678 ( .A1(n607), .A2(n606), .ZN(n610) );
  NAND2_X1 U679 ( .A1(n885), .A2(G135), .ZN(n608) );
  XOR2_X1 U680 ( .A(KEYINPUT76), .B(n608), .Z(n609) );
  NOR2_X1 U681 ( .A1(n610), .A2(n609), .ZN(n611) );
  NAND2_X1 U682 ( .A1(n612), .A2(n611), .ZN(n936) );
  XOR2_X1 U683 ( .A(G2096), .B(KEYINPUT77), .Z(n613) );
  XNOR2_X1 U684 ( .A(n936), .B(n613), .ZN(n614) );
  NOR2_X1 U685 ( .A1(G2100), .A2(n614), .ZN(n615) );
  XOR2_X1 U686 ( .A(KEYINPUT78), .B(n615), .Z(G156) );
  NAND2_X1 U687 ( .A1(G67), .A2(n646), .ZN(n617) );
  NAND2_X1 U688 ( .A1(G80), .A2(n649), .ZN(n616) );
  NAND2_X1 U689 ( .A1(n617), .A2(n616), .ZN(n621) );
  NAND2_X1 U690 ( .A1(G55), .A2(n655), .ZN(n619) );
  NAND2_X1 U691 ( .A1(G93), .A2(n644), .ZN(n618) );
  NAND2_X1 U692 ( .A1(n619), .A2(n618), .ZN(n620) );
  OR2_X1 U693 ( .A1(n621), .A2(n620), .ZN(n669) );
  NAND2_X1 U694 ( .A1(G559), .A2(n984), .ZN(n622) );
  XNOR2_X1 U695 ( .A(n622), .B(KEYINPUT79), .ZN(n666) );
  XOR2_X1 U696 ( .A(n666), .B(n989), .Z(n623) );
  NOR2_X1 U697 ( .A1(G860), .A2(n623), .ZN(n624) );
  XOR2_X1 U698 ( .A(n669), .B(n624), .Z(G145) );
  NAND2_X1 U699 ( .A1(G75), .A2(n649), .ZN(n626) );
  NAND2_X1 U700 ( .A1(G88), .A2(n644), .ZN(n625) );
  NAND2_X1 U701 ( .A1(n626), .A2(n625), .ZN(n630) );
  NAND2_X1 U702 ( .A1(G62), .A2(n646), .ZN(n628) );
  NAND2_X1 U703 ( .A1(G50), .A2(n655), .ZN(n627) );
  NAND2_X1 U704 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U705 ( .A1(n630), .A2(n629), .ZN(G166) );
  INV_X1 U706 ( .A(G166), .ZN(G303) );
  NAND2_X1 U707 ( .A1(G60), .A2(n646), .ZN(n632) );
  NAND2_X1 U708 ( .A1(G47), .A2(n655), .ZN(n631) );
  NAND2_X1 U709 ( .A1(n632), .A2(n631), .ZN(n633) );
  XNOR2_X1 U710 ( .A(KEYINPUT67), .B(n633), .ZN(n637) );
  NAND2_X1 U711 ( .A1(G72), .A2(n649), .ZN(n635) );
  NAND2_X1 U712 ( .A1(G85), .A2(n644), .ZN(n634) );
  AND2_X1 U713 ( .A1(n635), .A2(n634), .ZN(n636) );
  NAND2_X1 U714 ( .A1(n637), .A2(n636), .ZN(G290) );
  NAND2_X1 U715 ( .A1(G49), .A2(n655), .ZN(n639) );
  NAND2_X1 U716 ( .A1(G74), .A2(G651), .ZN(n638) );
  NAND2_X1 U717 ( .A1(n639), .A2(n638), .ZN(n640) );
  NOR2_X1 U718 ( .A1(n646), .A2(n640), .ZN(n643) );
  NAND2_X1 U719 ( .A1(n641), .A2(G87), .ZN(n642) );
  NAND2_X1 U720 ( .A1(n643), .A2(n642), .ZN(G288) );
  NAND2_X1 U721 ( .A1(n644), .A2(G86), .ZN(n645) );
  XNOR2_X1 U722 ( .A(n645), .B(KEYINPUT80), .ZN(n648) );
  NAND2_X1 U723 ( .A1(G61), .A2(n646), .ZN(n647) );
  NAND2_X1 U724 ( .A1(n648), .A2(n647), .ZN(n653) );
  NAND2_X1 U725 ( .A1(G73), .A2(n649), .ZN(n650) );
  XNOR2_X1 U726 ( .A(n650), .B(KEYINPUT2), .ZN(n651) );
  XNOR2_X1 U727 ( .A(n651), .B(KEYINPUT81), .ZN(n652) );
  NOR2_X1 U728 ( .A1(n653), .A2(n652), .ZN(n654) );
  XNOR2_X1 U729 ( .A(n654), .B(KEYINPUT82), .ZN(n657) );
  NAND2_X1 U730 ( .A1(G48), .A2(n655), .ZN(n656) );
  NAND2_X1 U731 ( .A1(n657), .A2(n656), .ZN(G305) );
  XOR2_X1 U732 ( .A(KEYINPUT19), .B(KEYINPUT83), .Z(n659) );
  XOR2_X1 U733 ( .A(G303), .B(KEYINPUT84), .Z(n658) );
  XNOR2_X1 U734 ( .A(n659), .B(n658), .ZN(n662) );
  XOR2_X1 U735 ( .A(G299), .B(G290), .Z(n660) );
  XNOR2_X1 U736 ( .A(n660), .B(G288), .ZN(n661) );
  XNOR2_X1 U737 ( .A(n662), .B(n661), .ZN(n664) );
  XOR2_X1 U738 ( .A(G305), .B(n669), .Z(n663) );
  XNOR2_X1 U739 ( .A(n664), .B(n663), .ZN(n665) );
  XOR2_X1 U740 ( .A(n665), .B(n989), .Z(n900) );
  XNOR2_X1 U741 ( .A(n666), .B(n900), .ZN(n667) );
  NOR2_X1 U742 ( .A1(n668), .A2(n667), .ZN(n671) );
  NOR2_X1 U743 ( .A1(G868), .A2(n669), .ZN(n670) );
  NOR2_X1 U744 ( .A1(n671), .A2(n670), .ZN(G295) );
  XOR2_X1 U745 ( .A(KEYINPUT21), .B(KEYINPUT85), .Z(n675) );
  NAND2_X1 U746 ( .A1(G2078), .A2(G2084), .ZN(n672) );
  XOR2_X1 U747 ( .A(KEYINPUT20), .B(n672), .Z(n673) );
  NAND2_X1 U748 ( .A1(n673), .A2(G2090), .ZN(n674) );
  XNOR2_X1 U749 ( .A(n675), .B(n674), .ZN(n676) );
  NAND2_X1 U750 ( .A1(n676), .A2(G2072), .ZN(n677) );
  XNOR2_X1 U751 ( .A(n677), .B(KEYINPUT86), .ZN(G158) );
  XNOR2_X1 U752 ( .A(KEYINPUT69), .B(G57), .ZN(G237) );
  XOR2_X1 U753 ( .A(KEYINPUT87), .B(G44), .Z(n678) );
  XNOR2_X1 U754 ( .A(KEYINPUT3), .B(n678), .ZN(G218) );
  NOR2_X1 U755 ( .A1(G235), .A2(G236), .ZN(n679) );
  XOR2_X1 U756 ( .A(KEYINPUT88), .B(n679), .Z(n680) );
  NOR2_X1 U757 ( .A1(G237), .A2(n680), .ZN(n681) );
  NAND2_X1 U758 ( .A1(G108), .A2(n681), .ZN(n829) );
  NAND2_X1 U759 ( .A1(n829), .A2(G567), .ZN(n686) );
  NOR2_X1 U760 ( .A1(G220), .A2(G219), .ZN(n682) );
  XOR2_X1 U761 ( .A(KEYINPUT22), .B(n682), .Z(n683) );
  NOR2_X1 U762 ( .A1(G218), .A2(n683), .ZN(n684) );
  NAND2_X1 U763 ( .A1(G96), .A2(n684), .ZN(n830) );
  NAND2_X1 U764 ( .A1(n830), .A2(G2106), .ZN(n685) );
  NAND2_X1 U765 ( .A1(n686), .A2(n685), .ZN(n831) );
  NAND2_X1 U766 ( .A1(G661), .A2(G483), .ZN(n687) );
  NOR2_X1 U767 ( .A1(n831), .A2(n687), .ZN(n828) );
  NAND2_X1 U768 ( .A1(n828), .A2(G36), .ZN(G176) );
  NOR2_X1 U769 ( .A1(G164), .A2(G1384), .ZN(n772) );
  NAND2_X1 U770 ( .A1(n688), .A2(G40), .ZN(n771) );
  INV_X1 U771 ( .A(KEYINPUT98), .ZN(n689) );
  XNOR2_X1 U772 ( .A(n771), .B(n689), .ZN(n690) );
  NAND2_X2 U773 ( .A1(n772), .A2(n690), .ZN(n732) );
  NAND2_X1 U774 ( .A1(G8), .A2(n732), .ZN(n767) );
  NOR2_X1 U775 ( .A1(G1976), .A2(G288), .ZN(n750) );
  NAND2_X1 U776 ( .A1(n750), .A2(KEYINPUT33), .ZN(n691) );
  NOR2_X1 U777 ( .A1(n767), .A2(n691), .ZN(n757) );
  AND2_X1 U778 ( .A1(G1341), .A2(n732), .ZN(n692) );
  NOR2_X1 U779 ( .A1(n692), .A2(n989), .ZN(n696) );
  INV_X1 U780 ( .A(n732), .ZN(n693) );
  NAND2_X1 U781 ( .A1(n693), .A2(G1996), .ZN(n694) );
  NAND2_X1 U782 ( .A1(n696), .A2(n695), .ZN(n703) );
  INV_X1 U783 ( .A(n984), .ZN(n702) );
  XNOR2_X1 U784 ( .A(n697), .B(KEYINPUT101), .ZN(n701) );
  INV_X1 U785 ( .A(n732), .ZN(n718) );
  NOR2_X1 U786 ( .A1(n718), .A2(G1348), .ZN(n699) );
  NOR2_X1 U787 ( .A1(G2067), .A2(n732), .ZN(n698) );
  NOR2_X1 U788 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U789 ( .A1(n701), .A2(n700), .ZN(n705) );
  NAND2_X1 U790 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U791 ( .A1(n705), .A2(n704), .ZN(n711) );
  NAND2_X1 U792 ( .A1(n718), .A2(G2072), .ZN(n706) );
  XNOR2_X1 U793 ( .A(KEYINPUT27), .B(n706), .ZN(n709) );
  NAND2_X1 U794 ( .A1(G1956), .A2(n732), .ZN(n707) );
  XOR2_X1 U795 ( .A(KEYINPUT100), .B(n707), .Z(n708) );
  NOR2_X1 U796 ( .A1(n709), .A2(n708), .ZN(n712) );
  NAND2_X1 U797 ( .A1(n973), .A2(n712), .ZN(n710) );
  NAND2_X1 U798 ( .A1(n711), .A2(n710), .ZN(n715) );
  NOR2_X1 U799 ( .A1(n973), .A2(n712), .ZN(n713) );
  XOR2_X1 U800 ( .A(n713), .B(KEYINPUT28), .Z(n714) );
  NAND2_X1 U801 ( .A1(n715), .A2(n714), .ZN(n717) );
  XOR2_X1 U802 ( .A(KEYINPUT29), .B(KEYINPUT102), .Z(n716) );
  XNOR2_X1 U803 ( .A(n717), .B(n716), .ZN(n722) );
  INV_X1 U804 ( .A(G1961), .ZN(n832) );
  NAND2_X1 U805 ( .A1(n732), .A2(n832), .ZN(n720) );
  XNOR2_X1 U806 ( .A(KEYINPUT25), .B(G2078), .ZN(n950) );
  NAND2_X1 U807 ( .A1(n718), .A2(n950), .ZN(n719) );
  NAND2_X1 U808 ( .A1(n720), .A2(n719), .ZN(n726) );
  NAND2_X1 U809 ( .A1(n726), .A2(G171), .ZN(n721) );
  NAND2_X1 U810 ( .A1(n722), .A2(n721), .ZN(n731) );
  NOR2_X1 U811 ( .A1(G1966), .A2(n767), .ZN(n744) );
  NOR2_X1 U812 ( .A1(G2084), .A2(n732), .ZN(n741) );
  NOR2_X1 U813 ( .A1(n744), .A2(n741), .ZN(n723) );
  NAND2_X1 U814 ( .A1(G8), .A2(n723), .ZN(n724) );
  XNOR2_X1 U815 ( .A(KEYINPUT30), .B(n724), .ZN(n725) );
  NOR2_X1 U816 ( .A1(G168), .A2(n725), .ZN(n728) );
  NOR2_X1 U817 ( .A1(G171), .A2(n726), .ZN(n727) );
  NOR2_X1 U818 ( .A1(n728), .A2(n727), .ZN(n729) );
  XOR2_X1 U819 ( .A(KEYINPUT31), .B(n729), .Z(n730) );
  NAND2_X1 U820 ( .A1(n731), .A2(n730), .ZN(n742) );
  NAND2_X1 U821 ( .A1(n742), .A2(G286), .ZN(n738) );
  NOR2_X1 U822 ( .A1(G1971), .A2(n767), .ZN(n734) );
  NOR2_X1 U823 ( .A1(G2090), .A2(n732), .ZN(n733) );
  NOR2_X1 U824 ( .A1(n734), .A2(n733), .ZN(n735) );
  XOR2_X1 U825 ( .A(KEYINPUT103), .B(n735), .Z(n736) );
  NAND2_X1 U826 ( .A1(n736), .A2(G303), .ZN(n737) );
  NAND2_X1 U827 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U828 ( .A1(n739), .A2(G8), .ZN(n740) );
  XNOR2_X1 U829 ( .A(n740), .B(KEYINPUT32), .ZN(n748) );
  NAND2_X1 U830 ( .A1(G8), .A2(n741), .ZN(n746) );
  INV_X1 U831 ( .A(n742), .ZN(n743) );
  NOR2_X1 U832 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U833 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U834 ( .A1(n748), .A2(n747), .ZN(n761) );
  NOR2_X1 U835 ( .A1(G1971), .A2(G303), .ZN(n749) );
  NOR2_X1 U836 ( .A1(n750), .A2(n749), .ZN(n977) );
  NAND2_X1 U837 ( .A1(n761), .A2(n977), .ZN(n751) );
  NAND2_X1 U838 ( .A1(G1976), .A2(G288), .ZN(n972) );
  NAND2_X1 U839 ( .A1(n751), .A2(n972), .ZN(n752) );
  XNOR2_X1 U840 ( .A(KEYINPUT104), .B(n752), .ZN(n753) );
  NOR2_X1 U841 ( .A1(n767), .A2(n753), .ZN(n754) );
  XNOR2_X1 U842 ( .A(n754), .B(KEYINPUT64), .ZN(n755) );
  NOR2_X1 U843 ( .A1(KEYINPUT33), .A2(n755), .ZN(n756) );
  NOR2_X1 U844 ( .A1(n757), .A2(n756), .ZN(n758) );
  XOR2_X1 U845 ( .A(G1981), .B(G305), .Z(n980) );
  NAND2_X1 U846 ( .A1(n758), .A2(n980), .ZN(n764) );
  NOR2_X1 U847 ( .A1(G2090), .A2(G303), .ZN(n759) );
  NAND2_X1 U848 ( .A1(G8), .A2(n759), .ZN(n760) );
  NAND2_X1 U849 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U850 ( .A1(n762), .A2(n767), .ZN(n763) );
  NAND2_X1 U851 ( .A1(n764), .A2(n763), .ZN(n770) );
  NOR2_X1 U852 ( .A1(G1981), .A2(G305), .ZN(n765) );
  XNOR2_X1 U853 ( .A(n765), .B(KEYINPUT99), .ZN(n766) );
  XNOR2_X1 U854 ( .A(n766), .B(KEYINPUT24), .ZN(n768) );
  NOR2_X1 U855 ( .A1(n768), .A2(n767), .ZN(n769) );
  NOR2_X1 U856 ( .A1(n772), .A2(n771), .ZN(n821) );
  NAND2_X1 U857 ( .A1(G104), .A2(n884), .ZN(n774) );
  NAND2_X1 U858 ( .A1(G140), .A2(n885), .ZN(n773) );
  NAND2_X1 U859 ( .A1(n774), .A2(n773), .ZN(n775) );
  XNOR2_X1 U860 ( .A(KEYINPUT34), .B(n775), .ZN(n783) );
  NAND2_X1 U861 ( .A1(G128), .A2(n890), .ZN(n778) );
  NAND2_X1 U862 ( .A1(n888), .A2(G116), .ZN(n776) );
  XOR2_X1 U863 ( .A(KEYINPUT89), .B(n776), .Z(n777) );
  NAND2_X1 U864 ( .A1(n778), .A2(n777), .ZN(n781) );
  XNOR2_X1 U865 ( .A(KEYINPUT90), .B(KEYINPUT91), .ZN(n779) );
  XNOR2_X1 U866 ( .A(n779), .B(KEYINPUT35), .ZN(n780) );
  XNOR2_X1 U867 ( .A(n781), .B(n780), .ZN(n782) );
  NOR2_X1 U868 ( .A1(n783), .A2(n782), .ZN(n784) );
  XNOR2_X1 U869 ( .A(n784), .B(KEYINPUT36), .ZN(n876) );
  XNOR2_X1 U870 ( .A(G2067), .B(KEYINPUT37), .ZN(n819) );
  NOR2_X1 U871 ( .A1(n876), .A2(n819), .ZN(n785) );
  XNOR2_X1 U872 ( .A(n785), .B(KEYINPUT92), .ZN(n939) );
  NAND2_X1 U873 ( .A1(n821), .A2(n939), .ZN(n817) );
  NAND2_X1 U874 ( .A1(G131), .A2(n885), .ZN(n787) );
  NAND2_X1 U875 ( .A1(G107), .A2(n888), .ZN(n786) );
  NAND2_X1 U876 ( .A1(n787), .A2(n786), .ZN(n793) );
  NAND2_X1 U877 ( .A1(G95), .A2(n884), .ZN(n788) );
  XNOR2_X1 U878 ( .A(n788), .B(KEYINPUT94), .ZN(n791) );
  NAND2_X1 U879 ( .A1(G119), .A2(n890), .ZN(n789) );
  XOR2_X1 U880 ( .A(KEYINPUT93), .B(n789), .Z(n790) );
  NAND2_X1 U881 ( .A1(n791), .A2(n790), .ZN(n792) );
  NOR2_X1 U882 ( .A1(n793), .A2(n792), .ZN(n877) );
  INV_X1 U883 ( .A(G1991), .ZN(n835) );
  NOR2_X1 U884 ( .A1(n877), .A2(n835), .ZN(n804) );
  XOR2_X1 U885 ( .A(KEYINPUT95), .B(KEYINPUT38), .Z(n795) );
  NAND2_X1 U886 ( .A1(G105), .A2(n884), .ZN(n794) );
  XNOR2_X1 U887 ( .A(n795), .B(n794), .ZN(n802) );
  NAND2_X1 U888 ( .A1(G129), .A2(n890), .ZN(n797) );
  NAND2_X1 U889 ( .A1(G117), .A2(n888), .ZN(n796) );
  NAND2_X1 U890 ( .A1(n797), .A2(n796), .ZN(n800) );
  NAND2_X1 U891 ( .A1(n885), .A2(G141), .ZN(n798) );
  XOR2_X1 U892 ( .A(KEYINPUT96), .B(n798), .Z(n799) );
  NOR2_X1 U893 ( .A1(n800), .A2(n799), .ZN(n801) );
  NAND2_X1 U894 ( .A1(n802), .A2(n801), .ZN(n878) );
  AND2_X1 U895 ( .A1(n878), .A2(G1996), .ZN(n803) );
  NOR2_X1 U896 ( .A1(n804), .A2(n803), .ZN(n923) );
  INV_X1 U897 ( .A(n923), .ZN(n805) );
  NAND2_X1 U898 ( .A1(n805), .A2(n821), .ZN(n809) );
  NAND2_X1 U899 ( .A1(n817), .A2(n809), .ZN(n806) );
  XOR2_X1 U900 ( .A(KEYINPUT97), .B(n806), .Z(n807) );
  XNOR2_X1 U901 ( .A(G1986), .B(G290), .ZN(n979) );
  NAND2_X1 U902 ( .A1(n525), .A2(n808), .ZN(n824) );
  NOR2_X1 U903 ( .A1(G1996), .A2(n878), .ZN(n929) );
  INV_X1 U904 ( .A(n809), .ZN(n813) );
  NOR2_X1 U905 ( .A1(G1986), .A2(G290), .ZN(n811) );
  AND2_X1 U906 ( .A1(n835), .A2(n877), .ZN(n810) );
  XOR2_X1 U907 ( .A(KEYINPUT105), .B(n810), .Z(n935) );
  NOR2_X1 U908 ( .A1(n811), .A2(n935), .ZN(n812) );
  NOR2_X1 U909 ( .A1(n813), .A2(n812), .ZN(n814) );
  XNOR2_X1 U910 ( .A(n814), .B(KEYINPUT106), .ZN(n815) );
  NOR2_X1 U911 ( .A1(n929), .A2(n815), .ZN(n816) );
  XNOR2_X1 U912 ( .A(n816), .B(KEYINPUT39), .ZN(n818) );
  NAND2_X1 U913 ( .A1(n818), .A2(n817), .ZN(n820) );
  NAND2_X1 U914 ( .A1(n819), .A2(n876), .ZN(n922) );
  NAND2_X1 U915 ( .A1(n820), .A2(n922), .ZN(n822) );
  NAND2_X1 U916 ( .A1(n822), .A2(n821), .ZN(n823) );
  NAND2_X1 U917 ( .A1(n824), .A2(n823), .ZN(n825) );
  XNOR2_X1 U918 ( .A(KEYINPUT40), .B(n825), .ZN(G329) );
  NAND2_X1 U919 ( .A1(G2106), .A2(n921), .ZN(G217) );
  AND2_X1 U920 ( .A1(G15), .A2(G2), .ZN(n826) );
  NAND2_X1 U921 ( .A1(G661), .A2(n826), .ZN(G259) );
  NAND2_X1 U922 ( .A1(G3), .A2(G1), .ZN(n827) );
  NAND2_X1 U923 ( .A1(n828), .A2(n827), .ZN(G188) );
  INV_X1 U925 ( .A(G108), .ZN(G238) );
  INV_X1 U926 ( .A(G96), .ZN(G221) );
  NOR2_X1 U927 ( .A1(n830), .A2(n829), .ZN(G325) );
  INV_X1 U928 ( .A(G325), .ZN(G261) );
  INV_X1 U929 ( .A(n831), .ZN(G319) );
  XNOR2_X1 U930 ( .A(G1981), .B(G2474), .ZN(n843) );
  XNOR2_X1 U931 ( .A(G1956), .B(n832), .ZN(n834) );
  XNOR2_X1 U932 ( .A(G1986), .B(G1966), .ZN(n833) );
  XNOR2_X1 U933 ( .A(n834), .B(n833), .ZN(n839) );
  XOR2_X1 U934 ( .A(G1976), .B(G1971), .Z(n837) );
  XOR2_X1 U935 ( .A(G1996), .B(n835), .Z(n836) );
  XNOR2_X1 U936 ( .A(n837), .B(n836), .ZN(n838) );
  XOR2_X1 U937 ( .A(n839), .B(n838), .Z(n841) );
  XNOR2_X1 U938 ( .A(KEYINPUT112), .B(KEYINPUT41), .ZN(n840) );
  XNOR2_X1 U939 ( .A(n841), .B(n840), .ZN(n842) );
  XNOR2_X1 U940 ( .A(n843), .B(n842), .ZN(G229) );
  XNOR2_X1 U941 ( .A(G2078), .B(G2072), .ZN(n844) );
  XNOR2_X1 U942 ( .A(n844), .B(KEYINPUT110), .ZN(n854) );
  XOR2_X1 U943 ( .A(KEYINPUT111), .B(G2678), .Z(n846) );
  XNOR2_X1 U944 ( .A(KEYINPUT43), .B(G2096), .ZN(n845) );
  XNOR2_X1 U945 ( .A(n846), .B(n845), .ZN(n850) );
  XOR2_X1 U946 ( .A(G2100), .B(G2090), .Z(n848) );
  XNOR2_X1 U947 ( .A(G2067), .B(G2084), .ZN(n847) );
  XNOR2_X1 U948 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U949 ( .A(n850), .B(n849), .Z(n852) );
  XNOR2_X1 U950 ( .A(KEYINPUT109), .B(KEYINPUT42), .ZN(n851) );
  XNOR2_X1 U951 ( .A(n852), .B(n851), .ZN(n853) );
  XNOR2_X1 U952 ( .A(n854), .B(n853), .ZN(G227) );
  NAND2_X1 U953 ( .A1(G100), .A2(n884), .ZN(n856) );
  NAND2_X1 U954 ( .A1(G112), .A2(n888), .ZN(n855) );
  NAND2_X1 U955 ( .A1(n856), .A2(n855), .ZN(n862) );
  NAND2_X1 U956 ( .A1(n890), .A2(G124), .ZN(n857) );
  XNOR2_X1 U957 ( .A(n857), .B(KEYINPUT44), .ZN(n859) );
  NAND2_X1 U958 ( .A1(G136), .A2(n885), .ZN(n858) );
  NAND2_X1 U959 ( .A1(n859), .A2(n858), .ZN(n860) );
  XOR2_X1 U960 ( .A(KEYINPUT113), .B(n860), .Z(n861) );
  NOR2_X1 U961 ( .A1(n862), .A2(n861), .ZN(G162) );
  NAND2_X1 U962 ( .A1(G130), .A2(n890), .ZN(n864) );
  NAND2_X1 U963 ( .A1(G118), .A2(n888), .ZN(n863) );
  NAND2_X1 U964 ( .A1(n864), .A2(n863), .ZN(n870) );
  NAND2_X1 U965 ( .A1(G106), .A2(n884), .ZN(n866) );
  NAND2_X1 U966 ( .A1(G142), .A2(n885), .ZN(n865) );
  NAND2_X1 U967 ( .A1(n866), .A2(n865), .ZN(n867) );
  XOR2_X1 U968 ( .A(KEYINPUT114), .B(n867), .Z(n868) );
  XNOR2_X1 U969 ( .A(KEYINPUT45), .B(n868), .ZN(n869) );
  NOR2_X1 U970 ( .A1(n870), .A2(n869), .ZN(n874) );
  XOR2_X1 U971 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n872) );
  XNOR2_X1 U972 ( .A(KEYINPUT118), .B(KEYINPUT115), .ZN(n871) );
  XNOR2_X1 U973 ( .A(n872), .B(n871), .ZN(n873) );
  XOR2_X1 U974 ( .A(n874), .B(n873), .Z(n875) );
  XNOR2_X1 U975 ( .A(n876), .B(n875), .ZN(n881) );
  XNOR2_X1 U976 ( .A(n878), .B(n877), .ZN(n879) );
  XNOR2_X1 U977 ( .A(n879), .B(n936), .ZN(n880) );
  XOR2_X1 U978 ( .A(n881), .B(n880), .Z(n883) );
  XNOR2_X1 U979 ( .A(G164), .B(G160), .ZN(n882) );
  XNOR2_X1 U980 ( .A(n883), .B(n882), .ZN(n898) );
  NAND2_X1 U981 ( .A1(G103), .A2(n884), .ZN(n887) );
  NAND2_X1 U982 ( .A1(G139), .A2(n885), .ZN(n886) );
  NAND2_X1 U983 ( .A1(n887), .A2(n886), .ZN(n896) );
  NAND2_X1 U984 ( .A1(n888), .A2(G115), .ZN(n889) );
  XNOR2_X1 U985 ( .A(KEYINPUT117), .B(n889), .ZN(n893) );
  NAND2_X1 U986 ( .A1(n890), .A2(G127), .ZN(n891) );
  XOR2_X1 U987 ( .A(KEYINPUT116), .B(n891), .Z(n892) );
  NOR2_X1 U988 ( .A1(n893), .A2(n892), .ZN(n894) );
  XNOR2_X1 U989 ( .A(n894), .B(KEYINPUT47), .ZN(n895) );
  NOR2_X1 U990 ( .A1(n896), .A2(n895), .ZN(n924) );
  XNOR2_X1 U991 ( .A(n924), .B(G162), .ZN(n897) );
  XNOR2_X1 U992 ( .A(n898), .B(n897), .ZN(n899) );
  NOR2_X1 U993 ( .A1(G37), .A2(n899), .ZN(G395) );
  XOR2_X1 U994 ( .A(G286), .B(n984), .Z(n901) );
  XNOR2_X1 U995 ( .A(n901), .B(n900), .ZN(n902) );
  XOR2_X1 U996 ( .A(n902), .B(G171), .Z(n903) );
  NOR2_X1 U997 ( .A1(G37), .A2(n903), .ZN(G397) );
  XNOR2_X1 U998 ( .A(G2451), .B(G2446), .ZN(n913) );
  XOR2_X1 U999 ( .A(G2430), .B(KEYINPUT108), .Z(n905) );
  XNOR2_X1 U1000 ( .A(G2454), .B(G2435), .ZN(n904) );
  XNOR2_X1 U1001 ( .A(n905), .B(n904), .ZN(n909) );
  XOR2_X1 U1002 ( .A(G2438), .B(KEYINPUT107), .Z(n907) );
  XNOR2_X1 U1003 ( .A(G1341), .B(G1348), .ZN(n906) );
  XNOR2_X1 U1004 ( .A(n907), .B(n906), .ZN(n908) );
  XOR2_X1 U1005 ( .A(n909), .B(n908), .Z(n911) );
  XNOR2_X1 U1006 ( .A(G2443), .B(G2427), .ZN(n910) );
  XNOR2_X1 U1007 ( .A(n911), .B(n910), .ZN(n912) );
  XNOR2_X1 U1008 ( .A(n913), .B(n912), .ZN(n914) );
  NAND2_X1 U1009 ( .A1(n914), .A2(G14), .ZN(n920) );
  NAND2_X1 U1010 ( .A1(G319), .A2(n920), .ZN(n917) );
  NOR2_X1 U1011 ( .A1(G229), .A2(G227), .ZN(n915) );
  XNOR2_X1 U1012 ( .A(KEYINPUT49), .B(n915), .ZN(n916) );
  NOR2_X1 U1013 ( .A1(n917), .A2(n916), .ZN(n919) );
  NOR2_X1 U1014 ( .A1(G395), .A2(G397), .ZN(n918) );
  NAND2_X1 U1015 ( .A1(n919), .A2(n918), .ZN(G225) );
  INV_X1 U1016 ( .A(G225), .ZN(G308) );
  INV_X1 U1017 ( .A(n920), .ZN(G401) );
  INV_X1 U1018 ( .A(n921), .ZN(G223) );
  NAND2_X1 U1019 ( .A1(n923), .A2(n922), .ZN(n944) );
  XOR2_X1 U1020 ( .A(G2072), .B(n924), .Z(n926) );
  XOR2_X1 U1021 ( .A(G164), .B(G2078), .Z(n925) );
  NOR2_X1 U1022 ( .A1(n926), .A2(n925), .ZN(n927) );
  XOR2_X1 U1023 ( .A(KEYINPUT50), .B(n927), .Z(n933) );
  XOR2_X1 U1024 ( .A(G2090), .B(G162), .Z(n928) );
  NOR2_X1 U1025 ( .A1(n929), .A2(n928), .ZN(n930) );
  XOR2_X1 U1026 ( .A(KEYINPUT51), .B(n930), .Z(n931) );
  XOR2_X1 U1027 ( .A(KEYINPUT120), .B(n931), .Z(n932) );
  NOR2_X1 U1028 ( .A1(n933), .A2(n932), .ZN(n942) );
  XOR2_X1 U1029 ( .A(G160), .B(G2084), .Z(n934) );
  NOR2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(n937) );
  NAND2_X1 U1031 ( .A1(n937), .A2(n936), .ZN(n938) );
  NOR2_X1 U1032 ( .A1(n939), .A2(n938), .ZN(n940) );
  XOR2_X1 U1033 ( .A(KEYINPUT119), .B(n940), .Z(n941) );
  NAND2_X1 U1034 ( .A1(n942), .A2(n941), .ZN(n943) );
  NOR2_X1 U1035 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1036 ( .A(KEYINPUT52), .B(n945), .ZN(n946) );
  XNOR2_X1 U1037 ( .A(KEYINPUT55), .B(KEYINPUT121), .ZN(n967) );
  NAND2_X1 U1038 ( .A1(n946), .A2(n967), .ZN(n947) );
  NAND2_X1 U1039 ( .A1(n947), .A2(G29), .ZN(n1025) );
  XNOR2_X1 U1040 ( .A(G2090), .B(G35), .ZN(n962) );
  XOR2_X1 U1041 ( .A(G25), .B(G1991), .Z(n948) );
  NAND2_X1 U1042 ( .A1(n948), .A2(G28), .ZN(n949) );
  XNOR2_X1 U1043 ( .A(KEYINPUT122), .B(n949), .ZN(n959) );
  XNOR2_X1 U1044 ( .A(G27), .B(n950), .ZN(n954) );
  XNOR2_X1 U1045 ( .A(G2067), .B(G26), .ZN(n952) );
  XNOR2_X1 U1046 ( .A(G1996), .B(G32), .ZN(n951) );
  NOR2_X1 U1047 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1048 ( .A1(n954), .A2(n953), .ZN(n956) );
  XNOR2_X1 U1049 ( .A(G33), .B(G2072), .ZN(n955) );
  NOR2_X1 U1050 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1051 ( .A(n957), .B(KEYINPUT123), .ZN(n958) );
  NOR2_X1 U1052 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1053 ( .A(KEYINPUT53), .B(n960), .ZN(n961) );
  NOR2_X1 U1054 ( .A1(n962), .A2(n961), .ZN(n965) );
  XOR2_X1 U1055 ( .A(G2084), .B(G34), .Z(n963) );
  XNOR2_X1 U1056 ( .A(KEYINPUT54), .B(n963), .ZN(n964) );
  NAND2_X1 U1057 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1058 ( .A(n967), .B(n966), .ZN(n969) );
  INV_X1 U1059 ( .A(G29), .ZN(n968) );
  NAND2_X1 U1060 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1061 ( .A1(G11), .A2(n970), .ZN(n1023) );
  INV_X1 U1062 ( .A(G16), .ZN(n1019) );
  XOR2_X1 U1063 ( .A(n1019), .B(KEYINPUT56), .Z(n995) );
  NAND2_X1 U1064 ( .A1(G1971), .A2(G303), .ZN(n971) );
  NAND2_X1 U1065 ( .A1(n972), .A2(n971), .ZN(n975) );
  XOR2_X1 U1066 ( .A(G1956), .B(n973), .Z(n974) );
  NOR2_X1 U1067 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1068 ( .A1(n977), .A2(n976), .ZN(n978) );
  NOR2_X1 U1069 ( .A1(n979), .A2(n978), .ZN(n993) );
  XNOR2_X1 U1070 ( .A(G1966), .B(G168), .ZN(n981) );
  NAND2_X1 U1071 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1072 ( .A(n982), .B(KEYINPUT124), .ZN(n983) );
  XNOR2_X1 U1073 ( .A(KEYINPUT57), .B(n983), .ZN(n988) );
  XOR2_X1 U1074 ( .A(G171), .B(G1961), .Z(n986) );
  XOR2_X1 U1075 ( .A(n984), .B(G1348), .Z(n985) );
  NOR2_X1 U1076 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1077 ( .A1(n988), .A2(n987), .ZN(n991) );
  XNOR2_X1 U1078 ( .A(G1341), .B(n989), .ZN(n990) );
  NOR2_X1 U1079 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1080 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1081 ( .A1(n995), .A2(n994), .ZN(n1021) );
  XOR2_X1 U1082 ( .A(G5), .B(G1961), .Z(n1008) );
  XNOR2_X1 U1083 ( .A(G1348), .B(KEYINPUT59), .ZN(n996) );
  XNOR2_X1 U1084 ( .A(n996), .B(G4), .ZN(n1000) );
  XNOR2_X1 U1085 ( .A(G1341), .B(G19), .ZN(n998) );
  XNOR2_X1 U1086 ( .A(G6), .B(G1981), .ZN(n997) );
  NOR2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1088 ( .A1(n1000), .A2(n999), .ZN(n1003) );
  XOR2_X1 U1089 ( .A(KEYINPUT125), .B(G1956), .Z(n1001) );
  XNOR2_X1 U1090 ( .A(G20), .B(n1001), .ZN(n1002) );
  NOR2_X1 U1091 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XOR2_X1 U1092 ( .A(KEYINPUT60), .B(n1004), .Z(n1006) );
  XNOR2_X1 U1093 ( .A(G1966), .B(G21), .ZN(n1005) );
  NOR2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1095 ( .A1(n1008), .A2(n1007), .ZN(n1016) );
  XNOR2_X1 U1096 ( .A(G1986), .B(G24), .ZN(n1010) );
  XNOR2_X1 U1097 ( .A(G23), .B(G1976), .ZN(n1009) );
  NOR2_X1 U1098 ( .A1(n1010), .A2(n1009), .ZN(n1013) );
  XOR2_X1 U1099 ( .A(G1971), .B(KEYINPUT126), .Z(n1011) );
  XNOR2_X1 U1100 ( .A(G22), .B(n1011), .ZN(n1012) );
  NAND2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1102 ( .A(KEYINPUT58), .B(n1014), .ZN(n1015) );
  NOR2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1104 ( .A(KEYINPUT61), .B(n1017), .ZN(n1018) );
  NAND2_X1 U1105 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1106 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NOR2_X1 U1107 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1108 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XNOR2_X1 U1109 ( .A(n1026), .B(KEYINPUT62), .ZN(n1027) );
  XOR2_X1 U1110 ( .A(KEYINPUT127), .B(n1027), .Z(G150) );
  INV_X1 U1111 ( .A(G150), .ZN(G311) );
  INV_X1 U1112 ( .A(G171), .ZN(G301) );
endmodule

