//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 0 0 1 1 1 0 1 1 1 0 0 1 1 0 1 0 1 0 0 0 0 0 1 0 0 0 1 1 1 0 1 0 1 1 0 0 1 1 1 1 1 0 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:26 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1290, new_n1291, new_n1292;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NOR2_X1   g0002(.A1(G58), .A2(G68), .ZN(new_n203));
  INV_X1    g0003(.A(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(G50), .ZN(new_n205));
  XNOR2_X1  g0005(.A(KEYINPUT64), .B(G20), .ZN(new_n206));
  NAND2_X1  g0006(.A1(G1), .A2(G13), .ZN(new_n207));
  NOR3_X1   g0007(.A1(new_n205), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G97), .A2(G257), .ZN(new_n210));
  INV_X1    g0010(.A(G68), .ZN(new_n211));
  INV_X1    g0011(.A(G238), .ZN(new_n212));
  OAI21_X1  g0012(.A(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n214));
  XOR2_X1   g0014(.A(new_n214), .B(KEYINPUT65), .Z(new_n215));
  AOI211_X1 g0015(.A(new_n213), .B(new_n215), .C1(G77), .C2(G244), .ZN(new_n216));
  INV_X1    g0016(.A(G58), .ZN(new_n217));
  INV_X1    g0017(.A(G232), .ZN(new_n218));
  INV_X1    g0018(.A(G87), .ZN(new_n219));
  INV_X1    g0019(.A(G250), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  AND2_X1   g0021(.A1(G107), .A2(G264), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n209), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT1), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n209), .A2(G13), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n225), .B(G250), .C1(G257), .C2(G264), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n226), .A2(KEYINPUT0), .ZN(new_n227));
  OR2_X1    g0027(.A1(new_n226), .A2(KEYINPUT0), .ZN(new_n228));
  AOI211_X1 g0028(.A(new_n208), .B(new_n224), .C1(new_n227), .C2(new_n228), .ZN(G361));
  XNOR2_X1  g0029(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G244), .ZN(new_n231));
  XOR2_X1   g0031(.A(G226), .B(G232), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT67), .B(G238), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n233), .B(new_n234), .Z(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G264), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n237), .B(G270), .Z(new_n238));
  XOR2_X1   g0038(.A(new_n235), .B(new_n238), .Z(G358));
  XNOR2_X1  g0039(.A(G87), .B(G97), .ZN(new_n240));
  INV_X1    g0040(.A(G107), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  INV_X1    g0042(.A(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G68), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  AND2_X1   g0048(.A1(KEYINPUT68), .A2(G223), .ZN(new_n249));
  NOR2_X1   g0049(.A1(KEYINPUT68), .A2(G223), .ZN(new_n250));
  OAI21_X1  g0050(.A(G1698), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT3), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G1698), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G222), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n251), .A2(new_n256), .A3(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G41), .ZN(new_n260));
  OAI211_X1 g0060(.A(G1), .B(G13), .C1(new_n253), .C2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  OAI211_X1 g0062(.A(new_n259), .B(new_n262), .C1(G77), .C2(new_n256), .ZN(new_n263));
  INV_X1    g0063(.A(G1), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n264), .B1(G41), .B2(G45), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n261), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G226), .ZN(new_n268));
  INV_X1    g0068(.A(G274), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n265), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n263), .A2(new_n268), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G200), .ZN(new_n273));
  INV_X1    g0073(.A(G190), .ZN(new_n274));
  INV_X1    g0074(.A(G20), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n275), .A2(G1), .ZN(new_n276));
  INV_X1    g0076(.A(G50), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  XOR2_X1   g0078(.A(new_n278), .B(KEYINPUT71), .Z(new_n279));
  NAND3_X1  g0079(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT69), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n280), .A2(new_n281), .A3(new_n207), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n281), .B1(new_n280), .B2(new_n207), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n276), .A2(G13), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n279), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  OAI21_X1  g0087(.A(G20), .B1(new_n204), .B2(G50), .ZN(new_n288));
  INV_X1    g0088(.A(G150), .ZN(new_n289));
  NOR2_X1   g0089(.A1(G20), .A2(G33), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n288), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT70), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(G58), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT8), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n294), .B(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n206), .A2(G33), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n292), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  OAI221_X1 g0100(.A(new_n287), .B1(G50), .B2(new_n286), .C1(new_n300), .C2(new_n285), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT9), .ZN(new_n302));
  OAI221_X1 g0102(.A(new_n273), .B1(new_n274), .B2(new_n272), .C1(new_n301), .C2(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n303), .B1(new_n302), .B2(new_n301), .ZN(new_n304));
  XOR2_X1   g0104(.A(new_n304), .B(KEYINPUT10), .Z(new_n305));
  NAND2_X1  g0105(.A1(new_n257), .A2(G223), .ZN(new_n306));
  NAND2_X1  g0106(.A1(G226), .A2(G1698), .ZN(new_n307));
  AOI22_X1  g0107(.A1(new_n254), .A2(new_n255), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n253), .A2(new_n219), .ZN(new_n309));
  OAI21_X1  g0109(.A(KEYINPUT80), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(G223), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n311), .A2(G1698), .ZN(new_n312));
  AND2_X1   g0112(.A1(G226), .A2(G1698), .ZN(new_n313));
  AND2_X1   g0113(.A1(KEYINPUT3), .A2(G33), .ZN(new_n314));
  NOR2_X1   g0114(.A1(KEYINPUT3), .A2(G33), .ZN(new_n315));
  OAI22_X1  g0115(.A1(new_n312), .A2(new_n313), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT80), .ZN(new_n317));
  INV_X1    g0117(.A(new_n309), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n316), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n310), .A2(new_n262), .A3(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(G179), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n271), .B1(new_n266), .B2(new_n218), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  AND3_X1   g0123(.A1(new_n320), .A2(new_n321), .A3(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(G169), .B1(new_n320), .B2(new_n323), .ZN(new_n325));
  OAI21_X1  g0125(.A(KEYINPUT81), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT81), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n320), .A2(new_n321), .A3(new_n323), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n307), .B1(new_n311), .B2(G1698), .ZN(new_n329));
  AOI211_X1 g0129(.A(KEYINPUT80), .B(new_n309), .C1(new_n256), .C2(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n317), .B1(new_n316), .B2(new_n318), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n322), .B1(new_n332), .B2(new_n262), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n327), .B(new_n328), .C1(new_n333), .C2(G169), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n326), .A2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT18), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n296), .A2(new_n286), .ZN(new_n338));
  NOR3_X1   g0138(.A1(new_n283), .A2(new_n284), .A3(new_n276), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n338), .B1(new_n339), .B2(new_n296), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(KEYINPUT79), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT79), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n338), .B(new_n342), .C1(new_n339), .C2(new_n296), .ZN(new_n343));
  AND2_X1   g0143(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT16), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n217), .A2(new_n211), .ZN(new_n346));
  OAI21_X1  g0146(.A(G20), .B1(new_n346), .B2(new_n203), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n290), .A2(G159), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AND2_X1   g0149(.A1(KEYINPUT64), .A2(G20), .ZN(new_n350));
  NOR2_X1   g0150(.A1(KEYINPUT64), .A2(G20), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n254), .B(new_n255), .C1(new_n350), .C2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT7), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(KEYINPUT78), .ZN(new_n355));
  NOR3_X1   g0155(.A1(new_n256), .A2(new_n353), .A3(G20), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT78), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n352), .A2(new_n358), .A3(new_n353), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n355), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  AOI211_X1 g0160(.A(new_n345), .B(new_n349), .C1(new_n360), .C2(G68), .ZN(new_n361));
  INV_X1    g0161(.A(new_n285), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n353), .B1(new_n256), .B2(G20), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n314), .A2(new_n315), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n364), .A2(new_n206), .A3(KEYINPUT7), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n349), .B1(new_n366), .B2(G68), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n362), .B1(new_n367), .B2(KEYINPUT16), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n344), .B1(new_n361), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n336), .A2(new_n337), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n341), .A2(new_n343), .ZN(new_n371));
  INV_X1    g0171(.A(new_n349), .ZN(new_n372));
  AND3_X1   g0172(.A1(new_n352), .A2(new_n358), .A3(new_n353), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n358), .B1(new_n352), .B2(new_n353), .ZN(new_n374));
  NOR3_X1   g0174(.A1(new_n373), .A2(new_n374), .A3(new_n356), .ZN(new_n375));
  OAI211_X1 g0175(.A(KEYINPUT16), .B(new_n372), .C1(new_n375), .C2(new_n211), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n352), .A2(new_n353), .ZN(new_n377));
  AOI21_X1  g0177(.A(KEYINPUT7), .B1(new_n364), .B2(new_n275), .ZN(new_n378));
  OAI21_X1  g0178(.A(G68), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(new_n372), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n285), .B1(new_n380), .B2(new_n345), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n371), .B1(new_n376), .B2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(G200), .ZN(new_n383));
  OR2_X1    g0183(.A1(new_n333), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n333), .A2(G190), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n382), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT17), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n382), .A2(KEYINPUT17), .A3(new_n384), .A4(new_n385), .ZN(new_n389));
  OAI21_X1  g0189(.A(KEYINPUT18), .B1(new_n335), .B2(new_n382), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n370), .A2(new_n388), .A3(new_n389), .A4(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(G169), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n272), .A2(new_n393), .ZN(new_n394));
  OR2_X1    g0194(.A1(new_n272), .A2(G179), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n301), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n286), .A2(G77), .ZN(new_n397));
  XOR2_X1   g0197(.A(KEYINPUT15), .B(G87), .Z(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(KEYINPUT73), .ZN(new_n399));
  XNOR2_X1  g0199(.A(KEYINPUT15), .B(G87), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT73), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n399), .A2(new_n402), .ZN(new_n403));
  OR3_X1    g0203(.A1(new_n403), .A2(KEYINPUT74), .A3(new_n298), .ZN(new_n404));
  XOR2_X1   g0204(.A(KEYINPUT8), .B(G58), .Z(new_n405));
  NOR2_X1   g0205(.A1(new_n350), .A2(new_n351), .ZN(new_n406));
  AOI22_X1  g0206(.A1(new_n405), .A2(new_n290), .B1(new_n406), .B2(G77), .ZN(new_n407));
  OAI21_X1  g0207(.A(KEYINPUT74), .B1(new_n403), .B2(new_n298), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n404), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n397), .B1(new_n409), .B2(new_n362), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n339), .A2(G77), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT72), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n413), .B1(new_n364), .B2(new_n218), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n256), .A2(KEYINPUT72), .A3(G232), .A4(new_n257), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n413), .B1(new_n256), .B2(G238), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n414), .B(new_n415), .C1(new_n416), .C2(new_n257), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n256), .A2(new_n241), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n262), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n267), .A2(G244), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n419), .A2(new_n271), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(new_n393), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n419), .A2(new_n321), .A3(new_n271), .A4(new_n420), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n412), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n305), .A2(new_n392), .A3(new_n396), .A4(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n256), .A2(G232), .A3(G1698), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(KEYINPUT75), .ZN(new_n427));
  NAND2_X1  g0227(.A1(G33), .A2(G97), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n256), .A2(G226), .A3(new_n257), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT75), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n256), .A2(new_n430), .A3(G232), .A4(G1698), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n427), .A2(new_n428), .A3(new_n429), .A4(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(new_n262), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n271), .B1(new_n266), .B2(new_n212), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(KEYINPUT13), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n434), .B1(new_n432), .B2(new_n262), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT13), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n437), .A2(KEYINPUT76), .A3(new_n440), .ZN(new_n441));
  OR3_X1    g0241(.A1(new_n438), .A2(KEYINPUT76), .A3(new_n439), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n441), .A2(G169), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(KEYINPUT14), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT14), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n441), .A2(new_n445), .A3(G169), .A4(new_n442), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT77), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n437), .A2(new_n440), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n447), .B1(new_n448), .B2(new_n321), .ZN(new_n449));
  INV_X1    g0249(.A(new_n448), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n450), .A2(KEYINPUT77), .A3(G179), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n444), .A2(new_n446), .A3(new_n449), .A4(new_n451), .ZN(new_n452));
  AOI22_X1  g0252(.A1(new_n299), .A2(G77), .B1(G50), .B2(new_n290), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n453), .B1(new_n275), .B2(G68), .ZN(new_n454));
  AND3_X1   g0254(.A1(new_n454), .A2(KEYINPUT11), .A3(new_n362), .ZN(new_n455));
  AOI21_X1  g0255(.A(KEYINPUT11), .B1(new_n454), .B2(new_n362), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n286), .A2(G68), .ZN(new_n457));
  XNOR2_X1  g0257(.A(new_n457), .B(KEYINPUT12), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n339), .A2(G68), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  OR4_X1    g0260(.A1(new_n455), .A2(new_n456), .A3(new_n458), .A4(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n452), .A2(new_n461), .ZN(new_n462));
  AND2_X1   g0262(.A1(new_n441), .A2(new_n442), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n461), .B1(new_n463), .B2(G200), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n450), .A2(G190), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AND2_X1   g0266(.A1(new_n421), .A2(G200), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n410), .B(new_n411), .C1(new_n274), .C2(new_n421), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n462), .B(new_n466), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n425), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n256), .A2(KEYINPUT4), .A3(G244), .A4(new_n257), .ZN(new_n471));
  OAI21_X1  g0271(.A(G244), .B1(new_n314), .B2(new_n315), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT4), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(G33), .A2(G283), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n471), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n256), .A2(G250), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n257), .B1(new_n477), .B2(KEYINPUT4), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n262), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(G45), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n480), .A2(G1), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n481), .B1(KEYINPUT5), .B2(new_n260), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n269), .B1(new_n482), .B2(KEYINPUT82), .ZN(new_n483));
  AND2_X1   g0283(.A1(new_n260), .A2(KEYINPUT5), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n262), .A2(new_n484), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n483), .B(new_n485), .C1(KEYINPUT82), .C2(new_n482), .ZN(new_n486));
  OAI211_X1 g0286(.A(G257), .B(new_n261), .C1(new_n482), .C2(new_n484), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n479), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n393), .ZN(new_n489));
  INV_X1    g0289(.A(new_n286), .ZN(new_n490));
  INV_X1    g0290(.A(G97), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n264), .A2(G33), .ZN(new_n493));
  AND3_X1   g0293(.A1(new_n285), .A2(new_n286), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(G97), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n241), .B1(new_n363), .B2(new_n365), .ZN(new_n496));
  INV_X1    g0296(.A(G77), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n291), .A2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT6), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n491), .A2(new_n241), .ZN(new_n500));
  NOR2_X1   g0300(.A1(G97), .A2(G107), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n241), .A2(KEYINPUT6), .A3(G97), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n206), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NOR3_X1   g0304(.A1(new_n496), .A2(new_n498), .A3(new_n504), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n492), .B(new_n495), .C1(new_n505), .C2(new_n285), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n479), .A2(new_n321), .A3(new_n486), .A4(new_n487), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n489), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(KEYINPUT83), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT83), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n489), .A2(new_n506), .A3(new_n510), .A4(new_n507), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  OR2_X1    g0312(.A1(KEYINPUT64), .A2(G20), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT23), .ZN(new_n514));
  NAND2_X1  g0314(.A1(KEYINPUT64), .A2(G20), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n513), .A2(new_n514), .A3(new_n241), .A4(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT89), .ZN(new_n517));
  XNOR2_X1  g0317(.A(new_n516), .B(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT88), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT22), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n256), .A2(new_n206), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n519), .B(new_n520), .C1(new_n521), .C2(new_n219), .ZN(new_n522));
  NAND2_X1  g0322(.A1(KEYINPUT23), .A2(G107), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n514), .B1(new_n253), .B2(new_n243), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n275), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n518), .A2(new_n522), .A3(new_n523), .A4(new_n525), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n519), .B1(new_n521), .B2(new_n219), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n256), .A2(new_n206), .A3(KEYINPUT88), .A4(G87), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n527), .A2(KEYINPUT22), .A3(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  OAI21_X1  g0330(.A(KEYINPUT24), .B1(new_n526), .B2(new_n530), .ZN(new_n531));
  AND3_X1   g0331(.A1(new_n522), .A2(new_n523), .A3(new_n525), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT24), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n532), .A2(new_n533), .A3(new_n529), .A4(new_n518), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n362), .ZN(new_n536));
  AND2_X1   g0336(.A1(new_n494), .A2(G107), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n490), .A2(new_n241), .ZN(new_n538));
  XNOR2_X1  g0338(.A(new_n538), .B(KEYINPUT25), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  OAI211_X1 g0340(.A(G257), .B(G1698), .C1(new_n314), .C2(new_n315), .ZN(new_n541));
  OAI211_X1 g0341(.A(G250), .B(new_n257), .C1(new_n314), .C2(new_n315), .ZN(new_n542));
  NAND2_X1  g0342(.A1(G33), .A2(G294), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n262), .ZN(new_n545));
  OAI211_X1 g0345(.A(G264), .B(new_n261), .C1(new_n482), .C2(new_n484), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n486), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(G200), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n548), .A2(G190), .A3(new_n486), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n536), .A2(new_n540), .A3(new_n550), .A4(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(new_n488), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n553), .A2(new_n383), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n488), .A2(new_n274), .ZN(new_n555));
  OR3_X1    g0355(.A1(new_n554), .A2(new_n506), .A3(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT19), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n557), .B1(new_n298), .B2(new_n491), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n256), .A2(new_n206), .A3(G68), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n428), .A2(new_n557), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n406), .A2(new_n560), .ZN(new_n561));
  NOR3_X1   g0361(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n562));
  XNOR2_X1  g0362(.A(new_n562), .B(KEYINPUT85), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n558), .B(new_n559), .C1(new_n561), .C2(new_n563), .ZN(new_n564));
  AOI22_X1  g0364(.A1(new_n564), .A2(new_n362), .B1(new_n490), .B2(new_n403), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n494), .A2(new_n402), .A3(new_n399), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n481), .A2(new_n269), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n220), .B1(new_n480), .B2(G1), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n568), .A2(new_n261), .A3(new_n569), .ZN(new_n570));
  OAI22_X1  g0370(.A1(new_n472), .A2(new_n257), .B1(new_n253), .B2(new_n243), .ZN(new_n571));
  OAI211_X1 g0371(.A(G238), .B(new_n257), .C1(new_n314), .C2(new_n315), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT84), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n256), .A2(KEYINPUT84), .A3(G238), .A4(new_n257), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n571), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n321), .B(new_n570), .C1(new_n576), .C2(new_n261), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n570), .B1(new_n576), .B2(new_n261), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n393), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n567), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n578), .A2(G200), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n494), .A2(G87), .ZN(new_n582));
  OAI211_X1 g0382(.A(G190), .B(new_n570), .C1(new_n576), .C2(new_n261), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n581), .A2(new_n565), .A3(new_n582), .A4(new_n583), .ZN(new_n584));
  AND2_X1   g0384(.A1(new_n580), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n512), .A2(new_n552), .A3(new_n556), .A4(new_n585), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n549), .A2(G179), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n587), .B1(new_n393), .B2(new_n549), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n285), .B1(new_n531), .B2(new_n534), .ZN(new_n589));
  INV_X1    g0389(.A(new_n540), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  OAI221_X1 g0391(.A(new_n475), .B1(G33), .B2(new_n491), .C1(new_n350), .C2(new_n351), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n280), .A2(new_n207), .B1(G20), .B2(new_n243), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT20), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n592), .A2(KEYINPUT20), .A3(new_n593), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n596), .A2(new_n597), .B1(new_n243), .B2(new_n490), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n494), .A2(G116), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n393), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  OAI211_X1 g0400(.A(G270), .B(new_n261), .C1(new_n482), .C2(new_n484), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  OAI211_X1 g0402(.A(G257), .B(new_n257), .C1(new_n314), .C2(new_n315), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT86), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n256), .A2(KEYINPUT86), .A3(G257), .A4(new_n257), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n256), .A2(G264), .A3(G1698), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n364), .A2(G303), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n605), .A2(new_n606), .A3(new_n607), .A4(new_n608), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n602), .B1(new_n609), .B2(new_n262), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n486), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT21), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(KEYINPUT87), .ZN(new_n613));
  AND3_X1   g0413(.A1(new_n600), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n613), .B1(new_n600), .B2(new_n611), .ZN(new_n615));
  AND2_X1   g0415(.A1(new_n598), .A2(new_n599), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n610), .A2(G179), .A3(new_n486), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NOR3_X1   g0418(.A1(new_n614), .A2(new_n615), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n611), .A2(G200), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n620), .B(new_n616), .C1(new_n274), .C2(new_n611), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n591), .A2(new_n619), .A3(new_n621), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n586), .A2(new_n622), .ZN(new_n623));
  AND2_X1   g0423(.A1(new_n470), .A2(new_n623), .ZN(G372));
  INV_X1    g0424(.A(new_n396), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n462), .A2(new_n424), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n388), .A2(new_n389), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n626), .A2(new_n627), .A3(new_n466), .ZN(new_n628));
  OAI21_X1  g0428(.A(KEYINPUT90), .B1(new_n335), .B2(new_n382), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT90), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n369), .A2(new_n630), .A3(new_n326), .A4(new_n334), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n632), .A2(new_n337), .ZN(new_n633));
  AOI21_X1  g0433(.A(KEYINPUT18), .B1(new_n629), .B2(new_n631), .ZN(new_n634));
  OR2_X1    g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n628), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n625), .B1(new_n636), .B2(new_n305), .ZN(new_n637));
  INV_X1    g0437(.A(new_n470), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n585), .A2(new_n509), .A3(new_n511), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(KEYINPUT26), .ZN(new_n640));
  INV_X1    g0440(.A(new_n508), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n585), .A2(new_n641), .ZN(new_n642));
  OAI211_X1 g0442(.A(new_n640), .B(new_n580), .C1(KEYINPUT26), .C2(new_n642), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n586), .B1(new_n619), .B2(new_n591), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n637), .B1(new_n638), .B2(new_n645), .ZN(G369));
  AND4_X1   g0446(.A1(new_n536), .A2(new_n540), .A3(new_n550), .A4(new_n551), .ZN(new_n647));
  INV_X1    g0447(.A(G13), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n406), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  OR3_X1    g0450(.A1(new_n650), .A2(KEYINPUT27), .A3(G1), .ZN(new_n651));
  OAI21_X1  g0451(.A(KEYINPUT27), .B1(new_n650), .B2(G1), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n651), .A2(new_n652), .A3(G213), .ZN(new_n653));
  INV_X1    g0453(.A(G343), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n656), .B1(new_n536), .B2(new_n540), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n591), .B1(new_n647), .B2(new_n657), .ZN(new_n658));
  OAI211_X1 g0458(.A(new_n588), .B(new_n656), .C1(new_n589), .C2(new_n590), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT91), .ZN(new_n661));
  OR2_X1    g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n660), .A2(new_n661), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n619), .ZN(new_n665));
  OR2_X1    g0465(.A1(new_n656), .A2(new_n616), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n665), .A2(new_n666), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n667), .A2(new_n621), .A3(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(G330), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n619), .A2(new_n655), .ZN(new_n672));
  OR2_X1    g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n664), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(new_n659), .ZN(G399));
  INV_X1    g0475(.A(new_n225), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n676), .A2(G41), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(G1), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n563), .A2(new_n243), .ZN(new_n680));
  OAI22_X1  g0480(.A1(new_n679), .A2(new_n680), .B1(new_n205), .B2(new_n678), .ZN(new_n681));
  XNOR2_X1  g0481(.A(new_n681), .B(KEYINPUT28), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT93), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n683), .B1(new_n623), .B2(new_n656), .ZN(new_n684));
  NOR4_X1   g0484(.A1(new_n586), .A2(new_n622), .A3(KEYINPUT93), .A4(new_n655), .ZN(new_n685));
  OR2_X1    g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n609), .A2(new_n262), .ZN(new_n687));
  AND4_X1   g0487(.A1(G179), .A2(new_n687), .A3(new_n486), .A4(new_n601), .ZN(new_n688));
  INV_X1    g0488(.A(new_n571), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n574), .A2(new_n575), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n261), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n570), .ZN(new_n692));
  NOR3_X1   g0492(.A1(new_n691), .A2(new_n547), .A3(new_n692), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n688), .A2(new_n553), .A3(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT30), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n688), .A2(new_n553), .A3(KEYINPUT30), .A4(new_n693), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n486), .B1(new_n548), .B2(new_n610), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n698), .A2(new_n321), .A3(new_n578), .A4(new_n488), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n696), .A2(new_n697), .A3(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(KEYINPUT31), .B1(new_n700), .B2(new_n655), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n701), .A2(KEYINPUT92), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n700), .A2(KEYINPUT31), .A3(new_n655), .ZN(new_n703));
  MUX2_X1   g0503(.A(KEYINPUT92), .B(new_n702), .S(new_n703), .Z(new_n704));
  AOI21_X1  g0504(.A(new_n670), .B1(new_n686), .B2(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n645), .A2(new_n655), .ZN(new_n706));
  OR2_X1    g0506(.A1(new_n706), .A2(KEYINPUT29), .ZN(new_n707));
  OR2_X1    g0507(.A1(new_n639), .A2(KEYINPUT26), .ZN(new_n708));
  INV_X1    g0508(.A(new_n580), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n709), .B1(new_n642), .B2(KEYINPUT26), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n591), .A2(new_n619), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n711), .B(KEYINPUT94), .ZN(new_n712));
  OAI211_X1 g0512(.A(new_n708), .B(new_n710), .C1(new_n712), .C2(new_n586), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n713), .A2(KEYINPUT29), .A3(new_n656), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n705), .B1(new_n707), .B2(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n682), .B1(new_n715), .B2(G1), .ZN(G364));
  INV_X1    g0516(.A(new_n671), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT95), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n718), .B1(new_n650), .B2(new_n480), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n649), .A2(KEYINPUT95), .A3(G45), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n719), .A2(G1), .A3(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(new_n677), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n669), .A2(new_n670), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n717), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n207), .B1(G20), .B2(new_n393), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n406), .A2(G179), .A3(G190), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(G200), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(G322), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n727), .A2(new_n383), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n256), .B1(new_n732), .B2(G326), .ZN(new_n733));
  INV_X1    g0533(.A(G303), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n383), .A2(G179), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n735), .A2(G20), .A3(G190), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n206), .A2(G190), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(G179), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(G200), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(G311), .ZN(new_n741));
  OAI221_X1 g0541(.A(new_n733), .B1(new_n734), .B2(new_n736), .C1(new_n740), .C2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n737), .A2(new_n735), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  AOI211_X1 g0544(.A(new_n731), .B(new_n742), .C1(G283), .C2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(G179), .A2(G200), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n737), .A2(new_n746), .ZN(new_n747));
  XOR2_X1   g0547(.A(new_n747), .B(KEYINPUT97), .Z(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(G329), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n746), .A2(G190), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n406), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(G294), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n738), .A2(new_n383), .ZN(new_n754));
  XNOR2_X1  g0554(.A(KEYINPUT33), .B(G317), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n745), .A2(new_n750), .A3(new_n753), .A4(new_n756), .ZN(new_n757));
  XNOR2_X1  g0557(.A(new_n757), .B(KEYINPUT98), .ZN(new_n758));
  AOI22_X1  g0558(.A1(new_n754), .A2(G68), .B1(G50), .B2(new_n732), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n759), .B1(new_n241), .B2(new_n743), .ZN(new_n760));
  INV_X1    g0560(.A(new_n747), .ZN(new_n761));
  XOR2_X1   g0561(.A(KEYINPUT96), .B(G159), .Z(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g0563(.A(new_n763), .B(KEYINPUT32), .ZN(new_n764));
  INV_X1    g0564(.A(new_n736), .ZN(new_n765));
  AOI211_X1 g0565(.A(new_n760), .B(new_n764), .C1(G87), .C2(new_n765), .ZN(new_n766));
  AOI22_X1  g0566(.A1(new_n728), .A2(G58), .B1(G97), .B2(new_n752), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n766), .A2(new_n256), .A3(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n768), .B1(G77), .B2(new_n739), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n726), .B1(new_n758), .B2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(G13), .A2(G33), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(G20), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n669), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n247), .A2(G45), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n676), .A2(new_n256), .ZN(new_n776));
  OAI211_X1 g0576(.A(new_n775), .B(new_n776), .C1(G45), .C2(new_n205), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n676), .A2(new_n364), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(G355), .ZN(new_n779));
  OAI211_X1 g0579(.A(new_n777), .B(new_n779), .C1(G116), .C2(new_n225), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n773), .A2(new_n726), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND4_X1  g0582(.A1(new_n770), .A2(new_n722), .A3(new_n774), .A4(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n725), .A2(new_n783), .ZN(G396));
  NOR2_X1   g0584(.A1(new_n468), .A2(new_n467), .ZN(new_n785));
  INV_X1    g0585(.A(KEYINPUT100), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n424), .A2(new_n786), .ZN(new_n787));
  NAND4_X1  g0587(.A1(new_n412), .A2(KEYINPUT100), .A3(new_n422), .A4(new_n423), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n785), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n412), .A2(new_n655), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n422), .A2(new_n423), .ZN(new_n791));
  OR3_X1    g0591(.A1(new_n790), .A2(KEYINPUT101), .A3(new_n791), .ZN(new_n792));
  OAI21_X1  g0592(.A(KEYINPUT101), .B1(new_n790), .B2(new_n791), .ZN(new_n793));
  AOI22_X1  g0593(.A1(new_n789), .A2(new_n790), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(KEYINPUT102), .B1(new_n706), .B2(new_n795), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n796), .B1(new_n706), .B2(new_n795), .ZN(new_n797));
  OAI211_X1 g0597(.A(KEYINPUT102), .B(new_n794), .C1(new_n645), .C2(new_n655), .ZN(new_n798));
  INV_X1    g0598(.A(new_n705), .ZN(new_n799));
  INV_X1    g0599(.A(KEYINPUT103), .ZN(new_n800));
  OAI211_X1 g0600(.A(new_n797), .B(new_n798), .C1(new_n799), .C2(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n799), .A2(new_n800), .ZN(new_n802));
  OR2_X1    g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n801), .A2(new_n802), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n803), .A2(new_n723), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n794), .A2(new_n771), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n726), .A2(new_n771), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(new_n497), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n754), .A2(G150), .B1(G143), .B2(new_n728), .ZN(new_n809));
  INV_X1    g0609(.A(G137), .ZN(new_n810));
  INV_X1    g0610(.A(new_n732), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n809), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n812), .B1(new_n739), .B2(new_n762), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n813), .B(KEYINPUT34), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n364), .B1(new_n749), .B2(G132), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n752), .A2(G58), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n744), .A2(G68), .B1(G50), .B2(new_n765), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n815), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n728), .A2(G294), .B1(G97), .B2(new_n752), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(KEYINPUT99), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n820), .B1(G303), .B2(new_n732), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n744), .A2(G87), .ZN(new_n822));
  AOI22_X1  g0622(.A1(new_n754), .A2(G283), .B1(G107), .B2(new_n765), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n739), .A2(G116), .ZN(new_n824));
  NAND4_X1  g0624(.A1(new_n821), .A2(new_n822), .A3(new_n823), .A4(new_n824), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n364), .B1(new_n748), .B2(new_n741), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n814), .A2(new_n818), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(new_n726), .ZN(new_n828));
  NAND4_X1  g0628(.A1(new_n806), .A2(new_n722), .A3(new_n808), .A4(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n805), .A2(new_n829), .ZN(G384));
  INV_X1    g0630(.A(KEYINPUT106), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n382), .A2(new_n653), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n376), .A2(new_n381), .ZN(new_n834));
  AND4_X1   g0634(.A1(new_n384), .A2(new_n834), .A3(new_n385), .A4(new_n344), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n835), .B1(new_n629), .B2(new_n631), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT105), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n833), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  AOI211_X1 g0638(.A(KEYINPUT105), .B(new_n835), .C1(new_n629), .C2(new_n631), .ZN(new_n839));
  OAI21_X1  g0639(.A(KEYINPUT37), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n835), .A2(KEYINPUT37), .ZN(new_n841));
  INV_X1    g0641(.A(new_n653), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n369), .B1(new_n336), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n627), .B1(new_n633), .B2(new_n634), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n840), .A2(new_n844), .B1(new_n832), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n831), .B1(new_n846), .B2(KEYINPUT38), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT38), .ZN(new_n848));
  INV_X1    g0648(.A(new_n844), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n632), .A2(new_n386), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(KEYINPUT105), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n836), .A2(new_n837), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n851), .A2(new_n833), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n849), .B1(new_n853), .B2(KEYINPUT37), .ZN(new_n854));
  AND2_X1   g0654(.A1(new_n845), .A2(new_n832), .ZN(new_n855));
  OAI211_X1 g0655(.A(KEYINPUT106), .B(new_n848), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n376), .A2(new_n362), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n349), .B1(new_n360), .B2(G68), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n858), .A2(KEYINPUT16), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n344), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(new_n842), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n391), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n336), .A2(new_n860), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n864), .A2(new_n861), .A3(new_n386), .ZN(new_n865));
  AND2_X1   g0665(.A1(new_n865), .A2(KEYINPUT37), .ZN(new_n866));
  OAI211_X1 g0666(.A(KEYINPUT38), .B(new_n863), .C1(new_n866), .C2(new_n849), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n847), .A2(new_n856), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(KEYINPUT110), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT108), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n701), .B1(new_n870), .B2(new_n703), .ZN(new_n871));
  AOI211_X1 g0671(.A(KEYINPUT108), .B(KEYINPUT31), .C1(new_n700), .C2(new_n655), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n873), .B1(new_n684), .B2(new_n685), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n461), .A2(new_n655), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n462), .A2(new_n466), .A3(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n452), .A2(new_n461), .A3(new_n655), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n794), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AND3_X1   g0678(.A1(new_n874), .A2(KEYINPUT40), .A3(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT110), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n847), .A2(new_n856), .A3(new_n880), .A4(new_n867), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n869), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  AND2_X1   g0682(.A1(new_n391), .A2(new_n862), .ZN(new_n883));
  AOI22_X1  g0683(.A1(new_n865), .A2(KEYINPUT37), .B1(new_n841), .B2(new_n843), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n848), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n867), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n874), .A2(new_n886), .A3(new_n878), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT40), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(KEYINPUT109), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT109), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n887), .A2(new_n891), .A3(new_n888), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n882), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n470), .A2(new_n874), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n894), .B(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(G330), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n707), .A2(new_n470), .A3(new_n714), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n637), .ZN(new_n901));
  XOR2_X1   g0701(.A(new_n901), .B(KEYINPUT107), .Z(new_n902));
  NAND2_X1  g0702(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  OR2_X1    g0704(.A1(new_n635), .A2(new_n842), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n706), .A2(new_n795), .ZN(new_n906));
  AND3_X1   g0706(.A1(new_n787), .A2(new_n656), .A3(new_n788), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n876), .A2(new_n877), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n886), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n905), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT39), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n868), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n912), .A2(KEYINPUT39), .ZN(new_n916));
  AND2_X1   g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n462), .A2(new_n655), .ZN(new_n918));
  XOR2_X1   g0718(.A(new_n918), .B(KEYINPUT104), .Z(new_n919));
  AOI21_X1  g0719(.A(new_n913), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n899), .A2(new_n902), .ZN(new_n922));
  OR3_X1    g0722(.A1(new_n904), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n921), .B1(new_n904), .B2(new_n922), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n923), .B(new_n924), .C1(new_n264), .C2(new_n649), .ZN(new_n925));
  AND2_X1   g0725(.A1(new_n502), .A2(new_n503), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT35), .ZN(new_n927));
  AOI211_X1 g0727(.A(new_n207), .B(new_n206), .C1(new_n926), .C2(new_n927), .ZN(new_n928));
  OAI211_X1 g0728(.A(new_n928), .B(G116), .C1(new_n927), .C2(new_n926), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n929), .B(KEYINPUT36), .ZN(new_n930));
  OAI21_X1  g0730(.A(G77), .B1(new_n217), .B2(new_n211), .ZN(new_n931));
  OAI22_X1  g0731(.A1(new_n205), .A2(new_n931), .B1(G50), .B2(new_n211), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n932), .A2(G1), .A3(new_n648), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n925), .A2(new_n930), .A3(new_n933), .ZN(G367));
  NAND2_X1  g0734(.A1(new_n664), .A2(new_n672), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n655), .A2(new_n506), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n512), .A2(new_n556), .A3(new_n936), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n937), .B(KEYINPUT111), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT42), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n941), .B(KEYINPUT112), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n939), .A2(new_n940), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n641), .A2(new_n655), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n938), .A2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n512), .B1(new_n946), .B2(new_n591), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n943), .B1(new_n656), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n942), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n565), .A2(new_n582), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(new_n655), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n585), .A2(new_n951), .ZN(new_n952));
  OR2_X1    g0752(.A1(new_n580), .A2(new_n951), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT43), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n954), .A2(KEYINPUT43), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n949), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  NAND4_X1  g0759(.A1(new_n942), .A2(new_n956), .A3(new_n955), .A4(new_n948), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n662), .A2(new_n663), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n962), .A2(new_n717), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n964), .A2(new_n946), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n961), .B(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(new_n721), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n935), .A2(new_n659), .A3(new_n945), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n968), .A2(KEYINPUT113), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(KEYINPUT113), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT45), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n945), .B1(new_n935), .B2(new_n659), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT44), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n969), .A2(KEYINPUT45), .A3(new_n970), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n973), .A2(new_n975), .A3(new_n964), .A4(new_n976), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n673), .B(new_n962), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n715), .A2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n977), .A2(new_n980), .ZN(new_n981));
  AND2_X1   g0781(.A1(new_n981), .A2(new_n715), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n677), .B(KEYINPUT41), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n967), .B1(new_n982), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n966), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n364), .B1(new_n739), .B2(G50), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n744), .A2(G77), .ZN(new_n988));
  OAI211_X1 g0788(.A(new_n987), .B(new_n988), .C1(new_n217), .C2(new_n736), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n754), .A2(new_n762), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n732), .A2(G143), .ZN(new_n991));
  OAI211_X1 g0791(.A(new_n990), .B(new_n991), .C1(new_n729), .C2(new_n289), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n747), .A2(new_n810), .ZN(new_n993));
  INV_X1    g0793(.A(new_n752), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n994), .A2(new_n211), .ZN(new_n995));
  NOR4_X1   g0795(.A1(new_n989), .A2(new_n992), .A3(new_n993), .A4(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n765), .A2(G116), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT46), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n744), .A2(G97), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n998), .A2(new_n364), .A3(new_n999), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(G283), .A2(new_n739), .B1(new_n754), .B2(G294), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n761), .A2(G317), .ZN(new_n1002));
  OAI211_X1 g0802(.A(new_n1001), .B(new_n1002), .C1(new_n241), .C2(new_n994), .ZN(new_n1003));
  AOI211_X1 g0803(.A(new_n1000), .B(new_n1003), .C1(G311), .C2(new_n732), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n728), .A2(G303), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n996), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n1006), .B(KEYINPUT47), .Z(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(new_n726), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n776), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n781), .B1(new_n225), .B2(new_n403), .C1(new_n238), .C2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1008), .A2(new_n722), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n773), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n954), .A2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n986), .A2(new_n1015), .ZN(G387));
  NAND2_X1  g0816(.A1(new_n978), .A2(new_n721), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n403), .A2(new_n994), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n754), .A2(new_n297), .B1(G159), .B2(new_n732), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n1019), .B1(new_n211), .B2(new_n740), .C1(new_n497), .C2(new_n736), .ZN(new_n1020));
  AOI211_X1 g0820(.A(new_n1018), .B(new_n1020), .C1(G150), .C2(new_n761), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n728), .A2(G50), .ZN(new_n1022));
  NAND4_X1  g0822(.A1(new_n1021), .A2(new_n256), .A3(new_n999), .A4(new_n1022), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n754), .A2(G311), .B1(G317), .B2(new_n728), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n1024), .B1(new_n734), .B2(new_n740), .C1(new_n730), .C2(new_n811), .ZN(new_n1025));
  XOR2_X1   g0825(.A(KEYINPUT114), .B(KEYINPUT48), .Z(new_n1026));
  XNOR2_X1  g0826(.A(new_n1025), .B(new_n1026), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(G294), .A2(new_n765), .B1(new_n752), .B2(G283), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1027), .A2(KEYINPUT49), .A3(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n744), .A2(G116), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n761), .A2(G326), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1029), .A2(new_n364), .A3(new_n1030), .A4(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(KEYINPUT49), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1023), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1009), .B1(new_n235), .B2(G45), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1035), .B1(new_n680), .B2(new_n778), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n405), .A2(new_n277), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT50), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n211), .A2(new_n497), .ZN(new_n1039));
  NOR4_X1   g0839(.A1(new_n1038), .A2(G45), .A3(new_n1039), .A4(new_n680), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n1036), .A2(new_n1040), .B1(G107), .B2(new_n225), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n1034), .A2(new_n726), .B1(new_n781), .B2(new_n1041), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n722), .B(new_n1042), .C1(new_n664), .C2(new_n1012), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n715), .A2(new_n978), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1044), .A2(KEYINPUT115), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(new_n677), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n979), .B1(new_n1044), .B2(KEYINPUT115), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n1017), .B(new_n1043), .C1(new_n1046), .C2(new_n1047), .ZN(G393));
  NAND3_X1  g0848(.A1(new_n973), .A2(new_n975), .A3(new_n976), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n963), .ZN(new_n1050));
  AND2_X1   g0850(.A1(new_n1050), .A2(new_n977), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(new_n721), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n946), .A2(new_n773), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(G150), .A2(new_n732), .B1(new_n728), .B2(G159), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT116), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n1055), .B(KEYINPUT51), .Z(new_n1056));
  NOR2_X1   g0856(.A1(new_n994), .A2(new_n497), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n364), .B(new_n1057), .C1(G143), .C2(new_n761), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n754), .A2(G50), .B1(G68), .B2(new_n765), .ZN(new_n1059));
  NAND4_X1  g0859(.A1(new_n1056), .A2(new_n822), .A3(new_n1058), .A4(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(new_n405), .B2(new_n739), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(G311), .A2(new_n728), .B1(new_n732), .B2(G317), .ZN(new_n1062));
  XOR2_X1   g0862(.A(new_n1062), .B(KEYINPUT52), .Z(new_n1063));
  NAND2_X1  g0863(.A1(new_n765), .A2(G283), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n739), .A2(G294), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1063), .A2(new_n364), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n994), .A2(new_n243), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n747), .A2(new_n730), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n754), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n1069), .A2(new_n734), .B1(new_n743), .B2(new_n241), .ZN(new_n1070));
  NOR4_X1   g0870(.A1(new_n1066), .A2(new_n1067), .A3(new_n1068), .A4(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n726), .B1(new_n1061), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n244), .A2(new_n776), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n1073), .B(new_n781), .C1(new_n491), .C2(new_n225), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n1053), .A2(new_n722), .A3(new_n1072), .A4(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1050), .A2(new_n977), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(new_n979), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n981), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n1052), .B(new_n1075), .C1(new_n1078), .C2(new_n678), .ZN(G390));
  OAI211_X1 g0879(.A(new_n900), .B(new_n637), .C1(new_n670), .C2(new_n895), .ZN(new_n1080));
  AND3_X1   g0880(.A1(new_n705), .A2(new_n795), .A3(new_n910), .ZN(new_n1081));
  AND2_X1   g0881(.A1(new_n874), .A2(G330), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n910), .B1(new_n1082), .B2(new_n795), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n713), .A2(new_n656), .A3(new_n795), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1084), .A2(new_n908), .ZN(new_n1085));
  OR3_X1    g0885(.A1(new_n1081), .A2(new_n1083), .A3(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n910), .B1(new_n705), .B2(new_n795), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n874), .A2(new_n878), .A3(G330), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n909), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1080), .B1(new_n1086), .B2(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n919), .B1(new_n1085), .B2(new_n910), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n869), .A2(new_n1093), .A3(new_n881), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n919), .B1(new_n909), .B2(new_n910), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(new_n915), .B2(new_n916), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1088), .B1(new_n1095), .B2(new_n1097), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n1094), .B(new_n1081), .C1(new_n917), .C2(new_n1096), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1092), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n1091), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1100), .A2(new_n1102), .A3(new_n677), .ZN(new_n1103));
  OAI221_X1 g0903(.A(new_n364), .B1(new_n497), .B2(new_n994), .C1(new_n729), .C2(new_n243), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n749), .A2(G294), .B1(G87), .B2(new_n765), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n754), .A2(G107), .B1(new_n744), .B2(G68), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1105), .B(new_n1106), .C1(new_n491), .C2(new_n740), .ZN(new_n1107));
  AOI211_X1 g0907(.A(new_n1104), .B(new_n1107), .C1(G283), .C2(new_n732), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n765), .A2(G150), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(new_n1109), .B(KEYINPUT53), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n749), .A2(G125), .ZN(new_n1111));
  INV_X1    g0911(.A(G159), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n743), .A2(new_n277), .B1(new_n994), .B2(new_n1112), .ZN(new_n1113));
  XOR2_X1   g0913(.A(KEYINPUT54), .B(G143), .Z(new_n1114));
  AOI21_X1  g0914(.A(new_n1113), .B1(new_n739), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n754), .A2(G137), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n364), .B1(new_n732), .B2(G128), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n1111), .A2(new_n1115), .A3(new_n1116), .A4(new_n1117), .ZN(new_n1118));
  AOI211_X1 g0918(.A(new_n1110), .B(new_n1118), .C1(G132), .C2(new_n728), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n726), .B1(new_n1108), .B2(new_n1119), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n722), .B(new_n1120), .C1(new_n917), .C2(new_n772), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1121), .B1(new_n296), .B2(new_n807), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1122), .B1(new_n721), .B2(new_n1101), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1103), .A2(new_n1123), .ZN(G378));
  NAND2_X1  g0924(.A1(new_n305), .A2(new_n396), .ZN(new_n1125));
  XOR2_X1   g0925(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1126));
  XOR2_X1   g0926(.A(new_n1125), .B(new_n1126), .Z(new_n1127));
  NAND2_X1  g0927(.A1(new_n301), .A2(new_n842), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(new_n1127), .B(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(new_n771), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n260), .B1(new_n740), .B2(new_n403), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n1069), .A2(new_n491), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n743), .A2(new_n217), .ZN(new_n1134));
  NOR4_X1   g0934(.A1(new_n1132), .A2(new_n1133), .A3(new_n1134), .A4(new_n995), .ZN(new_n1135));
  OAI221_X1 g0935(.A(new_n364), .B1(new_n497), .B2(new_n736), .C1(new_n729), .C2(new_n241), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(new_n749), .B2(G283), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n1135), .B(new_n1137), .C1(new_n243), .C2(new_n811), .ZN(new_n1138));
  XOR2_X1   g0938(.A(new_n1138), .B(KEYINPUT58), .Z(new_n1139));
  OAI21_X1  g0939(.A(new_n277), .B1(new_n314), .B2(G41), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n754), .A2(G132), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n728), .A2(G128), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n732), .A2(G125), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n765), .A2(new_n1114), .B1(new_n752), .B2(G150), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1141), .A2(new_n1142), .A3(new_n1143), .A4(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1145), .B1(G137), .B2(new_n739), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT59), .ZN(new_n1147));
  AOI21_X1  g0947(.A(G33), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n744), .A2(new_n762), .ZN(new_n1149));
  AOI21_X1  g0949(.A(G41), .B1(new_n761), .B2(G124), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1148), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1140), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n726), .B1(new_n1139), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n807), .A2(new_n277), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n1131), .A2(new_n722), .A3(new_n1154), .A4(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1080), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1102), .A2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n670), .B1(new_n890), .B2(new_n892), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n882), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT117), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n882), .A2(new_n1160), .A3(KEYINPUT117), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1163), .A2(new_n1164), .A3(new_n1129), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1130), .A2(KEYINPUT117), .A3(new_n882), .A4(new_n1160), .ZN(new_n1166));
  AND3_X1   g0966(.A1(new_n1165), .A2(new_n921), .A3(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n921), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1159), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT57), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n678), .A2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1157), .B1(new_n1169), .B2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1080), .B1(new_n1101), .B2(new_n1091), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n677), .A2(new_n1170), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n967), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT118), .ZN(new_n1176));
  AND3_X1   g0976(.A1(new_n882), .A2(new_n1160), .A3(KEYINPUT117), .ZN(new_n1177));
  AOI21_X1  g0977(.A(KEYINPUT117), .B1(new_n882), .B2(new_n1160), .ZN(new_n1178));
  NOR3_X1   g0978(.A1(new_n1177), .A2(new_n1178), .A3(new_n1130), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1166), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n920), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1165), .A2(new_n921), .A3(new_n1166), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1176), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(new_n1176), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1175), .B1(new_n1183), .B2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1172), .A2(new_n1186), .ZN(G375));
  NAND3_X1  g0987(.A1(new_n1086), .A2(new_n1080), .A3(new_n1090), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1092), .A2(new_n983), .A3(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n967), .B1(new_n1086), .B2(new_n1090), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n910), .A2(new_n772), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n739), .A2(G107), .B1(G294), .B2(new_n732), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1192), .B1(new_n243), .B2(new_n1069), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(new_n1193), .B(KEYINPUT120), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1018), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n728), .A2(G283), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1195), .A2(new_n1196), .A3(new_n988), .ZN(new_n1197));
  AOI211_X1 g0997(.A(new_n256), .B(new_n1197), .C1(G97), .C2(new_n765), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1194), .B(new_n1198), .C1(new_n734), .C2(new_n748), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n736), .A2(new_n1112), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1134), .A2(new_n364), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(new_n1201), .B(KEYINPUT121), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n1200), .B(new_n1202), .C1(G50), .C2(new_n752), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1203), .B1(new_n289), .B2(new_n740), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(G128), .B2(new_n749), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(new_n1205), .B(KEYINPUT122), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n754), .A2(new_n1114), .B1(G132), .B2(new_n732), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1207), .B1(new_n810), .B2(new_n729), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1199), .B1(new_n1206), .B2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1191), .B1(new_n1209), .B2(new_n726), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n723), .B1(new_n211), .B2(new_n807), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(new_n1211), .B(KEYINPUT119), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1190), .B1(new_n1210), .B2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1189), .A2(new_n1213), .ZN(G381));
  AOI21_X1  g1014(.A(new_n1014), .B1(new_n966), .B2(new_n985), .ZN(new_n1215));
  NOR3_X1   g1015(.A1(G390), .A2(G396), .A3(G393), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(G381), .A2(G384), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(G375), .A2(G378), .ZN(new_n1218));
  AND4_X1   g1018(.A1(new_n1215), .A2(new_n1216), .A3(new_n1217), .A4(new_n1218), .ZN(new_n1219));
  AND2_X1   g1019(.A1(new_n1219), .A2(KEYINPUT123), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1219), .A2(KEYINPUT123), .ZN(new_n1221));
  OR2_X1    g1021(.A1(new_n1220), .A2(new_n1221), .ZN(G407));
  INV_X1    g1022(.A(G213), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n654), .A2(G213), .ZN(new_n1224));
  XOR2_X1   g1024(.A(new_n1224), .B(KEYINPUT124), .Z(new_n1225));
  NOR3_X1   g1025(.A1(G375), .A2(G378), .A3(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1223), .B1(new_n1226), .B2(KEYINPUT125), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n1227), .B1(KEYINPUT125), .B2(new_n1226), .C1(new_n1220), .C2(new_n1221), .ZN(G409));
  XOR2_X1   g1028(.A(G393), .B(G396), .Z(new_n1229));
  INV_X1    g1029(.A(KEYINPUT127), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1052), .A2(new_n1075), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1078), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1232), .B1(new_n1233), .B2(new_n677), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1231), .B1(G387), .B2(new_n1234), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1215), .A2(G390), .A3(new_n1229), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(G387), .A2(new_n1234), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1238), .A2(new_n1231), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1239), .A2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1225), .ZN(new_n1243));
  INV_X1    g1043(.A(G378), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1159), .A2(new_n983), .ZN(new_n1245));
  OAI21_X1  g1045(.A(KEYINPUT118), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1245), .B1(new_n1246), .B2(new_n1184), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(new_n721), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(new_n1156), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1244), .B1(new_n1247), .B2(new_n1250), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1172), .A2(new_n1186), .A3(G378), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1243), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT60), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n678), .B1(new_n1188), .B2(new_n1254), .ZN(new_n1255));
  OAI211_X1 g1055(.A(new_n1255), .B(new_n1092), .C1(new_n1254), .C2(new_n1188), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(new_n1213), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1257), .A2(new_n805), .A3(new_n829), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1256), .A2(G384), .A3(new_n1213), .ZN(new_n1259));
  AND2_X1   g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  AND2_X1   g1060(.A1(new_n1260), .A2(KEYINPUT63), .ZN(new_n1261));
  AOI21_X1  g1061(.A(KEYINPUT61), .B1(new_n1253), .B2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT63), .ZN(new_n1263));
  AND3_X1   g1063(.A1(new_n1172), .A2(new_n1186), .A3(G378), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1173), .A2(new_n984), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1265), .B1(new_n1183), .B2(new_n1185), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1157), .B1(new_n1248), .B2(new_n721), .ZN(new_n1267));
  AOI21_X1  g1067(.A(G378), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  OAI21_X1  g1068(.A(KEYINPUT126), .B1(new_n1264), .B2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT126), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1251), .A2(new_n1270), .A3(new_n1252), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1269), .A2(new_n1224), .A3(new_n1271), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1260), .A2(new_n1225), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n654), .A2(G213), .A3(G2897), .ZN(new_n1274));
  AOI22_X1  g1074(.A1(new_n1273), .A2(G2897), .B1(new_n1260), .B2(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1263), .B1(new_n1272), .B2(new_n1275), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1269), .A2(new_n1224), .A3(new_n1260), .A4(new_n1271), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  OAI211_X1 g1078(.A(new_n1242), .B(new_n1262), .C1(new_n1276), .C2(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1240), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1258), .A2(KEYINPUT62), .A3(new_n1259), .ZN(new_n1281));
  AOI211_X1 g1081(.A(new_n1243), .B(new_n1281), .C1(new_n1251), .C2(new_n1252), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT62), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1282), .B1(new_n1277), .B2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT61), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1275), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1285), .B1(new_n1286), .B2(new_n1253), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1280), .B1(new_n1284), .B2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1279), .A2(new_n1288), .ZN(G405));
  NAND2_X1  g1089(.A1(G375), .A2(new_n1244), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1290), .A2(new_n1252), .ZN(new_n1291));
  XNOR2_X1  g1091(.A(new_n1291), .B(new_n1260), .ZN(new_n1292));
  XNOR2_X1  g1092(.A(new_n1280), .B(new_n1292), .ZN(G402));
endmodule


