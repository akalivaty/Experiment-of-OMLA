

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588;

  NOR2_X1 U320 ( .A1(n472), .A2(n518), .ZN(n570) );
  XNOR2_X1 U321 ( .A(n371), .B(n444), .ZN(n372) );
  XNOR2_X1 U322 ( .A(n368), .B(n367), .ZN(n369) );
  NOR2_X1 U323 ( .A1(n476), .A2(n475), .ZN(n566) );
  XOR2_X1 U324 ( .A(n377), .B(n376), .Z(n528) );
  XOR2_X1 U325 ( .A(KEYINPUT48), .B(KEYINPUT64), .Z(n288) );
  XNOR2_X1 U326 ( .A(n366), .B(n365), .ZN(n368) );
  INV_X1 U327 ( .A(n442), .ZN(n446) );
  INV_X1 U328 ( .A(KEYINPUT98), .ZN(n404) );
  XNOR2_X1 U329 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U330 ( .A(n468), .B(n288), .ZN(n527) );
  XNOR2_X1 U331 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U332 ( .A(n373), .B(n372), .ZN(n375) );
  INV_X1 U333 ( .A(G190GAT), .ZN(n477) );
  XOR2_X1 U334 ( .A(n473), .B(KEYINPUT28), .Z(n530) );
  XOR2_X1 U335 ( .A(n348), .B(n347), .Z(n518) );
  XNOR2_X1 U336 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U337 ( .A(G50GAT), .B(KEYINPUT106), .ZN(n454) );
  XNOR2_X1 U338 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n452) );
  XNOR2_X1 U339 ( .A(n480), .B(n479), .ZN(G1351GAT) );
  XNOR2_X1 U340 ( .A(n455), .B(n454), .ZN(G1331GAT) );
  XOR2_X1 U341 ( .A(KEYINPUT87), .B(KEYINPUT85), .Z(n290) );
  XNOR2_X1 U342 ( .A(KEYINPUT12), .B(KEYINPUT86), .ZN(n289) );
  XNOR2_X1 U343 ( .A(n290), .B(n289), .ZN(n308) );
  XOR2_X1 U344 ( .A(G155GAT), .B(G211GAT), .Z(n292) );
  XNOR2_X1 U345 ( .A(G22GAT), .B(G78GAT), .ZN(n291) );
  XNOR2_X1 U346 ( .A(n292), .B(n291), .ZN(n296) );
  XOR2_X1 U347 ( .A(KEYINPUT14), .B(KEYINPUT84), .Z(n294) );
  XNOR2_X1 U348 ( .A(G8GAT), .B(G64GAT), .ZN(n293) );
  XNOR2_X1 U349 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U350 ( .A(n296), .B(n295), .Z(n306) );
  XNOR2_X1 U351 ( .A(G15GAT), .B(G1GAT), .ZN(n297) );
  XNOR2_X1 U352 ( .A(n297), .B(KEYINPUT71), .ZN(n427) );
  XOR2_X1 U353 ( .A(n427), .B(KEYINPUT15), .Z(n299) );
  NAND2_X1 U354 ( .A1(G231GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U355 ( .A(n299), .B(n298), .ZN(n304) );
  XOR2_X1 U356 ( .A(G183GAT), .B(KEYINPUT83), .Z(n384) );
  XNOR2_X1 U357 ( .A(G57GAT), .B(KEYINPUT74), .ZN(n300) );
  XNOR2_X1 U358 ( .A(n300), .B(KEYINPUT13), .ZN(n438) );
  XOR2_X1 U359 ( .A(n384), .B(n438), .Z(n302) );
  XNOR2_X1 U360 ( .A(G71GAT), .B(G127GAT), .ZN(n301) );
  XNOR2_X1 U361 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U362 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U363 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U364 ( .A(n308), .B(n307), .Z(n483) );
  INV_X1 U365 ( .A(n483), .ZN(n581) );
  XOR2_X1 U366 ( .A(KEYINPUT11), .B(KEYINPUT81), .Z(n310) );
  XNOR2_X1 U367 ( .A(KEYINPUT9), .B(KEYINPUT65), .ZN(n309) );
  XNOR2_X1 U368 ( .A(n310), .B(n309), .ZN(n313) );
  XOR2_X1 U369 ( .A(G85GAT), .B(G92GAT), .Z(n312) );
  XNOR2_X1 U370 ( .A(G99GAT), .B(G106GAT), .ZN(n311) );
  XNOR2_X1 U371 ( .A(n312), .B(n311), .ZN(n439) );
  XOR2_X1 U372 ( .A(n313), .B(n439), .Z(n315) );
  XOR2_X1 U373 ( .A(G190GAT), .B(G134GAT), .Z(n366) );
  XOR2_X1 U374 ( .A(G218GAT), .B(G162GAT), .Z(n350) );
  XNOR2_X1 U375 ( .A(n366), .B(n350), .ZN(n314) );
  XNOR2_X1 U376 ( .A(n315), .B(n314), .ZN(n319) );
  XOR2_X1 U377 ( .A(KEYINPUT10), .B(KEYINPUT67), .Z(n317) );
  NAND2_X1 U378 ( .A1(G232GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U379 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U380 ( .A(n319), .B(n318), .Z(n325) );
  XNOR2_X1 U381 ( .A(G36GAT), .B(KEYINPUT8), .ZN(n320) );
  XNOR2_X1 U382 ( .A(n320), .B(G29GAT), .ZN(n321) );
  XOR2_X1 U383 ( .A(n321), .B(KEYINPUT7), .Z(n323) );
  XNOR2_X1 U384 ( .A(G43GAT), .B(G50GAT), .ZN(n322) );
  XNOR2_X1 U385 ( .A(n323), .B(n322), .ZN(n431) );
  XNOR2_X1 U386 ( .A(n431), .B(KEYINPUT80), .ZN(n324) );
  XNOR2_X1 U387 ( .A(n325), .B(n324), .ZN(n556) );
  XOR2_X1 U388 ( .A(KEYINPUT82), .B(n556), .Z(n538) );
  XNOR2_X1 U389 ( .A(KEYINPUT36), .B(n538), .ZN(n584) );
  XOR2_X1 U390 ( .A(KEYINPUT6), .B(G57GAT), .Z(n327) );
  XNOR2_X1 U391 ( .A(G1GAT), .B(G148GAT), .ZN(n326) );
  XNOR2_X1 U392 ( .A(n327), .B(n326), .ZN(n348) );
  XOR2_X1 U393 ( .A(G85GAT), .B(G134GAT), .Z(n329) );
  XNOR2_X1 U394 ( .A(G141GAT), .B(G120GAT), .ZN(n328) );
  XNOR2_X1 U395 ( .A(n329), .B(n328), .ZN(n331) );
  XOR2_X1 U396 ( .A(G29GAT), .B(G162GAT), .Z(n330) );
  XNOR2_X1 U397 ( .A(n331), .B(n330), .ZN(n344) );
  XNOR2_X1 U398 ( .A(KEYINPUT5), .B(KEYINPUT1), .ZN(n332) );
  XNOR2_X1 U399 ( .A(n332), .B(KEYINPUT4), .ZN(n333) );
  XOR2_X1 U400 ( .A(n333), .B(KEYINPUT91), .Z(n342) );
  INV_X1 U401 ( .A(G127GAT), .ZN(n334) );
  NAND2_X1 U402 ( .A1(n334), .A2(KEYINPUT0), .ZN(n337) );
  INV_X1 U403 ( .A(KEYINPUT0), .ZN(n335) );
  NAND2_X1 U404 ( .A1(G127GAT), .A2(n335), .ZN(n336) );
  NAND2_X1 U405 ( .A1(n337), .A2(n336), .ZN(n339) );
  XNOR2_X1 U406 ( .A(G113GAT), .B(KEYINPUT89), .ZN(n338) );
  XNOR2_X1 U407 ( .A(n339), .B(n338), .ZN(n367) );
  XNOR2_X1 U408 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n340) );
  XNOR2_X1 U409 ( .A(n340), .B(KEYINPUT2), .ZN(n349) );
  XNOR2_X1 U410 ( .A(n367), .B(n349), .ZN(n341) );
  XNOR2_X1 U411 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U412 ( .A(n344), .B(n343), .ZN(n346) );
  NAND2_X1 U413 ( .A1(G225GAT), .A2(G233GAT), .ZN(n345) );
  XNOR2_X1 U414 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U415 ( .A(n350), .B(n349), .Z(n352) );
  NAND2_X1 U416 ( .A1(G228GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U417 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U418 ( .A(n353), .B(KEYINPUT23), .Z(n356) );
  XNOR2_X1 U419 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n354) );
  XNOR2_X1 U420 ( .A(n354), .B(G211GAT), .ZN(n381) );
  XNOR2_X1 U421 ( .A(n381), .B(G204GAT), .ZN(n355) );
  XNOR2_X1 U422 ( .A(n356), .B(n355), .ZN(n360) );
  XOR2_X1 U423 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n358) );
  XNOR2_X1 U424 ( .A(G50GAT), .B(G106GAT), .ZN(n357) );
  XNOR2_X1 U425 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U426 ( .A(n360), .B(n359), .Z(n362) );
  XOR2_X1 U427 ( .A(G141GAT), .B(G22GAT), .Z(n415) );
  XOR2_X1 U428 ( .A(G148GAT), .B(G78GAT), .Z(n443) );
  XNOR2_X1 U429 ( .A(n415), .B(n443), .ZN(n361) );
  XNOR2_X1 U430 ( .A(n362), .B(n361), .ZN(n473) );
  XOR2_X1 U431 ( .A(KEYINPUT90), .B(KEYINPUT20), .Z(n364) );
  XNOR2_X1 U432 ( .A(G15GAT), .B(G183GAT), .ZN(n363) );
  XNOR2_X1 U433 ( .A(n364), .B(n363), .ZN(n377) );
  AND2_X1 U434 ( .A1(G227GAT), .A2(G233GAT), .ZN(n365) );
  XOR2_X1 U435 ( .A(G176GAT), .B(n369), .Z(n373) );
  XNOR2_X1 U436 ( .A(KEYINPUT17), .B(KEYINPUT19), .ZN(n370) );
  XNOR2_X1 U437 ( .A(n370), .B(KEYINPUT18), .ZN(n392) );
  XNOR2_X1 U438 ( .A(G169GAT), .B(n392), .ZN(n371) );
  XOR2_X1 U439 ( .A(G120GAT), .B(G71GAT), .Z(n444) );
  XOR2_X1 U440 ( .A(G43GAT), .B(G99GAT), .Z(n374) );
  XNOR2_X1 U441 ( .A(n375), .B(n374), .ZN(n376) );
  NOR2_X1 U442 ( .A1(n473), .A2(n528), .ZN(n378) );
  XNOR2_X1 U443 ( .A(n378), .B(KEYINPUT26), .ZN(n571) );
  XOR2_X1 U444 ( .A(G64GAT), .B(KEYINPUT78), .Z(n380) );
  XNOR2_X1 U445 ( .A(G176GAT), .B(G204GAT), .ZN(n379) );
  XNOR2_X1 U446 ( .A(n380), .B(n379), .ZN(n442) );
  XNOR2_X1 U447 ( .A(n381), .B(n442), .ZN(n396) );
  XOR2_X1 U448 ( .A(KEYINPUT95), .B(KEYINPUT93), .Z(n383) );
  XNOR2_X1 U449 ( .A(G190GAT), .B(G92GAT), .ZN(n382) );
  XNOR2_X1 U450 ( .A(n383), .B(n382), .ZN(n388) );
  XOR2_X1 U451 ( .A(n384), .B(G218GAT), .Z(n386) );
  XOR2_X1 U452 ( .A(G169GAT), .B(G8GAT), .Z(n414) );
  XNOR2_X1 U453 ( .A(G36GAT), .B(n414), .ZN(n385) );
  XNOR2_X1 U454 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U455 ( .A(n388), .B(n387), .Z(n390) );
  NAND2_X1 U456 ( .A1(G226GAT), .A2(G233GAT), .ZN(n389) );
  XNOR2_X1 U457 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U458 ( .A(n391), .B(KEYINPUT94), .Z(n394) );
  XNOR2_X1 U459 ( .A(n392), .B(KEYINPUT92), .ZN(n393) );
  XNOR2_X1 U460 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U461 ( .A(n396), .B(n395), .ZN(n520) );
  XNOR2_X1 U462 ( .A(n520), .B(KEYINPUT27), .ZN(n406) );
  AND2_X1 U463 ( .A1(n571), .A2(n406), .ZN(n397) );
  XNOR2_X1 U464 ( .A(KEYINPUT96), .B(n397), .ZN(n402) );
  NAND2_X1 U465 ( .A1(n520), .A2(n528), .ZN(n398) );
  NAND2_X1 U466 ( .A1(n398), .A2(n473), .ZN(n399) );
  XNOR2_X1 U467 ( .A(n399), .B(KEYINPUT97), .ZN(n400) );
  XOR2_X1 U468 ( .A(KEYINPUT25), .B(n400), .Z(n401) );
  NOR2_X1 U469 ( .A1(n402), .A2(n401), .ZN(n403) );
  NOR2_X1 U470 ( .A1(n518), .A2(n403), .ZN(n405) );
  XNOR2_X1 U471 ( .A(n405), .B(n404), .ZN(n409) );
  NAND2_X1 U472 ( .A1(n518), .A2(n406), .ZN(n526) );
  NOR2_X1 U473 ( .A1(n530), .A2(n526), .ZN(n407) );
  INV_X1 U474 ( .A(n528), .ZN(n476) );
  NAND2_X1 U475 ( .A1(n407), .A2(n476), .ZN(n408) );
  NAND2_X1 U476 ( .A1(n409), .A2(n408), .ZN(n486) );
  NAND2_X1 U477 ( .A1(n584), .A2(n486), .ZN(n410) );
  NOR2_X1 U478 ( .A1(n581), .A2(n410), .ZN(n411) );
  XNOR2_X1 U479 ( .A(n411), .B(KEYINPUT37), .ZN(n517) );
  XOR2_X1 U480 ( .A(KEYINPUT30), .B(KEYINPUT70), .Z(n413) );
  XNOR2_X1 U481 ( .A(KEYINPUT69), .B(KEYINPUT29), .ZN(n412) );
  XNOR2_X1 U482 ( .A(n413), .B(n412), .ZN(n419) );
  XOR2_X1 U483 ( .A(G197GAT), .B(G113GAT), .Z(n417) );
  XNOR2_X1 U484 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U485 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U486 ( .A(n419), .B(n418), .Z(n421) );
  NAND2_X1 U487 ( .A1(G229GAT), .A2(G233GAT), .ZN(n420) );
  XNOR2_X1 U488 ( .A(n421), .B(n420), .ZN(n423) );
  INV_X1 U489 ( .A(KEYINPUT72), .ZN(n422) );
  NAND2_X1 U490 ( .A1(n423), .A2(n422), .ZN(n426) );
  INV_X1 U491 ( .A(n423), .ZN(n424) );
  NAND2_X1 U492 ( .A1(n424), .A2(KEYINPUT72), .ZN(n425) );
  NAND2_X1 U493 ( .A1(n426), .A2(n425), .ZN(n429) );
  XNOR2_X1 U494 ( .A(n427), .B(KEYINPUT68), .ZN(n428) );
  XNOR2_X1 U495 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U496 ( .A(n431), .B(n430), .Z(n505) );
  XOR2_X1 U497 ( .A(KEYINPUT73), .B(n505), .Z(n531) );
  XOR2_X1 U498 ( .A(KEYINPUT76), .B(KEYINPUT75), .Z(n433) );
  XNOR2_X1 U499 ( .A(KEYINPUT31), .B(KEYINPUT32), .ZN(n432) );
  XNOR2_X1 U500 ( .A(n433), .B(n432), .ZN(n450) );
  XOR2_X1 U501 ( .A(KEYINPUT33), .B(KEYINPUT79), .Z(n435) );
  NAND2_X1 U502 ( .A1(G230GAT), .A2(G233GAT), .ZN(n434) );
  XNOR2_X1 U503 ( .A(n435), .B(n434), .ZN(n437) );
  INV_X1 U504 ( .A(KEYINPUT77), .ZN(n436) );
  XNOR2_X1 U505 ( .A(n437), .B(n436), .ZN(n441) );
  XNOR2_X1 U506 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U507 ( .A(n441), .B(n440), .ZN(n448) );
  XNOR2_X1 U508 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U509 ( .A(n450), .B(n449), .Z(n576) );
  OR2_X1 U510 ( .A1(n531), .A2(n576), .ZN(n488) );
  NOR2_X1 U511 ( .A1(n517), .A2(n488), .ZN(n451) );
  XNOR2_X1 U512 ( .A(KEYINPUT38), .B(n451), .ZN(n503) );
  NAND2_X1 U513 ( .A1(n503), .A2(n528), .ZN(n453) );
  XNOR2_X1 U514 ( .A(n453), .B(n452), .ZN(G1330GAT) );
  NAND2_X1 U515 ( .A1(n503), .A2(n530), .ZN(n455) );
  XOR2_X1 U516 ( .A(KEYINPUT54), .B(KEYINPUT117), .Z(n471) );
  XOR2_X1 U517 ( .A(KEYINPUT66), .B(KEYINPUT110), .Z(n456) );
  XNOR2_X1 U518 ( .A(KEYINPUT45), .B(n456), .ZN(n458) );
  NAND2_X1 U519 ( .A1(n581), .A2(n584), .ZN(n457) );
  XOR2_X1 U520 ( .A(n458), .B(n457), .Z(n459) );
  NOR2_X1 U521 ( .A1(n576), .A2(n459), .ZN(n460) );
  NAND2_X1 U522 ( .A1(n460), .A2(n531), .ZN(n467) );
  INV_X1 U523 ( .A(KEYINPUT41), .ZN(n461) );
  XNOR2_X1 U524 ( .A(n461), .B(n576), .ZN(n548) );
  INV_X1 U525 ( .A(n505), .ZN(n573) );
  NAND2_X1 U526 ( .A1(n548), .A2(n573), .ZN(n462) );
  XNOR2_X1 U527 ( .A(n462), .B(KEYINPUT46), .ZN(n463) );
  AND2_X1 U528 ( .A1(n463), .A2(n556), .ZN(n464) );
  AND2_X1 U529 ( .A1(n483), .A2(n464), .ZN(n465) );
  XNOR2_X1 U530 ( .A(n465), .B(KEYINPUT47), .ZN(n466) );
  NAND2_X1 U531 ( .A1(n467), .A2(n466), .ZN(n468) );
  INV_X1 U532 ( .A(n527), .ZN(n469) );
  NAND2_X1 U533 ( .A1(n520), .A2(n469), .ZN(n470) );
  XNOR2_X1 U534 ( .A(n471), .B(n470), .ZN(n472) );
  NAND2_X1 U535 ( .A1(n473), .A2(n570), .ZN(n474) );
  XOR2_X1 U536 ( .A(KEYINPUT55), .B(n474), .Z(n475) );
  NAND2_X1 U537 ( .A1(n566), .A2(n538), .ZN(n480) );
  XOR2_X1 U538 ( .A(KEYINPUT120), .B(KEYINPUT58), .Z(n478) );
  XNOR2_X1 U539 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n481) );
  XNOR2_X1 U540 ( .A(n481), .B(KEYINPUT100), .ZN(n482) );
  XOR2_X1 U541 ( .A(KEYINPUT99), .B(n482), .Z(n490) );
  XNOR2_X1 U542 ( .A(KEYINPUT88), .B(KEYINPUT16), .ZN(n485) );
  NOR2_X1 U543 ( .A1(n538), .A2(n483), .ZN(n484) );
  XNOR2_X1 U544 ( .A(n485), .B(n484), .ZN(n487) );
  NAND2_X1 U545 ( .A1(n487), .A2(n486), .ZN(n507) );
  NOR2_X1 U546 ( .A1(n488), .A2(n507), .ZN(n497) );
  NAND2_X1 U547 ( .A1(n497), .A2(n518), .ZN(n489) );
  XNOR2_X1 U548 ( .A(n490), .B(n489), .ZN(G1324GAT) );
  XOR2_X1 U549 ( .A(G8GAT), .B(KEYINPUT101), .Z(n492) );
  NAND2_X1 U550 ( .A1(n497), .A2(n520), .ZN(n491) );
  XNOR2_X1 U551 ( .A(n492), .B(n491), .ZN(G1325GAT) );
  XOR2_X1 U552 ( .A(KEYINPUT35), .B(KEYINPUT103), .Z(n494) );
  NAND2_X1 U553 ( .A1(n497), .A2(n528), .ZN(n493) );
  XNOR2_X1 U554 ( .A(n494), .B(n493), .ZN(n496) );
  XOR2_X1 U555 ( .A(G15GAT), .B(KEYINPUT102), .Z(n495) );
  XNOR2_X1 U556 ( .A(n496), .B(n495), .ZN(G1326GAT) );
  NAND2_X1 U557 ( .A1(n497), .A2(n530), .ZN(n498) );
  XNOR2_X1 U558 ( .A(n498), .B(KEYINPUT104), .ZN(n499) );
  XNOR2_X1 U559 ( .A(G22GAT), .B(n499), .ZN(G1327GAT) );
  NAND2_X1 U560 ( .A1(n503), .A2(n518), .ZN(n502) );
  XNOR2_X1 U561 ( .A(G29GAT), .B(KEYINPUT105), .ZN(n500) );
  XNOR2_X1 U562 ( .A(n500), .B(KEYINPUT39), .ZN(n501) );
  XNOR2_X1 U563 ( .A(n502), .B(n501), .ZN(G1328GAT) );
  NAND2_X1 U564 ( .A1(n503), .A2(n520), .ZN(n504) );
  XNOR2_X1 U565 ( .A(n504), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U566 ( .A(KEYINPUT107), .B(KEYINPUT42), .Z(n509) );
  XNOR2_X1 U567 ( .A(n548), .B(KEYINPUT108), .ZN(n563) );
  NAND2_X1 U568 ( .A1(n563), .A2(n505), .ZN(n506) );
  XOR2_X1 U569 ( .A(KEYINPUT109), .B(n506), .Z(n516) );
  NOR2_X1 U570 ( .A1(n516), .A2(n507), .ZN(n513) );
  NAND2_X1 U571 ( .A1(n513), .A2(n518), .ZN(n508) );
  XNOR2_X1 U572 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U573 ( .A(G57GAT), .B(n510), .ZN(G1332GAT) );
  NAND2_X1 U574 ( .A1(n513), .A2(n520), .ZN(n511) );
  XNOR2_X1 U575 ( .A(n511), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U576 ( .A1(n513), .A2(n528), .ZN(n512) );
  XNOR2_X1 U577 ( .A(n512), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U578 ( .A(G78GAT), .B(KEYINPUT43), .Z(n515) );
  NAND2_X1 U579 ( .A1(n513), .A2(n530), .ZN(n514) );
  XNOR2_X1 U580 ( .A(n515), .B(n514), .ZN(G1335GAT) );
  NOR2_X1 U581 ( .A1(n517), .A2(n516), .ZN(n523) );
  NAND2_X1 U582 ( .A1(n518), .A2(n523), .ZN(n519) );
  XNOR2_X1 U583 ( .A(G85GAT), .B(n519), .ZN(G1336GAT) );
  NAND2_X1 U584 ( .A1(n523), .A2(n520), .ZN(n521) );
  XNOR2_X1 U585 ( .A(n521), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U586 ( .A1(n523), .A2(n528), .ZN(n522) );
  XNOR2_X1 U587 ( .A(n522), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U588 ( .A1(n523), .A2(n530), .ZN(n524) );
  XNOR2_X1 U589 ( .A(n524), .B(KEYINPUT44), .ZN(n525) );
  XNOR2_X1 U590 ( .A(G106GAT), .B(n525), .ZN(G1339GAT) );
  XOR2_X1 U591 ( .A(G113GAT), .B(KEYINPUT111), .Z(n533) );
  NOR2_X1 U592 ( .A1(n527), .A2(n526), .ZN(n544) );
  NAND2_X1 U593 ( .A1(n528), .A2(n544), .ZN(n529) );
  NOR2_X1 U594 ( .A1(n530), .A2(n529), .ZN(n539) );
  INV_X1 U595 ( .A(n531), .ZN(n558) );
  NAND2_X1 U596 ( .A1(n539), .A2(n558), .ZN(n532) );
  XNOR2_X1 U597 ( .A(n533), .B(n532), .ZN(G1340GAT) );
  XOR2_X1 U598 ( .A(G120GAT), .B(KEYINPUT49), .Z(n535) );
  NAND2_X1 U599 ( .A1(n539), .A2(n563), .ZN(n534) );
  XNOR2_X1 U600 ( .A(n535), .B(n534), .ZN(G1341GAT) );
  NAND2_X1 U601 ( .A1(n581), .A2(n539), .ZN(n536) );
  XNOR2_X1 U602 ( .A(n536), .B(KEYINPUT50), .ZN(n537) );
  XNOR2_X1 U603 ( .A(G127GAT), .B(n537), .ZN(G1342GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT112), .B(KEYINPUT51), .Z(n541) );
  NAND2_X1 U605 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U606 ( .A(n541), .B(n540), .ZN(n543) );
  XOR2_X1 U607 ( .A(G134GAT), .B(KEYINPUT113), .Z(n542) );
  XNOR2_X1 U608 ( .A(n543), .B(n542), .ZN(G1343GAT) );
  XOR2_X1 U609 ( .A(G141GAT), .B(KEYINPUT115), .Z(n547) );
  NAND2_X1 U610 ( .A1(n544), .A2(n571), .ZN(n545) );
  XNOR2_X1 U611 ( .A(KEYINPUT114), .B(n545), .ZN(n555) );
  INV_X1 U612 ( .A(n555), .ZN(n553) );
  NAND2_X1 U613 ( .A1(n553), .A2(n573), .ZN(n546) );
  XNOR2_X1 U614 ( .A(n547), .B(n546), .ZN(G1344GAT) );
  XNOR2_X1 U615 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n552) );
  XOR2_X1 U616 ( .A(KEYINPUT116), .B(KEYINPUT53), .Z(n550) );
  NAND2_X1 U617 ( .A1(n548), .A2(n553), .ZN(n549) );
  XNOR2_X1 U618 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n552), .B(n551), .ZN(G1345GAT) );
  NAND2_X1 U620 ( .A1(n553), .A2(n581), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n554), .B(G155GAT), .ZN(G1346GAT) );
  NOR2_X1 U622 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U623 ( .A(G162GAT), .B(n557), .Z(G1347GAT) );
  NAND2_X1 U624 ( .A1(n566), .A2(n558), .ZN(n559) );
  XNOR2_X1 U625 ( .A(G169GAT), .B(n559), .ZN(G1348GAT) );
  XOR2_X1 U626 ( .A(KEYINPUT57), .B(KEYINPUT119), .Z(n561) );
  XNOR2_X1 U627 ( .A(G176GAT), .B(KEYINPUT118), .ZN(n560) );
  XNOR2_X1 U628 ( .A(n561), .B(n560), .ZN(n562) );
  XOR2_X1 U629 ( .A(KEYINPUT56), .B(n562), .Z(n565) );
  NAND2_X1 U630 ( .A1(n566), .A2(n563), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(G1349GAT) );
  NAND2_X1 U632 ( .A1(n581), .A2(n566), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n567), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U634 ( .A(G197GAT), .B(KEYINPUT122), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n568), .B(KEYINPUT60), .ZN(n569) );
  XOR2_X1 U636 ( .A(KEYINPUT59), .B(n569), .Z(n575) );
  NAND2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n572), .B(KEYINPUT121), .ZN(n585) );
  NAND2_X1 U639 ( .A1(n585), .A2(n573), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(G1352GAT) );
  XOR2_X1 U641 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n578) );
  NAND2_X1 U642 ( .A1(n585), .A2(n576), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(n580) );
  XOR2_X1 U644 ( .A(G204GAT), .B(KEYINPUT123), .Z(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1353GAT) );
  XOR2_X1 U646 ( .A(G211GAT), .B(KEYINPUT125), .Z(n583) );
  NAND2_X1 U647 ( .A1(n585), .A2(n581), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(G1354GAT) );
  XOR2_X1 U649 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n587) );
  NAND2_X1 U650 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n587), .B(n586), .ZN(n588) );
  XOR2_X1 U652 ( .A(G218GAT), .B(n588), .Z(G1355GAT) );
endmodule

