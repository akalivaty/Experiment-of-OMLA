//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 1 1 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 0 0 1 0 0 1 0 1 1 1 0 1 0 1 1 1 1 0 0 1 0 1 1 0 1 0 0 0 0 1 0 0 1 1 1 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:36 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1289, new_n1290, new_n1291,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1361, new_n1362, new_n1363, new_n1364, new_n1365,
    new_n1366, new_n1367, new_n1368, new_n1369, new_n1370, new_n1371;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NOR2_X1   g0002(.A1(G58), .A2(G68), .ZN(new_n203));
  AND3_X1   g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n207));
  INV_X1    g0007(.A(G68), .ZN(new_n208));
  INV_X1    g0008(.A(G238), .ZN(new_n209));
  INV_X1    g0009(.A(G87), .ZN(new_n210));
  INV_X1    g0010(.A(G250), .ZN(new_n211));
  OAI221_X1 g0011(.A(new_n207), .B1(new_n208), .B2(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n206), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT66), .Z(new_n217));
  INV_X1    g0017(.A(KEYINPUT1), .ZN(new_n218));
  OR2_X1    g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n217), .A2(new_n218), .ZN(new_n220));
  INV_X1    g0020(.A(KEYINPUT65), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n221), .B1(new_n206), .B2(G13), .ZN(new_n222));
  INV_X1    g0022(.A(G13), .ZN(new_n223));
  NAND4_X1  g0023(.A1(new_n223), .A2(KEYINPUT65), .A3(G1), .A4(G20), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n225), .B(G250), .C1(G257), .C2(G264), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT0), .Z(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  INV_X1    g0028(.A(G20), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(G50), .B1(G58), .B2(G68), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n227), .B1(new_n230), .B2(new_n232), .ZN(new_n233));
  AND3_X1   g0033(.A1(new_n219), .A2(new_n220), .A3(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  INV_X1    g0035(.A(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XOR2_X1   g0043(.A(G68), .B(G77), .Z(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G58), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G107), .B(G116), .Z(new_n247));
  XNOR2_X1  g0047(.A(G87), .B(G97), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  INV_X1    g0050(.A(G169), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT13), .ZN(new_n252));
  INV_X1    g0052(.A(G274), .ZN(new_n253));
  AND2_X1   g0053(.A1(G1), .A2(G13), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G33), .A2(G41), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n253), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NOR2_X1   g0056(.A1(G41), .A2(G45), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n257), .A2(G1), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(KEYINPUT72), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT72), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n256), .A2(new_n261), .A3(new_n258), .ZN(new_n262));
  NAND2_X1  g0062(.A1(G33), .A2(G97), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n236), .A2(G1698), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n264), .B1(G226), .B2(G1698), .ZN(new_n265));
  AND2_X1   g0065(.A1(KEYINPUT3), .A2(G33), .ZN(new_n266));
  NOR2_X1   g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n263), .B1(new_n265), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n254), .A2(new_n255), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  AOI22_X1  g0071(.A1(new_n260), .A2(new_n262), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  OAI21_X1  g0072(.A(KEYINPUT67), .B1(new_n257), .B2(G1), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT67), .ZN(new_n274));
  INV_X1    g0074(.A(G1), .ZN(new_n275));
  OAI211_X1 g0075(.A(new_n274), .B(new_n275), .C1(G41), .C2(G45), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n273), .A2(new_n270), .A3(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT73), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND4_X1  g0079(.A1(new_n273), .A2(KEYINPUT73), .A3(new_n270), .A4(new_n276), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n279), .A2(G238), .A3(new_n280), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n252), .B1(new_n272), .B2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n272), .A2(new_n252), .A3(new_n281), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n251), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT14), .ZN(new_n286));
  INV_X1    g0086(.A(new_n284), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n287), .A2(new_n282), .ZN(new_n288));
  AOI22_X1  g0088(.A1(new_n285), .A2(new_n286), .B1(new_n288), .B2(G179), .ZN(new_n289));
  NOR3_X1   g0089(.A1(new_n285), .A2(KEYINPUT74), .A3(new_n286), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT74), .ZN(new_n291));
  OAI21_X1  g0091(.A(G169), .B1(new_n287), .B2(new_n282), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n291), .B1(new_n292), .B2(KEYINPUT14), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n289), .B1(new_n290), .B2(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n275), .A2(G13), .A3(G20), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(new_n208), .ZN(new_n297));
  XNOR2_X1  g0097(.A(new_n297), .B(KEYINPUT12), .ZN(new_n298));
  NAND3_X1  g0098(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(new_n228), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n296), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n275), .A2(G20), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n301), .A2(G68), .A3(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G33), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n304), .A2(G20), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n306), .A2(new_n202), .ZN(new_n307));
  NOR2_X1   g0107(.A1(G20), .A2(G33), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G50), .ZN(new_n310));
  OAI22_X1  g0110(.A1(new_n309), .A2(new_n310), .B1(new_n229), .B2(G68), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n300), .B1(new_n307), .B2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT11), .ZN(new_n313));
  OAI211_X1 g0113(.A(new_n298), .B(new_n303), .C1(new_n312), .C2(new_n313), .ZN(new_n314));
  AND2_X1   g0114(.A1(new_n312), .A2(new_n313), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n294), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n288), .A2(G190), .ZN(new_n319));
  OAI21_X1  g0119(.A(G200), .B1(new_n287), .B2(new_n282), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n319), .A2(new_n316), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n318), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g0122(.A(KEYINPUT3), .B(G33), .ZN(new_n323));
  INV_X1    g0123(.A(G1698), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n323), .A2(G222), .A3(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n323), .A2(G223), .A3(G1698), .ZN(new_n326));
  OAI211_X1 g0126(.A(new_n325), .B(new_n326), .C1(new_n202), .C2(new_n323), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(new_n271), .ZN(new_n328));
  INV_X1    g0128(.A(G226), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n259), .B1(new_n277), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(KEYINPUT68), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT68), .ZN(new_n332));
  OAI211_X1 g0132(.A(new_n332), .B(new_n259), .C1(new_n277), .C2(new_n329), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n328), .A2(new_n331), .A3(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT69), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n328), .A2(new_n331), .A3(KEYINPUT69), .A4(new_n333), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(G190), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n336), .A2(G200), .A3(new_n337), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT71), .ZN(new_n341));
  XNOR2_X1  g0141(.A(KEYINPUT8), .B(G58), .ZN(new_n342));
  INV_X1    g0142(.A(G150), .ZN(new_n343));
  OAI22_X1  g0143(.A1(new_n342), .A2(new_n306), .B1(new_n343), .B2(new_n309), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n229), .B1(new_n201), .B2(new_n203), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n300), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n296), .A2(new_n310), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n301), .A2(G50), .A3(new_n302), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  OR2_X1    g0149(.A1(new_n349), .A2(KEYINPUT9), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(KEYINPUT9), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n341), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n339), .A2(new_n340), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(KEYINPUT10), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT10), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n339), .A2(new_n355), .A3(new_n340), .A4(new_n352), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(G179), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n338), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n336), .A2(new_n251), .A3(new_n337), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n359), .A2(new_n349), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n357), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n342), .B1(new_n275), .B2(G20), .ZN(new_n363));
  AOI22_X1  g0163(.A1(new_n363), .A2(new_n301), .B1(new_n296), .B2(new_n342), .ZN(new_n364));
  INV_X1    g0164(.A(G58), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n365), .A2(new_n208), .ZN(new_n366));
  OAI21_X1  g0166(.A(G20), .B1(new_n366), .B2(new_n203), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n308), .A2(G159), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g0169(.A(KEYINPUT7), .B1(new_n268), .B2(new_n229), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT3), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(new_n304), .ZN(new_n372));
  NAND2_X1  g0172(.A1(KEYINPUT3), .A2(G33), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n372), .A2(KEYINPUT7), .A3(new_n229), .A4(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(G68), .B1(new_n370), .B2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT75), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n369), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n372), .A2(new_n229), .A3(new_n373), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT7), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n208), .B1(new_n381), .B2(new_n374), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(KEYINPUT75), .ZN(new_n383));
  AOI21_X1  g0183(.A(KEYINPUT16), .B1(new_n378), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n369), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n376), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT16), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n300), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n364), .B1(new_n384), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(KEYINPUT76), .ZN(new_n390));
  OAI211_X1 g0190(.A(G223), .B(new_n324), .C1(new_n266), .C2(new_n267), .ZN(new_n391));
  OAI211_X1 g0191(.A(G226), .B(G1698), .C1(new_n266), .C2(new_n267), .ZN(new_n392));
  NAND2_X1  g0192(.A1(G33), .A2(G87), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n391), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(new_n271), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n273), .A2(G232), .A3(new_n270), .A4(new_n276), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n259), .ZN(new_n398));
  NOR3_X1   g0198(.A1(new_n396), .A2(G179), .A3(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(KEYINPUT77), .B1(new_n396), .B2(new_n398), .ZN(new_n400));
  AND2_X1   g0200(.A1(new_n397), .A2(new_n259), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT77), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n401), .A2(new_n395), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n400), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n399), .B1(new_n404), .B2(new_n251), .ZN(new_n405));
  INV_X1    g0205(.A(new_n364), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n385), .B1(new_n382), .B2(KEYINPUT75), .ZN(new_n407));
  AOI211_X1 g0207(.A(new_n377), .B(new_n208), .C1(new_n381), .C2(new_n374), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n387), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n300), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n382), .A2(new_n369), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n410), .B1(new_n411), .B2(KEYINPUT16), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n406), .B1(new_n409), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT76), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n390), .A2(new_n405), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(KEYINPUT18), .ZN(new_n417));
  INV_X1    g0217(.A(G200), .ZN(new_n418));
  AND3_X1   g0218(.A1(new_n401), .A2(new_n395), .A3(new_n402), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n402), .B1(new_n401), .B2(new_n395), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n418), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NOR3_X1   g0221(.A1(new_n396), .A2(G190), .A3(new_n398), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  AND3_X1   g0224(.A1(new_n424), .A2(KEYINPUT17), .A3(new_n413), .ZN(new_n425));
  AOI21_X1  g0225(.A(KEYINPUT17), .B1(new_n424), .B2(new_n413), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT18), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n390), .A2(new_n415), .A3(new_n428), .A4(new_n405), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n210), .A2(KEYINPUT15), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT15), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(G87), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n430), .A2(new_n432), .A3(KEYINPUT70), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(KEYINPUT70), .B1(new_n430), .B2(new_n432), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(new_n305), .ZN(new_n437));
  INV_X1    g0237(.A(new_n342), .ZN(new_n438));
  AOI22_X1  g0238(.A1(new_n438), .A2(new_n308), .B1(G20), .B2(G77), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n410), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n301), .A2(G77), .A3(new_n302), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n441), .B1(G77), .B2(new_n295), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(G244), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n259), .B1(new_n277), .B2(new_n445), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n323), .A2(G238), .A3(G1698), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n323), .A2(G232), .A3(new_n324), .ZN(new_n448));
  INV_X1    g0248(.A(G107), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n447), .B(new_n448), .C1(new_n449), .C2(new_n323), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n446), .B1(new_n450), .B2(new_n271), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(new_n358), .ZN(new_n452));
  OR2_X1    g0252(.A1(new_n451), .A2(G169), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n444), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n451), .A2(G190), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n443), .B(new_n455), .C1(new_n418), .C2(new_n451), .ZN(new_n456));
  AND2_X1   g0256(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n417), .A2(new_n427), .A3(new_n429), .A4(new_n457), .ZN(new_n458));
  NOR3_X1   g0258(.A1(new_n322), .A2(new_n362), .A3(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT83), .ZN(new_n461));
  INV_X1    g0261(.A(G41), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n461), .A2(new_n462), .A3(KEYINPUT5), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT5), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n464), .B1(KEYINPUT83), .B2(G41), .ZN(new_n465));
  INV_X1    g0265(.A(G45), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n466), .A2(G1), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n463), .A2(new_n465), .A3(new_n467), .ZN(new_n468));
  AND2_X1   g0268(.A1(new_n468), .A2(new_n270), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(G257), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n256), .A2(new_n467), .A3(new_n465), .A4(new_n463), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  OAI211_X1 g0273(.A(G250), .B(G1698), .C1(new_n266), .C2(new_n267), .ZN(new_n474));
  NAND2_X1  g0274(.A1(G33), .A2(G283), .ZN(new_n475));
  OAI211_X1 g0275(.A(G244), .B(new_n324), .C1(new_n266), .C2(new_n267), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT4), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n474), .B(new_n475), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n476), .A2(KEYINPUT80), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT80), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n323), .A2(new_n480), .A3(G244), .A4(new_n324), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n479), .A2(new_n481), .A3(new_n477), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT81), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n478), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n479), .A2(new_n481), .A3(KEYINPUT81), .A4(new_n477), .ZN(new_n485));
  AOI211_X1 g0285(.A(KEYINPUT82), .B(new_n270), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT82), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n482), .A2(new_n483), .ZN(new_n488));
  INV_X1    g0288(.A(new_n478), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n488), .A2(new_n485), .A3(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n487), .B1(new_n490), .B2(new_n271), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n358), .B(new_n473), .C1(new_n486), .C2(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n472), .B1(new_n490), .B2(new_n271), .ZN(new_n493));
  OR2_X1    g0293(.A1(new_n493), .A2(G169), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT6), .ZN(new_n495));
  AND2_X1   g0295(.A1(G97), .A2(G107), .ZN(new_n496));
  NOR2_X1   g0296(.A1(G97), .A2(G107), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  AND2_X1   g0298(.A1(KEYINPUT78), .A2(G97), .ZN(new_n499));
  NOR2_X1   g0299(.A1(KEYINPUT78), .A2(G97), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n449), .A2(KEYINPUT6), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n498), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  AOI22_X1  g0303(.A1(new_n503), .A2(G20), .B1(G77), .B2(new_n308), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT79), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n449), .B1(new_n381), .B2(new_n374), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  AND2_X1   g0307(.A1(new_n506), .A2(new_n505), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n300), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n295), .A2(G97), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n304), .A2(G1), .ZN(new_n511));
  NOR3_X1   g0311(.A1(new_n296), .A2(new_n300), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n510), .B1(new_n512), .B2(G97), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n509), .A2(new_n513), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n514), .A2(KEYINPUT84), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT84), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n516), .B1(new_n509), .B2(new_n513), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n492), .B(new_n494), .C1(new_n515), .C2(new_n517), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n514), .B1(G190), .B2(new_n493), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n490), .A2(new_n271), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(KEYINPUT82), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n490), .A2(new_n487), .A3(new_n271), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n472), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n519), .B1(new_n523), .B2(new_n418), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n518), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n323), .A2(G238), .A3(new_n324), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n323), .A2(G244), .A3(G1698), .ZN(new_n527));
  NAND2_X1  g0327(.A1(G33), .A2(G116), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n271), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n270), .B(G250), .C1(G1), .C2(new_n466), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n256), .A2(new_n467), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n530), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(G200), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n430), .A2(new_n432), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT70), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n295), .B1(new_n539), .B2(new_n433), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT19), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n541), .B1(new_n501), .B2(new_n306), .ZN(new_n542));
  OR2_X1    g0342(.A1(KEYINPUT78), .A2(G97), .ZN(new_n543));
  NAND2_X1  g0343(.A1(KEYINPUT78), .A2(G97), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n543), .A2(new_n210), .A3(new_n449), .A4(new_n544), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n229), .B1(new_n263), .B2(new_n541), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n323), .A2(new_n229), .A3(G68), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n542), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n540), .B1(new_n549), .B2(new_n300), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n533), .B1(new_n529), .B2(new_n271), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(G190), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n512), .A2(G87), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n536), .A2(new_n550), .A3(new_n552), .A4(new_n553), .ZN(new_n554));
  AND3_X1   g0354(.A1(new_n539), .A2(KEYINPUT85), .A3(new_n433), .ZN(new_n555));
  AOI21_X1  g0355(.A(KEYINPUT85), .B1(new_n539), .B2(new_n433), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(new_n512), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n550), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n535), .A2(new_n251), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n551), .A2(new_n358), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT86), .ZN(new_n563));
  AND3_X1   g0363(.A1(new_n554), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n563), .B1(new_n554), .B2(new_n562), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n525), .A2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n528), .A2(G20), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT23), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n570), .B1(new_n229), .B2(G107), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n449), .A2(KEYINPUT23), .A3(G20), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n569), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n323), .A2(new_n229), .A3(G87), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(KEYINPUT22), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT22), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n323), .A2(new_n577), .A3(new_n229), .A4(G87), .ZN(new_n578));
  AOI211_X1 g0378(.A(KEYINPUT24), .B(new_n574), .C1(new_n576), .C2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT24), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n576), .A2(new_n578), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n580), .B1(new_n581), .B2(new_n573), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n300), .B1(new_n579), .B2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT25), .ZN(new_n584));
  NOR3_X1   g0384(.A1(new_n295), .A2(new_n584), .A3(G107), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n584), .B1(new_n295), .B2(G107), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n512), .A2(G107), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n323), .A2(G257), .A3(G1698), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n323), .A2(G250), .A3(new_n324), .ZN(new_n590));
  XNOR2_X1  g0390(.A(KEYINPUT88), .B(G294), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(G33), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n589), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n271), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n469), .A2(G264), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n594), .A2(G190), .A3(new_n471), .A4(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n594), .A2(new_n471), .A3(new_n595), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(G200), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n583), .A2(new_n588), .A3(new_n596), .A4(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n588), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n581), .A2(new_n573), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(KEYINPUT24), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n581), .A2(new_n580), .A3(new_n573), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n600), .B1(new_n604), .B2(new_n300), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n597), .A2(new_n251), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n606), .B1(G179), .B2(new_n597), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n599), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(G116), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n296), .A2(KEYINPUT87), .A3(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT87), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n611), .B1(new_n295), .B2(G116), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n512), .A2(G116), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n299), .A2(new_n228), .B1(G20), .B2(new_n609), .ZN(new_n614));
  AOI21_X1  g0414(.A(G33), .B1(new_n543), .B2(new_n544), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n475), .A2(new_n229), .ZN(new_n616));
  OAI211_X1 g0416(.A(KEYINPUT20), .B(new_n614), .C1(new_n615), .C2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n616), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n619), .B1(new_n501), .B2(G33), .ZN(new_n620));
  AOI21_X1  g0420(.A(KEYINPUT20), .B1(new_n620), .B2(new_n614), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n613), .B1(new_n618), .B2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n468), .A2(G270), .A3(new_n270), .ZN(new_n624));
  AND2_X1   g0424(.A1(new_n624), .A2(new_n471), .ZN(new_n625));
  OAI211_X1 g0425(.A(G264), .B(G1698), .C1(new_n266), .C2(new_n267), .ZN(new_n626));
  OAI211_X1 g0426(.A(G257), .B(new_n324), .C1(new_n266), .C2(new_n267), .ZN(new_n627));
  INV_X1    g0427(.A(G303), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n626), .B(new_n627), .C1(new_n628), .C2(new_n323), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(new_n271), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n625), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(G200), .ZN(new_n632));
  INV_X1    g0432(.A(G190), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n623), .B(new_n632), .C1(new_n633), .C2(new_n631), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n251), .B1(new_n625), .B2(new_n630), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(new_n622), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT21), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n624), .A2(new_n471), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n639), .B1(new_n271), .B2(new_n629), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n622), .A2(new_n640), .A3(G179), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n635), .A2(KEYINPUT21), .A3(new_n622), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n634), .A2(new_n638), .A3(new_n641), .A4(new_n642), .ZN(new_n643));
  NOR4_X1   g0443(.A1(new_n460), .A2(new_n568), .A3(new_n608), .A4(new_n643), .ZN(G372));
  OAI21_X1  g0444(.A(new_n251), .B1(new_n419), .B2(new_n420), .ZN(new_n645));
  INV_X1    g0445(.A(new_n399), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n647), .A2(new_n413), .ZN(new_n648));
  XNOR2_X1  g0448(.A(new_n648), .B(new_n428), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n321), .A2(new_n452), .A3(new_n444), .A4(new_n453), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n283), .A2(G179), .A3(new_n284), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n651), .B1(new_n292), .B2(KEYINPUT14), .ZN(new_n652));
  OAI21_X1  g0452(.A(KEYINPUT74), .B1(new_n285), .B2(new_n286), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n292), .A2(new_n291), .A3(KEYINPUT14), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n652), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n650), .B1(new_n655), .B2(new_n316), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n649), .B1(new_n656), .B2(new_n427), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT90), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n357), .B1(new_n657), .B2(new_n658), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n361), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n642), .A2(new_n641), .ZN(new_n663));
  AOI21_X1  g0463(.A(KEYINPUT21), .B1(new_n635), .B2(new_n622), .ZN(new_n664));
  OAI21_X1  g0464(.A(KEYINPUT89), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT89), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n638), .A2(new_n666), .A3(new_n641), .A4(new_n642), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n607), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n583), .A2(new_n588), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  AND2_X1   g0472(.A1(new_n554), .A2(new_n562), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n673), .A2(new_n599), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n672), .A2(new_n524), .A3(new_n518), .A4(new_n674), .ZN(new_n675));
  AND3_X1   g0475(.A1(new_n514), .A2(new_n554), .A3(new_n562), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT26), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n676), .A2(new_n677), .A3(new_n492), .A4(new_n494), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n678), .A2(new_n562), .ZN(new_n679));
  OAI21_X1  g0479(.A(KEYINPUT26), .B1(new_n518), .B2(new_n566), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n675), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n459), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n662), .A2(new_n682), .ZN(G369));
  NAND3_X1  g0483(.A1(new_n275), .A2(new_n229), .A3(G13), .ZN(new_n684));
  OR2_X1    g0484(.A1(new_n684), .A2(KEYINPUT27), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(KEYINPUT27), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n685), .A2(G213), .A3(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(G343), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n622), .A2(new_n689), .ZN(new_n690));
  OR3_X1    g0490(.A1(new_n668), .A2(KEYINPUT91), .A3(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n663), .A2(new_n664), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n692), .A2(new_n634), .A3(new_n690), .ZN(new_n693));
  OAI211_X1 g0493(.A(KEYINPUT91), .B(new_n693), .C1(new_n668), .C2(new_n690), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n691), .A2(G330), .A3(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT92), .ZN(new_n697));
  INV_X1    g0497(.A(new_n689), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n697), .B1(new_n671), .B2(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n605), .A2(new_n607), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n700), .A2(KEYINPUT92), .A3(new_n689), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  OAI211_X1 g0502(.A(new_n671), .B(new_n599), .C1(new_n605), .C2(new_n698), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n696), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n692), .A2(new_n689), .ZN(new_n706));
  AOI22_X1  g0506(.A1(new_n704), .A2(new_n706), .B1(new_n700), .B2(new_n698), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n705), .A2(new_n707), .ZN(G399));
  INV_X1    g0508(.A(new_n225), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(G41), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n545), .A2(G116), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR3_X1   g0512(.A1(new_n710), .A2(new_n712), .A3(new_n275), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n713), .B1(new_n232), .B2(new_n710), .ZN(new_n714));
  XOR2_X1   g0514(.A(new_n714), .B(KEYINPUT28), .Z(new_n715));
  AND2_X1   g0515(.A1(new_n492), .A2(new_n494), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n554), .A2(new_n562), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(KEYINPUT86), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n554), .A2(new_n562), .A3(new_n563), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  OR2_X1    g0520(.A1(new_n515), .A2(new_n517), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n716), .A2(new_n720), .A3(new_n721), .A4(new_n677), .ZN(new_n722));
  INV_X1    g0522(.A(new_n562), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n676), .A2(new_n494), .A3(new_n492), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n723), .B1(new_n724), .B2(KEYINPUT26), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n671), .A2(new_n692), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n674), .A2(new_n726), .ZN(new_n727));
  OAI211_X1 g0527(.A(new_n722), .B(new_n725), .C1(new_n525), .C2(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n728), .A2(KEYINPUT29), .A3(new_n698), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(KEYINPUT94), .ZN(new_n730));
  AOI21_X1  g0530(.A(KEYINPUT29), .B1(new_n681), .B2(new_n698), .ZN(new_n731));
  OR2_X1    g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n597), .ZN(new_n733));
  OAI21_X1  g0533(.A(KEYINPUT93), .B1(new_n523), .B2(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n473), .B1(new_n486), .B2(new_n491), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT93), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n735), .A2(new_n736), .A3(new_n597), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n535), .A2(new_n631), .A3(new_n358), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n734), .A2(new_n737), .A3(new_n739), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n551), .A2(new_n595), .A3(new_n594), .ZN(new_n741));
  NOR3_X1   g0541(.A1(new_n741), .A2(new_n358), .A3(new_n631), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(new_n493), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT30), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n742), .A2(KEYINPUT30), .A3(new_n493), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n740), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT31), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n698), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  NOR3_X1   g0552(.A1(new_n608), .A2(new_n643), .A3(new_n689), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n753), .A2(new_n720), .A3(new_n518), .A4(new_n524), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n698), .B1(new_n740), .B2(new_n748), .ZN(new_n755));
  OAI211_X1 g0555(.A(new_n752), .B(new_n754), .C1(KEYINPUT31), .C2(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G330), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT94), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n728), .A2(new_n758), .A3(KEYINPUT29), .A4(new_n698), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n732), .A2(new_n757), .A3(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n715), .B1(new_n761), .B2(G1), .ZN(G364));
  NOR2_X1   g0562(.A1(new_n223), .A2(G20), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n275), .B1(new_n763), .B2(G45), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n710), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n695), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(G330), .B1(new_n691), .B2(new_n694), .ZN(new_n769));
  NOR2_X1   g0569(.A1(G13), .A2(G33), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(G20), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n773), .B1(new_n691), .B2(new_n694), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n228), .B1(G20), .B2(new_n251), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n229), .A2(G179), .ZN(new_n776));
  NOR2_X1   g0576(.A1(G190), .A2(G200), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(G159), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n776), .A2(new_n633), .A3(G200), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI22_X1  g0582(.A1(new_n780), .A2(KEYINPUT32), .B1(G107), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(G20), .A2(G179), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n785), .A2(G190), .A3(G200), .ZN(new_n786));
  INV_X1    g0586(.A(G97), .ZN(new_n787));
  NOR3_X1   g0587(.A1(new_n633), .A2(G179), .A3(G200), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(new_n229), .ZN(new_n789));
  OAI221_X1 g0589(.A(new_n783), .B1(new_n310), .B2(new_n786), .C1(new_n787), .C2(new_n789), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n776), .A2(G190), .A3(G200), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(new_n210), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n785), .A2(new_n633), .A3(G200), .ZN(new_n794));
  OAI221_X1 g0594(.A(new_n793), .B1(new_n208), .B2(new_n794), .C1(new_n780), .C2(KEYINPUT32), .ZN(new_n795));
  NOR3_X1   g0595(.A1(new_n784), .A2(G190), .A3(G200), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NOR3_X1   g0597(.A1(new_n784), .A2(new_n633), .A3(G200), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  OAI221_X1 g0599(.A(new_n323), .B1(new_n797), .B2(new_n202), .C1(new_n365), .C2(new_n799), .ZN(new_n800));
  NOR3_X1   g0600(.A1(new_n790), .A2(new_n795), .A3(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n794), .ZN(new_n802));
  INV_X1    g0602(.A(G317), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(KEYINPUT33), .ZN(new_n804));
  OR2_X1    g0604(.A1(new_n803), .A2(KEYINPUT33), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n802), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(G326), .ZN(new_n807));
  OAI221_X1 g0607(.A(new_n806), .B1(new_n628), .B2(new_n791), .C1(new_n807), .C2(new_n786), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n779), .A2(G329), .B1(G322), .B2(new_n798), .ZN(new_n809));
  INV_X1    g0609(.A(G311), .ZN(new_n810));
  OAI211_X1 g0610(.A(new_n809), .B(new_n268), .C1(new_n810), .C2(new_n797), .ZN(new_n811));
  INV_X1    g0611(.A(new_n591), .ZN(new_n812));
  INV_X1    g0612(.A(G283), .ZN(new_n813));
  OAI22_X1  g0613(.A1(new_n789), .A2(new_n812), .B1(new_n781), .B2(new_n813), .ZN(new_n814));
  NOR3_X1   g0614(.A1(new_n808), .A2(new_n811), .A3(new_n814), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n775), .B1(new_n801), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n232), .A2(new_n466), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n709), .A2(new_n323), .ZN(new_n818));
  OAI211_X1 g0618(.A(new_n817), .B(new_n818), .C1(new_n246), .C2(new_n466), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n709), .A2(new_n268), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n820), .A2(G355), .B1(new_n609), .B2(new_n709), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n772), .A2(new_n775), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n767), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n816), .A2(new_n824), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n768), .A2(new_n769), .B1(new_n774), .B2(new_n825), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n826), .B(KEYINPUT95), .ZN(G396));
  NAND2_X1  g0627(.A1(new_n681), .A2(new_n698), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n456), .B1(new_n443), .B2(new_n698), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(new_n454), .ZN(new_n830));
  OR2_X1    g0630(.A1(new_n454), .A2(new_n689), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n828), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n832), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n681), .A2(new_n698), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n766), .B1(new_n836), .B2(new_n757), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(new_n757), .B2(new_n836), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n775), .A2(new_n770), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n839), .B(KEYINPUT96), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n767), .B1(new_n841), .B2(new_n202), .ZN(new_n842));
  INV_X1    g0642(.A(new_n775), .ZN(new_n843));
  INV_X1    g0643(.A(new_n786), .ZN(new_n844));
  AOI22_X1  g0644(.A1(G87), .A2(new_n782), .B1(new_n844), .B2(G303), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n845), .B1(new_n449), .B2(new_n791), .ZN(new_n846));
  AOI22_X1  g0646(.A1(G116), .A2(new_n796), .B1(new_n798), .B2(G294), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n847), .B(new_n268), .C1(new_n810), .C2(new_n778), .ZN(new_n848));
  OAI22_X1  g0648(.A1(new_n789), .A2(new_n787), .B1(new_n794), .B2(new_n813), .ZN(new_n849));
  NOR3_X1   g0649(.A1(new_n846), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(G132), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n323), .B1(new_n778), .B2(new_n851), .C1(new_n208), .C2(new_n781), .ZN(new_n852));
  OAI22_X1  g0652(.A1(new_n789), .A2(new_n365), .B1(new_n791), .B2(new_n310), .ZN(new_n853));
  AOI22_X1  g0653(.A1(G143), .A2(new_n798), .B1(new_n796), .B2(G159), .ZN(new_n854));
  INV_X1    g0654(.A(G137), .ZN(new_n855));
  OAI221_X1 g0655(.A(new_n854), .B1(new_n855), .B2(new_n786), .C1(new_n343), .C2(new_n794), .ZN(new_n856));
  XNOR2_X1  g0656(.A(new_n856), .B(KEYINPUT97), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT34), .ZN(new_n858));
  AOI211_X1 g0658(.A(new_n852), .B(new_n853), .C1(new_n857), .C2(new_n858), .ZN(new_n859));
  OR2_X1    g0659(.A1(new_n857), .A2(new_n858), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n850), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  OAI221_X1 g0661(.A(new_n842), .B1(new_n843), .B2(new_n861), .C1(new_n834), .C2(new_n771), .ZN(new_n862));
  AND2_X1   g0662(.A1(new_n838), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(G384));
  OR2_X1    g0664(.A1(new_n503), .A2(KEYINPUT35), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n503), .A2(KEYINPUT35), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n865), .A2(G116), .A3(new_n230), .A4(new_n866), .ZN(new_n867));
  XOR2_X1   g0667(.A(new_n867), .B(KEYINPUT36), .Z(new_n868));
  NOR3_X1   g0668(.A1(new_n366), .A2(new_n231), .A3(new_n202), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT98), .ZN(new_n870));
  OR2_X1    g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n869), .A2(new_n870), .B1(G68), .B2(new_n201), .ZN(new_n872));
  AOI211_X1 g0672(.A(new_n275), .B(G13), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n868), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n759), .B1(new_n730), .B2(new_n731), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n459), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(new_n662), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT39), .ZN(new_n878));
  XOR2_X1   g0678(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n405), .A2(new_n389), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n424), .A2(new_n413), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT100), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n687), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n390), .A2(new_n415), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n883), .B1(new_n881), .B2(new_n882), .ZN(new_n888));
  OAI21_X1  g0688(.A(KEYINPUT37), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(KEYINPUT37), .B1(new_n424), .B2(new_n413), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n416), .A2(new_n886), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n409), .A2(new_n412), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n414), .B1(new_n893), .B2(new_n364), .ZN(new_n894));
  AOI211_X1 g0694(.A(KEYINPUT76), .B(new_n406), .C1(new_n409), .C2(new_n412), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n427), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n896), .B(new_n885), .C1(new_n649), .C2(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n880), .B1(new_n892), .B2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT38), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n411), .A2(KEYINPUT16), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n388), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n885), .B1(new_n902), .B2(new_n406), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n902), .A2(new_n406), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n882), .B(new_n903), .C1(new_n647), .C2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(KEYINPUT37), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n417), .A2(new_n429), .A3(new_n427), .ZN(new_n907));
  INV_X1    g0707(.A(new_n903), .ZN(new_n908));
  AOI221_X4 g0708(.A(new_n900), .B1(new_n891), .B2(new_n906), .C1(new_n907), .C2(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n878), .B1(new_n899), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n907), .A2(new_n908), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n891), .A2(new_n906), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n900), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n911), .A2(KEYINPUT38), .A3(new_n912), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n914), .A2(KEYINPUT39), .A3(new_n915), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n318), .A2(new_n689), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n910), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n321), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n317), .B(new_n689), .C1(new_n294), .C2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n317), .A2(new_n689), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n321), .B(new_n921), .C1(new_n655), .C2(new_n316), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n924), .B1(new_n835), .B2(new_n831), .ZN(new_n925));
  AOI21_X1  g0725(.A(KEYINPUT38), .B1(new_n911), .B2(new_n912), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n925), .B1(new_n909), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n649), .A2(new_n687), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n918), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n877), .B(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n832), .B1(new_n920), .B2(new_n922), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n756), .B(new_n931), .C1(new_n899), .C2(new_n909), .ZN(new_n932));
  AOI21_X1  g0732(.A(KEYINPUT40), .B1(new_n914), .B2(new_n915), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n923), .A2(new_n834), .ZN(new_n934));
  AOI21_X1  g0734(.A(KEYINPUT31), .B1(new_n749), .B2(new_n689), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n735), .A2(new_n597), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n738), .B1(new_n937), .B2(KEYINPUT93), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n747), .B1(new_n938), .B2(new_n737), .ZN(new_n939));
  INV_X1    g0739(.A(new_n751), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n754), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n934), .B1(new_n936), .B2(new_n942), .ZN(new_n943));
  AOI22_X1  g0743(.A1(KEYINPUT40), .A2(new_n932), .B1(new_n933), .B2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n756), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n944), .B1(new_n460), .B2(new_n945), .ZN(new_n946));
  AND2_X1   g0746(.A1(new_n933), .A2(new_n943), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT40), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n422), .B1(new_n404), .B2(new_n418), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n949), .A2(new_n389), .ZN(new_n950));
  OAI21_X1  g0750(.A(KEYINPUT100), .B1(new_n950), .B2(new_n648), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n951), .A2(new_n886), .A3(new_n884), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT37), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n949), .B2(new_n389), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n954), .B1(new_n896), .B2(new_n405), .ZN(new_n955));
  AOI22_X1  g0755(.A1(new_n952), .A2(KEYINPUT37), .B1(new_n886), .B2(new_n955), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n648), .B(KEYINPUT18), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n886), .B1(new_n957), .B2(new_n427), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n879), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(new_n915), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n948), .B1(new_n943), .B2(new_n960), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n459), .B(new_n756), .C1(new_n947), .C2(new_n961), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n946), .A2(new_n962), .A3(G330), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n930), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(new_n275), .B2(new_n763), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n930), .A2(new_n963), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n874), .B1(new_n965), .B2(new_n966), .ZN(G367));
  INV_X1    g0767(.A(KEYINPUT104), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n705), .A2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT45), .ZN(new_n971));
  INV_X1    g0771(.A(new_n707), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n514), .A2(new_n689), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n525), .A2(new_n973), .ZN(new_n974));
  OR2_X1    g0774(.A1(new_n716), .A2(new_n973), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n971), .B1(new_n972), .B2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n976), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n978), .A2(new_n707), .A3(KEYINPUT45), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n705), .A2(new_n968), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  NAND4_X1  g0783(.A1(new_n972), .A2(KEYINPUT102), .A3(KEYINPUT44), .A4(new_n976), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT102), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT44), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n978), .A2(new_n707), .B1(new_n985), .B2(new_n986), .ZN(new_n988));
  AND3_X1   g0788(.A1(new_n984), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n970), .B1(new_n983), .B2(new_n989), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n984), .A2(new_n987), .A3(new_n988), .ZN(new_n991));
  NAND4_X1  g0791(.A1(new_n991), .A2(new_n980), .A3(new_n969), .A4(new_n982), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT103), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(new_n704), .B2(new_n706), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(new_n696), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n995), .A2(new_n696), .ZN(new_n998));
  INV_X1    g0798(.A(new_n704), .ZN(new_n999));
  INV_X1    g0799(.A(new_n706), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n997), .A2(new_n998), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n998), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n999), .A2(new_n1000), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n1002), .A2(new_n1003), .A3(new_n996), .ZN(new_n1004));
  AND2_X1   g0804(.A1(new_n1001), .A2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n1005), .A2(new_n760), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n760), .B1(new_n993), .B2(new_n1006), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n710), .B(KEYINPUT41), .Z(new_n1008));
  OAI21_X1  g0808(.A(new_n764), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n550), .A2(new_n553), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1010), .A2(new_n689), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n562), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  OR2_X1    g0813(.A1(new_n1013), .A2(KEYINPUT101), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n1011), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n1013), .B(KEYINPUT101), .C1(new_n717), .C2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT43), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1017), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1020), .A2(KEYINPUT43), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1003), .A2(new_n978), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT42), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n978), .A2(new_n700), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n689), .B1(new_n1024), .B2(new_n518), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n1019), .B(new_n1021), .C1(new_n1023), .C2(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT42), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1022), .B(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1025), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1028), .A2(new_n1018), .A3(new_n1017), .A4(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1026), .A2(new_n1030), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n705), .A2(new_n976), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1031), .B(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1009), .A2(new_n1033), .ZN(new_n1034));
  XOR2_X1   g0834(.A(KEYINPUT105), .B(KEYINPUT46), .Z(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n791), .B2(new_n609), .ZN(new_n1036));
  XOR2_X1   g0836(.A(new_n1036), .B(KEYINPUT106), .Z(new_n1037));
  NOR2_X1   g0837(.A1(new_n791), .A2(new_n609), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n1038), .A2(KEYINPUT46), .B1(new_n802), .B2(new_n591), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n1040), .A2(KEYINPUT107), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(KEYINPUT107), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n268), .B1(new_n778), .B2(new_n803), .C1(new_n501), .C2(new_n781), .ZN(new_n1043));
  AND2_X1   g0843(.A1(new_n1043), .A2(KEYINPUT108), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n1043), .A2(KEYINPUT108), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(G283), .A2(new_n796), .B1(new_n798), .B2(G303), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1046), .B1(new_n449), .B2(new_n789), .C1(new_n810), .C2(new_n786), .ZN(new_n1047));
  NOR3_X1   g0847(.A1(new_n1044), .A2(new_n1045), .A3(new_n1047), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1041), .A2(new_n1042), .A3(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(G159), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n781), .A2(new_n202), .B1(new_n794), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n791), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1051), .B1(G58), .B2(new_n1052), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n789), .A2(new_n208), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(G143), .B2(new_n844), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n201), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n268), .B1(new_n1056), .B2(new_n796), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n779), .A2(G137), .B1(G150), .B2(new_n798), .ZN(new_n1058));
  NAND4_X1  g0858(.A1(new_n1053), .A2(new_n1055), .A3(new_n1057), .A4(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1049), .A2(new_n1059), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT47), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(new_n775), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n772), .B(new_n775), .C1(new_n436), .C2(new_n709), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n818), .A2(new_n242), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n767), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1062), .B(new_n1065), .C1(new_n773), .C2(new_n1020), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1034), .A2(new_n1066), .ZN(G387));
  INV_X1    g0867(.A(new_n710), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n1006), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1005), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1069), .B1(new_n761), .B2(new_n1070), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(G303), .A2(new_n796), .B1(new_n798), .B2(G317), .ZN(new_n1072));
  INV_X1    g0872(.A(G322), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n1072), .B1(new_n810), .B2(new_n794), .C1(new_n1073), .C2(new_n786), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT48), .ZN(new_n1075));
  OR2_X1    g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n789), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n1078), .A2(G283), .B1(new_n1052), .B2(new_n591), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1076), .A2(new_n1077), .A3(new_n1079), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1080), .B(KEYINPUT112), .ZN(new_n1081));
  OR2_X1    g0881(.A1(new_n1081), .A2(KEYINPUT49), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1081), .A2(KEYINPUT49), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n268), .B1(new_n778), .B2(new_n807), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(G116), .B2(new_n782), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1082), .A2(new_n1083), .A3(new_n1085), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n791), .A2(new_n202), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(G150), .B2(new_n779), .ZN(new_n1088));
  XOR2_X1   g0888(.A(new_n1088), .B(KEYINPUT111), .Z(new_n1089));
  OAI22_X1  g0889(.A1(new_n781), .A2(new_n787), .B1(new_n786), .B2(new_n1050), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n323), .B1(new_n797), .B2(new_n208), .C1(new_n310), .C2(new_n799), .ZN(new_n1091));
  AOI211_X1 g0891(.A(new_n1090), .B(new_n1091), .C1(new_n438), .C2(new_n802), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n1089), .B(new_n1092), .C1(new_n557), .C2(new_n789), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n843), .B1(new_n1086), .B2(new_n1093), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n820), .A2(new_n712), .B1(new_n449), .B2(new_n709), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n239), .A2(G45), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1096), .B(KEYINPUT109), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n342), .A2(G50), .ZN(new_n1098));
  XOR2_X1   g0898(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n1099));
  XNOR2_X1  g0899(.A(new_n1098), .B(new_n1099), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n711), .B(new_n466), .C1(new_n208), .C2(new_n202), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n818), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1095), .B1(new_n1097), .B2(new_n1102), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n767), .B(new_n1094), .C1(new_n823), .C2(new_n1103), .ZN(new_n1104));
  AND2_X1   g0904(.A1(new_n1104), .A2(KEYINPUT113), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1104), .A2(KEYINPUT113), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n704), .A2(new_n773), .ZN(new_n1107));
  NOR3_X1   g0907(.A1(new_n1105), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1108), .B1(new_n765), .B2(new_n1070), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1071), .A2(new_n1109), .ZN(G393));
  NAND2_X1  g0910(.A1(new_n993), .A2(new_n1006), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n990), .B(new_n992), .C1(new_n760), .C2(new_n1005), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1111), .A2(new_n710), .A3(new_n1112), .ZN(new_n1113));
  NOR3_X1   g0913(.A1(new_n249), .A2(new_n709), .A3(new_n323), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n823), .B1(new_n225), .B2(new_n501), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n799), .A2(new_n810), .B1(new_n786), .B2(new_n803), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1116), .B(KEYINPUT52), .ZN(new_n1117));
  INV_X1    g0917(.A(G294), .ZN(new_n1118));
  OAI221_X1 g0918(.A(new_n268), .B1(new_n778), .B2(new_n1073), .C1(new_n797), .C2(new_n1118), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n781), .A2(new_n449), .B1(new_n794), .B2(new_n628), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n789), .A2(new_n609), .B1(new_n791), .B2(new_n813), .ZN(new_n1121));
  NOR3_X1   g0921(.A1(new_n1119), .A2(new_n1120), .A3(new_n1121), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n799), .A2(new_n1050), .B1(new_n786), .B2(new_n343), .ZN(new_n1123));
  XOR2_X1   g0923(.A(KEYINPUT114), .B(KEYINPUT51), .Z(new_n1124));
  XNOR2_X1  g0924(.A(new_n1123), .B(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(G143), .ZN(new_n1126));
  OAI221_X1 g0926(.A(new_n323), .B1(new_n778), .B2(new_n1126), .C1(new_n797), .C2(new_n342), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n781), .A2(new_n210), .B1(new_n794), .B2(new_n201), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n789), .A2(new_n202), .B1(new_n791), .B2(new_n208), .ZN(new_n1129));
  NOR3_X1   g0929(.A1(new_n1127), .A2(new_n1128), .A3(new_n1129), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(new_n1117), .A2(new_n1122), .B1(new_n1125), .B2(new_n1130), .ZN(new_n1131));
  OAI221_X1 g0931(.A(new_n766), .B1(new_n1114), .B2(new_n1115), .C1(new_n1131), .C2(new_n843), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1132), .B1(new_n976), .B2(new_n772), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1133), .B1(new_n993), .B2(new_n765), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1113), .A2(new_n1134), .ZN(G390));
  NOR3_X1   g0935(.A1(new_n909), .A2(new_n926), .A3(new_n878), .ZN(new_n1136));
  AOI21_X1  g0936(.A(KEYINPUT39), .B1(new_n959), .B2(new_n915), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n1136), .A2(new_n1137), .B1(new_n925), .B2(new_n917), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n917), .B1(new_n959), .B2(new_n915), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n728), .A2(new_n698), .A3(new_n830), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n831), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1139), .B1(new_n1142), .B2(new_n924), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n756), .A2(G330), .A3(new_n834), .A4(new_n923), .ZN(new_n1144));
  AND3_X1   g0944(.A1(new_n1138), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1144), .B1(new_n1138), .B2(new_n1143), .ZN(new_n1146));
  NOR3_X1   g0946(.A1(new_n1145), .A2(new_n1146), .A3(new_n764), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n770), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n789), .A2(new_n1050), .B1(new_n794), .B2(new_n855), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(KEYINPUT54), .B(G143), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n1151), .A2(new_n796), .B1(G132), .B2(new_n798), .ZN(new_n1152));
  INV_X1    g0952(.A(G125), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1152), .B1(new_n1153), .B2(new_n778), .ZN(new_n1154));
  AOI211_X1 g0954(.A(new_n1149), .B(new_n1154), .C1(G128), .C2(new_n844), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1052), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT53), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1157), .B1(new_n791), .B2(new_n343), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n323), .B1(new_n781), .B2(new_n201), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT116), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n1156), .A2(new_n1158), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n1155), .B(new_n1161), .C1(new_n1160), .C2(new_n1159), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n789), .A2(new_n202), .B1(new_n799), .B2(new_n609), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(new_n1163), .B(KEYINPUT117), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n268), .B1(new_n778), .B2(new_n1118), .C1(new_n797), .C2(new_n501), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n449), .A2(new_n794), .B1(new_n786), .B2(new_n813), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n781), .A2(new_n208), .ZN(new_n1167));
  NOR4_X1   g0967(.A1(new_n1165), .A2(new_n1166), .A3(new_n792), .A4(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1164), .A2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n843), .B1(new_n1162), .B2(new_n1169), .ZN(new_n1170));
  AOI211_X1 g0970(.A(new_n767), .B(new_n1170), .C1(new_n342), .C2(new_n841), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(new_n1171), .B(KEYINPUT118), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1148), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  OAI21_X1  g0974(.A(KEYINPUT119), .B1(new_n1147), .B2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT119), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1138), .A2(new_n1143), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1144), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1138), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1176), .B(new_n1173), .C1(new_n1181), .C2(new_n764), .ZN(new_n1182));
  OAI211_X1 g0982(.A(G330), .B(new_n834), .C1(new_n935), .C2(new_n941), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1183), .A2(new_n924), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT115), .ZN(new_n1185));
  NAND4_X1  g0985(.A1(new_n1184), .A2(new_n1142), .A3(new_n1144), .A4(new_n1185), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1184), .A2(new_n1144), .A3(new_n1142), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1187), .A2(KEYINPUT115), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n1184), .A2(new_n1144), .B1(new_n831), .B2(new_n835), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1186), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n756), .A2(G330), .A3(new_n459), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n876), .A2(new_n662), .A3(new_n1191), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n1190), .A2(new_n1192), .B1(new_n1146), .B2(new_n1145), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1193), .A2(new_n710), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1191), .ZN(new_n1195));
  AOI211_X1 g0995(.A(new_n661), .B(new_n1195), .C1(new_n459), .C2(new_n875), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1196), .B(new_n1186), .C1(new_n1189), .C2(new_n1188), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1197), .A2(new_n1181), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1175), .B(new_n1182), .C1(new_n1194), .C2(new_n1198), .ZN(G378));
  INV_X1    g0999(.A(new_n349), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1200), .A2(new_n687), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n362), .A2(new_n1201), .ZN(new_n1202));
  AND2_X1   g1002(.A1(new_n362), .A2(new_n1201), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  OR3_X1    g1005(.A1(new_n1202), .A2(new_n1203), .A3(new_n1205), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1205), .B1(new_n1203), .B2(new_n1202), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(G330), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1209), .B1(new_n944), .B2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n929), .ZN(new_n1212));
  OAI211_X1 g1012(.A(G330), .B(new_n1208), .C1(new_n947), .C2(new_n961), .ZN(new_n1213));
  AND3_X1   g1013(.A1(new_n1211), .A2(new_n1212), .A3(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1212), .B1(new_n1211), .B2(new_n1213), .ZN(new_n1215));
  OAI21_X1  g1015(.A(KEYINPUT57), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1186), .ZN(new_n1218));
  AND2_X1   g1018(.A1(new_n1187), .A2(KEYINPUT115), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1189), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1218), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1192), .B1(new_n1217), .B2(new_n1221), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n710), .B1(new_n1216), .B2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1211), .A2(new_n1213), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1224), .A2(new_n929), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1211), .A2(new_n1213), .A3(new_n1212), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1196), .B1(new_n1181), .B2(new_n1190), .ZN(new_n1228));
  AOI21_X1  g1028(.A(KEYINPUT57), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  OR2_X1    g1029(.A1(new_n1223), .A2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1209), .A2(new_n770), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n766), .B1(new_n840), .B2(new_n1056), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(G58), .A2(new_n782), .B1(new_n844), .B2(G116), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1233), .B1(new_n787), .B2(new_n794), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n323), .A2(G41), .ZN(new_n1235));
  OAI221_X1 g1035(.A(new_n1235), .B1(new_n813), .B2(new_n778), .C1(new_n449), .C2(new_n799), .ZN(new_n1236));
  NOR4_X1   g1036(.A1(new_n1234), .A2(new_n1236), .A3(new_n1054), .A4(new_n1087), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1237), .B1(new_n557), .B2(new_n797), .ZN(new_n1238));
  XOR2_X1   g1038(.A(new_n1238), .B(KEYINPUT120), .Z(new_n1239));
  OR2_X1    g1039(.A1(new_n1239), .A2(KEYINPUT58), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(KEYINPUT58), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(G33), .A2(G41), .ZN(new_n1242));
  NOR3_X1   g1042(.A1(new_n1235), .A2(G50), .A3(new_n1242), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n1153), .A2(new_n786), .B1(new_n794), .B2(new_n851), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(G150), .B2(new_n1078), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(G128), .A2(new_n798), .B1(new_n796), .B2(G137), .ZN(new_n1246));
  OAI211_X1 g1046(.A(new_n1245), .B(new_n1246), .C1(new_n791), .C2(new_n1150), .ZN(new_n1247));
  OR2_X1    g1047(.A1(new_n1247), .A2(KEYINPUT59), .ZN(new_n1248));
  INV_X1    g1048(.A(G124), .ZN(new_n1249));
  OAI221_X1 g1049(.A(new_n1242), .B1(new_n778), .B2(new_n1249), .C1(new_n1050), .C2(new_n781), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1250), .B1(new_n1247), .B2(KEYINPUT59), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1243), .B1(new_n1248), .B2(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1240), .A2(new_n1241), .A3(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1232), .B1(new_n1253), .B2(new_n775), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n1227), .A2(new_n765), .B1(new_n1231), .B2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1230), .A2(new_n1255), .ZN(G375));
  NAND2_X1  g1056(.A1(new_n1190), .A2(new_n1192), .ZN(new_n1257));
  XOR2_X1   g1057(.A(new_n1008), .B(KEYINPUT121), .Z(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1197), .A2(new_n1257), .A3(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n924), .A2(new_n770), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n766), .B1(new_n840), .B2(G68), .ZN(new_n1262));
  OAI22_X1  g1062(.A1(new_n789), .A2(new_n310), .B1(new_n791), .B2(new_n1050), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1263), .B1(G132), .B2(new_n844), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n268), .B1(G137), .B2(new_n798), .ZN(new_n1265));
  AOI22_X1  g1065(.A1(new_n779), .A2(G128), .B1(G150), .B2(new_n796), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(G58), .A2(new_n782), .B1(new_n802), .B2(new_n1151), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1264), .A2(new_n1265), .A3(new_n1266), .A4(new_n1267), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n557), .A2(new_n789), .ZN(new_n1269));
  AOI22_X1  g1069(.A1(G77), .A2(new_n782), .B1(new_n802), .B2(G116), .ZN(new_n1270));
  AOI22_X1  g1070(.A1(G97), .A2(new_n1052), .B1(new_n844), .B2(G294), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n323), .B1(new_n779), .B2(G303), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(G107), .A2(new_n796), .B1(new_n798), .B2(G283), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1270), .A2(new_n1271), .A3(new_n1272), .A4(new_n1273), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1268), .B1(new_n1269), .B2(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1262), .B1(new_n1275), .B2(new_n775), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1261), .A2(new_n1276), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1277), .B1(new_n1190), .B2(new_n764), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1260), .A2(new_n1279), .ZN(G381));
  NOR4_X1   g1080(.A1(G390), .A2(G393), .A3(G396), .A4(G384), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1281), .A2(new_n1034), .A3(new_n1066), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1173), .B1(new_n1181), .B2(new_n764), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1068), .B1(new_n1197), .B2(new_n1181), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1217), .A2(new_n1221), .A3(new_n1196), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1283), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  OR4_X1    g1087(.A1(G375), .A2(new_n1282), .A3(G381), .A4(new_n1287), .ZN(G407));
  NAND2_X1  g1088(.A1(new_n688), .A2(G213), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1286), .A2(new_n1290), .ZN(new_n1291));
  OAI211_X1 g1091(.A(G407), .B(G213), .C1(G375), .C2(new_n1291), .ZN(G409));
  XNOR2_X1  g1092(.A(G393), .B(G396), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1066), .ZN(new_n1294));
  AOI221_X4 g1094(.A(new_n1294), .B1(new_n1113), .B2(new_n1134), .C1(new_n1009), .C2(new_n1033), .ZN(new_n1295));
  AOI21_X1  g1095(.A(G390), .B1(new_n1034), .B2(new_n1066), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1293), .B1(new_n1295), .B2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(G390), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1032), .ZN(new_n1299));
  XNOR2_X1  g1099(.A(new_n1031), .B(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1008), .ZN(new_n1301));
  AOI211_X1 g1101(.A(new_n760), .B(new_n1005), .C1(new_n990), .C2(new_n992), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1301), .B1(new_n1302), .B2(new_n760), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1300), .B1(new_n1303), .B2(new_n764), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1298), .B1(new_n1304), .B2(new_n1294), .ZN(new_n1305));
  INV_X1    g1105(.A(G396), .ZN(new_n1306));
  XNOR2_X1  g1106(.A(G393), .B(new_n1306), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1034), .A2(new_n1066), .A3(G390), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1305), .A2(new_n1307), .A3(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1297), .A2(new_n1309), .ZN(new_n1310));
  OAI211_X1 g1110(.A(G378), .B(new_n1255), .C1(new_n1223), .C2(new_n1229), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1312));
  NOR3_X1   g1112(.A1(new_n1312), .A2(new_n1222), .A3(new_n1258), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1231), .A2(new_n1254), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1314), .B1(new_n1312), .B2(new_n764), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1286), .B1(new_n1313), .B2(new_n1315), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1290), .B1(new_n1311), .B2(new_n1316), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1190), .A2(KEYINPUT60), .A3(new_n1192), .ZN(new_n1318));
  AND2_X1   g1118(.A1(new_n1318), .A2(new_n710), .ZN(new_n1319));
  OAI21_X1  g1119(.A(KEYINPUT60), .B1(new_n1190), .B2(new_n1192), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1320), .A2(new_n1257), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1278), .B1(new_n1319), .B2(new_n1321), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1322), .A2(G384), .ZN(new_n1323));
  AOI211_X1 g1123(.A(new_n863), .B(new_n1278), .C1(new_n1319), .C2(new_n1321), .ZN(new_n1324));
  NOR2_X1   g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  AND3_X1   g1125(.A1(new_n1317), .A2(KEYINPUT62), .A3(new_n1325), .ZN(new_n1326));
  XNOR2_X1  g1126(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1327), .B1(new_n1317), .B2(new_n1325), .ZN(new_n1328));
  NOR3_X1   g1128(.A1(new_n1326), .A2(new_n1328), .A3(KEYINPUT126), .ZN(new_n1329));
  XNOR2_X1  g1129(.A(KEYINPUT124), .B(KEYINPUT61), .ZN(new_n1330));
  AND2_X1   g1130(.A1(new_n1319), .A2(new_n1321), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n863), .B1(new_n1331), .B2(new_n1278), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1322), .A2(G384), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1290), .A2(G2897), .ZN(new_n1334));
  INV_X1    g1134(.A(new_n1334), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1332), .A2(new_n1333), .A3(new_n1335), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1334), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1336), .A2(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1311), .A2(new_n1316), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1339), .A2(new_n1289), .ZN(new_n1340));
  AOI21_X1  g1140(.A(new_n1330), .B1(new_n1338), .B2(new_n1340), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1339), .A2(new_n1325), .A3(new_n1289), .ZN(new_n1342));
  INV_X1    g1142(.A(new_n1327), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1342), .A2(KEYINPUT126), .A3(new_n1343), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1341), .A2(new_n1344), .ZN(new_n1345));
  OAI21_X1  g1145(.A(new_n1310), .B1(new_n1329), .B2(new_n1345), .ZN(new_n1346));
  NOR2_X1   g1146(.A1(new_n1338), .A2(KEYINPUT123), .ZN(new_n1347));
  INV_X1    g1147(.A(KEYINPUT123), .ZN(new_n1348));
  AOI21_X1  g1148(.A(new_n1348), .B1(new_n1336), .B2(new_n1337), .ZN(new_n1349));
  AND2_X1   g1149(.A1(new_n1317), .A2(KEYINPUT122), .ZN(new_n1350));
  NOR2_X1   g1150(.A1(new_n1317), .A2(KEYINPUT122), .ZN(new_n1351));
  OAI22_X1  g1151(.A1(new_n1347), .A2(new_n1349), .B1(new_n1350), .B2(new_n1351), .ZN(new_n1352));
  INV_X1    g1152(.A(KEYINPUT61), .ZN(new_n1353));
  AND3_X1   g1153(.A1(new_n1297), .A2(new_n1309), .A3(new_n1353), .ZN(new_n1354));
  NAND3_X1  g1154(.A1(new_n1317), .A2(KEYINPUT63), .A3(new_n1325), .ZN(new_n1355));
  AND2_X1   g1155(.A1(new_n1354), .A2(new_n1355), .ZN(new_n1356));
  INV_X1    g1156(.A(KEYINPUT63), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1342), .A2(new_n1357), .ZN(new_n1358));
  NAND3_X1  g1158(.A1(new_n1352), .A2(new_n1356), .A3(new_n1358), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1346), .A2(new_n1359), .ZN(G405));
  AOI21_X1  g1160(.A(new_n1287), .B1(new_n1230), .B2(new_n1255), .ZN(new_n1361));
  INV_X1    g1161(.A(new_n1311), .ZN(new_n1362));
  NOR2_X1   g1162(.A1(new_n1361), .A2(new_n1362), .ZN(new_n1363));
  INV_X1    g1163(.A(KEYINPUT127), .ZN(new_n1364));
  NAND3_X1  g1164(.A1(new_n1363), .A2(new_n1364), .A3(new_n1325), .ZN(new_n1365));
  INV_X1    g1165(.A(new_n1310), .ZN(new_n1366));
  NAND2_X1  g1166(.A1(new_n1325), .A2(new_n1364), .ZN(new_n1367));
  OAI21_X1  g1167(.A(KEYINPUT127), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1368));
  OAI211_X1 g1168(.A(new_n1367), .B(new_n1368), .C1(new_n1361), .C2(new_n1362), .ZN(new_n1369));
  AND3_X1   g1169(.A1(new_n1365), .A2(new_n1366), .A3(new_n1369), .ZN(new_n1370));
  AOI21_X1  g1170(.A(new_n1366), .B1(new_n1365), .B2(new_n1369), .ZN(new_n1371));
  NOR2_X1   g1171(.A1(new_n1370), .A2(new_n1371), .ZN(G402));
endmodule


