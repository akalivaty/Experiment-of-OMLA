//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 0 1 1 0 1 0 0 0 1 0 0 1 0 0 1 0 0 0 1 0 0 1 0 1 0 1 0 0 0 0 1 1 1 0 1 0 1 0 0 0 1 1 0 0 1 0 0 1 1 1 0 0 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:12 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n773,
    new_n774, new_n775, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n846, new_n847, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1033, new_n1034, new_n1035,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073;
  OAI21_X1  g000(.A(KEYINPUT74), .B1(G472), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  NOR3_X1   g002(.A1(KEYINPUT74), .A2(G472), .A3(G902), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G143), .ZN(new_n193));
  INV_X1    g007(.A(G143), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G146), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n193), .A2(new_n195), .A3(G128), .ZN(new_n196));
  XNOR2_X1  g010(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n197));
  OAI21_X1  g011(.A(KEYINPUT66), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  AND2_X1   g012(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n199));
  NOR2_X1   g013(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  XNOR2_X1  g015(.A(G143), .B(G146), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT66), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n201), .A2(new_n202), .A3(new_n203), .A4(G128), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n198), .A2(new_n204), .ZN(new_n205));
  XNOR2_X1  g019(.A(KEYINPUT67), .B(G128), .ZN(new_n206));
  INV_X1    g020(.A(new_n193), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n206), .B1(new_n201), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(new_n202), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n205), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(KEYINPUT69), .ZN(new_n212));
  INV_X1    g026(.A(G134), .ZN(new_n213));
  OAI21_X1  g027(.A(KEYINPUT11), .B1(new_n213), .B2(G137), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT11), .ZN(new_n215));
  INV_X1    g029(.A(G137), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n215), .A2(new_n216), .A3(G134), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n214), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G131), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n213), .A2(G137), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(KEYINPUT64), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT64), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n223), .A2(new_n213), .A3(G137), .ZN(new_n224));
  AOI22_X1  g038(.A1(new_n222), .A2(new_n224), .B1(G134), .B2(new_n216), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n221), .B1(new_n225), .B2(new_n219), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  AOI22_X1  g041(.A1(new_n198), .A2(new_n204), .B1(new_n208), .B2(new_n209), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT69), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n212), .A2(new_n227), .A3(new_n230), .ZN(new_n231));
  XOR2_X1   g045(.A(G116), .B(G119), .Z(new_n232));
  XNOR2_X1  g046(.A(KEYINPUT2), .B(G113), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(G113), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(KEYINPUT2), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT2), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(G113), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  XNOR2_X1  g053(.A(G116), .B(G119), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT68), .ZN(new_n241));
  AND3_X1   g055(.A1(new_n239), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n241), .B1(new_n239), .B2(new_n240), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n234), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n244), .A2(KEYINPUT70), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT70), .ZN(new_n246));
  OAI21_X1  g060(.A(KEYINPUT68), .B1(new_n232), .B2(new_n233), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n239), .A2(new_n240), .A3(new_n241), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n246), .B1(new_n249), .B2(new_n234), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n245), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(KEYINPUT0), .A2(G128), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n202), .A2(new_n252), .ZN(new_n253));
  XOR2_X1   g067(.A(KEYINPUT0), .B(G128), .Z(new_n254));
  OAI21_X1  g068(.A(new_n253), .B1(new_n202), .B2(new_n254), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n216), .A2(G134), .ZN(new_n256));
  AOI211_X1 g070(.A(G131), .B(new_n256), .C1(new_n214), .C2(new_n217), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n219), .B1(new_n218), .B2(new_n220), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n255), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n231), .A2(new_n251), .A3(new_n259), .ZN(new_n260));
  NOR2_X1   g074(.A1(G237), .A2(G953), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G210), .ZN(new_n262));
  XOR2_X1   g076(.A(new_n262), .B(KEYINPUT27), .Z(new_n263));
  XNOR2_X1  g077(.A(KEYINPUT26), .B(G101), .ZN(new_n264));
  XOR2_X1   g078(.A(new_n263), .B(new_n264), .Z(new_n265));
  INV_X1    g079(.A(KEYINPUT30), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n259), .B(new_n266), .C1(new_n228), .C2(new_n226), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n231), .A2(new_n259), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n268), .B1(new_n269), .B2(KEYINPUT30), .ZN(new_n270));
  INV_X1    g084(.A(new_n244), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n260), .B(new_n265), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT71), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n266), .B1(new_n231), .B2(new_n259), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n244), .B1(new_n275), .B2(new_n268), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n276), .A2(KEYINPUT71), .A3(new_n260), .A4(new_n265), .ZN(new_n277));
  AND3_X1   g091(.A1(new_n274), .A2(KEYINPUT31), .A3(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT31), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n276), .A2(new_n279), .A3(new_n260), .A4(new_n265), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT28), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n259), .B1(new_n228), .B2(new_n226), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT72), .ZN(new_n283));
  AND3_X1   g097(.A1(new_n282), .A2(new_n283), .A3(new_n244), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n283), .B1(new_n282), .B2(new_n244), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n281), .B1(new_n286), .B2(new_n260), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n231), .A2(KEYINPUT73), .A3(new_n259), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(KEYINPUT73), .B1(new_n231), .B2(new_n259), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n251), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n287), .B1(new_n281), .B2(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n280), .B1(new_n292), .B2(new_n265), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n191), .B1(new_n278), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT32), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n282), .A2(new_n244), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(KEYINPUT72), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n282), .A2(new_n283), .A3(new_n244), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n260), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(KEYINPUT28), .ZN(new_n301));
  INV_X1    g115(.A(new_n251), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT73), .ZN(new_n303));
  AND3_X1   g117(.A1(new_n205), .A2(new_n229), .A3(new_n210), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n229), .B1(new_n205), .B2(new_n210), .ZN(new_n305));
  NOR3_X1   g119(.A1(new_n304), .A2(new_n305), .A3(new_n226), .ZN(new_n306));
  INV_X1    g120(.A(new_n259), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n303), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n302), .B1(new_n308), .B2(new_n288), .ZN(new_n309));
  OAI211_X1 g123(.A(new_n301), .B(new_n265), .C1(new_n309), .C2(KEYINPUT28), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(KEYINPUT75), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n291), .A2(new_n281), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT75), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n312), .A2(new_n313), .A3(new_n265), .A4(new_n301), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n265), .B1(new_n276), .B2(new_n260), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n315), .A2(KEYINPUT29), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n311), .A2(new_n314), .A3(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n260), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n251), .B1(new_n231), .B2(new_n259), .ZN(new_n319));
  OAI21_X1  g133(.A(KEYINPUT28), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n320), .B1(new_n309), .B2(KEYINPUT28), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  AND2_X1   g136(.A1(new_n265), .A2(KEYINPUT29), .ZN(new_n323));
  AOI21_X1  g137(.A(G902), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n317), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(G472), .ZN(new_n326));
  INV_X1    g140(.A(new_n265), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n301), .B1(new_n309), .B2(KEYINPUT28), .ZN(new_n328));
  AND3_X1   g142(.A1(new_n276), .A2(new_n260), .A3(new_n265), .ZN(new_n329));
  AOI22_X1  g143(.A1(new_n327), .A2(new_n328), .B1(new_n329), .B2(new_n279), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n274), .A2(KEYINPUT31), .A3(new_n277), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n190), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(KEYINPUT32), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n296), .A2(new_n326), .A3(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT25), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT77), .ZN(new_n336));
  AND2_X1   g150(.A1(KEYINPUT67), .A2(G128), .ZN(new_n337));
  NOR2_X1   g151(.A1(KEYINPUT67), .A2(G128), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n339), .A2(KEYINPUT23), .A3(G119), .ZN(new_n340));
  INV_X1    g154(.A(G119), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(G128), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(KEYINPUT23), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n343), .B1(new_n341), .B2(G128), .ZN(new_n344));
  INV_X1    g158(.A(G110), .ZN(new_n345));
  AND3_X1   g159(.A1(new_n340), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  XOR2_X1   g160(.A(KEYINPUT24), .B(G110), .Z(new_n347));
  NAND2_X1  g161(.A1(new_n339), .A2(G119), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n347), .B1(new_n348), .B2(new_n342), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n336), .B1(new_n346), .B2(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n340), .A2(new_n344), .A3(new_n345), .ZN(new_n351));
  AND2_X1   g165(.A1(new_n348), .A2(new_n342), .ZN(new_n352));
  OAI211_X1 g166(.A(new_n351), .B(KEYINPUT77), .C1(new_n352), .C2(new_n347), .ZN(new_n353));
  XNOR2_X1  g167(.A(G125), .B(G140), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(KEYINPUT16), .ZN(new_n355));
  INV_X1    g169(.A(G140), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(G125), .ZN(new_n357));
  OR2_X1    g171(.A1(new_n357), .A2(KEYINPUT16), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n355), .A2(G146), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n354), .A2(new_n192), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n350), .A2(new_n353), .A3(new_n359), .A4(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n355), .A2(new_n358), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(new_n192), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(new_n359), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n352), .A2(new_n347), .ZN(new_n365));
  AND2_X1   g179(.A1(new_n340), .A2(new_n344), .ZN(new_n366));
  OAI211_X1 g180(.A(new_n364), .B(new_n365), .C1(new_n345), .C2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n361), .A2(new_n367), .ZN(new_n368));
  XNOR2_X1  g182(.A(KEYINPUT22), .B(G137), .ZN(new_n369));
  INV_X1    g183(.A(G221), .ZN(new_n370));
  INV_X1    g184(.A(G234), .ZN(new_n371));
  NOR3_X1   g185(.A1(new_n370), .A2(new_n371), .A3(G953), .ZN(new_n372));
  XOR2_X1   g186(.A(new_n369), .B(new_n372), .Z(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n368), .A2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT78), .ZN(new_n376));
  AND3_X1   g190(.A1(new_n361), .A2(new_n367), .A3(new_n376), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n376), .B1(new_n361), .B2(new_n367), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n375), .B1(new_n379), .B2(new_n374), .ZN(new_n380));
  INV_X1    g194(.A(G902), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n335), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n368), .A2(KEYINPUT78), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n361), .A2(new_n367), .A3(new_n376), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n383), .A2(new_n374), .A3(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n375), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n385), .A2(new_n386), .A3(new_n335), .A4(new_n381), .ZN(new_n387));
  OAI21_X1  g201(.A(G217), .B1(new_n371), .B2(G902), .ZN(new_n388));
  XNOR2_X1  g202(.A(new_n388), .B(KEYINPUT76), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n382), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n388), .A2(new_n381), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  AND2_X1   g207(.A1(new_n380), .A2(new_n393), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n391), .A2(new_n394), .ZN(new_n395));
  AND2_X1   g209(.A1(new_n334), .A2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(G469), .ZN(new_n397));
  XNOR2_X1  g211(.A(G110), .B(G140), .ZN(new_n398));
  INV_X1    g212(.A(G953), .ZN(new_n399));
  AND2_X1   g213(.A1(new_n399), .A2(G227), .ZN(new_n400));
  XOR2_X1   g214(.A(new_n398), .B(new_n400), .Z(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(G107), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(KEYINPUT79), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT79), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(G107), .ZN(new_n406));
  AOI21_X1  g220(.A(G104), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(G104), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n408), .A2(G107), .ZN(new_n409));
  OAI21_X1  g223(.A(G101), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT3), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n411), .B1(new_n403), .B2(G104), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n403), .A2(G104), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n408), .A2(KEYINPUT3), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n415), .A2(new_n404), .A3(new_n406), .ZN(new_n416));
  INV_X1    g230(.A(G101), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n414), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n410), .A2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT80), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n410), .A2(KEYINPUT80), .A3(new_n418), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n423), .A2(new_n212), .A3(KEYINPUT10), .A4(new_n230), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT10), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT1), .ZN(new_n426));
  OAI22_X1  g240(.A1(new_n202), .A2(G128), .B1(new_n426), .B2(new_n195), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n427), .B1(new_n198), .B2(new_n204), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n425), .B1(new_n428), .B2(new_n419), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n417), .B1(new_n414), .B2(new_n416), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT4), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n418), .A2(KEYINPUT4), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n432), .B(new_n255), .C1(new_n433), .C2(new_n430), .ZN(new_n434));
  AND2_X1   g248(.A1(new_n429), .A2(new_n434), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n257), .A2(new_n258), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n424), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT81), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n424), .A2(new_n435), .A3(KEYINPUT81), .A4(new_n436), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n402), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(new_n436), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT82), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n228), .A2(new_n443), .A3(new_n419), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n444), .B1(new_n419), .B2(new_n428), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n443), .B1(new_n228), .B2(new_n419), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n442), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT12), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n448), .B1(new_n436), .B2(KEYINPUT83), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n442), .B(new_n449), .C1(new_n445), .C2(new_n446), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AND2_X1   g267(.A1(new_n441), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n439), .A2(new_n440), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n429), .A2(new_n434), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n304), .A2(new_n305), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n425), .B1(new_n421), .B2(new_n422), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n456), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  OR2_X1    g273(.A1(new_n459), .A2(new_n436), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n401), .B1(new_n455), .B2(new_n460), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n397), .B(new_n381), .C1(new_n454), .C2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n455), .A2(new_n453), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(new_n402), .ZN(new_n464));
  AOI21_X1  g278(.A(KEYINPUT81), .B1(new_n459), .B2(new_n436), .ZN(new_n465));
  INV_X1    g279(.A(new_n440), .ZN(new_n466));
  OAI211_X1 g280(.A(KEYINPUT84), .B(new_n401), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(new_n460), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n441), .A2(KEYINPUT84), .ZN(new_n469));
  OAI211_X1 g283(.A(G469), .B(new_n464), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n397), .A2(new_n381), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n462), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  XNOR2_X1  g287(.A(KEYINPUT9), .B(G234), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n370), .B1(new_n475), .B2(new_n381), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n473), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT94), .ZN(new_n479));
  INV_X1    g293(.A(G122), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(G116), .ZN(new_n481));
  INV_X1    g295(.A(G116), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(G122), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n404), .A2(new_n406), .A3(new_n481), .A4(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n338), .ZN(new_n485));
  NAND2_X1  g299(.A1(KEYINPUT67), .A2(G128), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n485), .A2(G143), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n194), .A2(G128), .ZN(new_n488));
  AND3_X1   g302(.A1(new_n487), .A2(new_n213), .A3(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n213), .B1(new_n487), .B2(new_n488), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n484), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(KEYINPUT14), .B1(new_n480), .B2(G116), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n480), .A2(G116), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT92), .ZN(new_n494));
  NOR3_X1   g308(.A1(new_n492), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n483), .A2(KEYINPUT14), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n494), .B1(new_n492), .B2(new_n493), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n403), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n491), .A2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT91), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n404), .A2(new_n406), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n481), .A2(new_n483), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT90), .ZN(new_n505));
  AND3_X1   g319(.A1(new_n504), .A2(new_n505), .A3(new_n484), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n505), .B1(new_n504), .B2(new_n484), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n487), .A2(KEYINPUT13), .A3(new_n488), .ZN(new_n509));
  INV_X1    g323(.A(new_n488), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT13), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n213), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n510), .B1(new_n339), .B2(G143), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(new_n213), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n501), .B1(new_n508), .B2(new_n516), .ZN(new_n517));
  AND4_X1   g331(.A1(new_n404), .A2(new_n406), .A3(new_n481), .A4(new_n483), .ZN(new_n518));
  AOI22_X1  g332(.A1(new_n404), .A2(new_n406), .B1(new_n481), .B2(new_n483), .ZN(new_n519));
  OAI21_X1  g333(.A(KEYINPUT90), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n504), .A2(new_n505), .A3(new_n484), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI22_X1  g336(.A1(new_n509), .A2(new_n512), .B1(new_n514), .B2(new_n213), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n522), .A2(KEYINPUT91), .A3(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n500), .B1(new_n517), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n475), .A2(G217), .A3(new_n399), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n479), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  OR2_X1    g342(.A1(new_n491), .A2(new_n499), .ZN(new_n529));
  AND3_X1   g343(.A1(new_n522), .A2(KEYINPUT91), .A3(new_n523), .ZN(new_n530));
  AOI21_X1  g344(.A(KEYINPUT91), .B1(new_n522), .B2(new_n523), .ZN(new_n531));
  OAI211_X1 g345(.A(new_n529), .B(new_n527), .C1(new_n530), .C2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(KEYINPUT93), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n534), .A2(KEYINPUT94), .A3(new_n526), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n517), .A2(new_n524), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT93), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n536), .A2(new_n537), .A3(new_n529), .A4(new_n527), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n528), .A2(new_n533), .A3(new_n535), .A4(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(new_n381), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(KEYINPUT96), .ZN(new_n541));
  XOR2_X1   g355(.A(KEYINPUT95), .B(KEYINPUT15), .Z(new_n542));
  INV_X1    g356(.A(G478), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT96), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n539), .A2(new_n546), .A3(new_n381), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n541), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n539), .A2(new_n546), .A3(new_n381), .A4(new_n544), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AND2_X1   g364(.A1(new_n399), .A2(G952), .ZN(new_n551));
  INV_X1    g365(.A(G237), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n551), .B1(new_n371), .B2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  OAI211_X1 g368(.A(G902), .B(G953), .C1(new_n371), .C2(new_n552), .ZN(new_n555));
  XOR2_X1   g369(.A(new_n555), .B(KEYINPUT97), .Z(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  XNOR2_X1  g371(.A(KEYINPUT21), .B(G898), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n554), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(G475), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n552), .A2(new_n399), .A3(G214), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(new_n194), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n261), .A2(G143), .A3(G214), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n565), .A2(KEYINPUT18), .A3(G131), .ZN(new_n566));
  NAND2_X1  g380(.A1(KEYINPUT18), .A2(G131), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n563), .A2(new_n564), .A3(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(G125), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(G140), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n357), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(G146), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(new_n360), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n566), .A2(new_n568), .A3(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT88), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n564), .ZN(new_n577));
  AOI21_X1  g391(.A(G143), .B1(new_n261), .B2(G214), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AOI22_X1  g393(.A1(new_n579), .A2(new_n567), .B1(new_n360), .B2(new_n572), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n580), .A2(KEYINPUT88), .A3(new_n566), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n576), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n565), .A2(G131), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT17), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n563), .A2(new_n219), .A3(new_n564), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n565), .A2(KEYINPUT17), .A3(G131), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n586), .A2(new_n363), .A3(new_n587), .A4(new_n359), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n582), .A2(new_n588), .ZN(new_n589));
  XNOR2_X1  g403(.A(G113), .B(G122), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(new_n408), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(KEYINPUT88), .B1(new_n580), .B2(new_n566), .ZN(new_n594));
  AND4_X1   g408(.A1(KEYINPUT88), .A2(new_n566), .A3(new_n568), .A4(new_n573), .ZN(new_n595));
  OAI211_X1 g409(.A(new_n591), .B(new_n588), .C1(new_n594), .C2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n561), .B1(new_n597), .B2(new_n381), .ZN(new_n598));
  INV_X1    g412(.A(new_n596), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n354), .B(KEYINPUT19), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n192), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n583), .A2(new_n585), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n601), .A2(new_n359), .A3(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n591), .B1(new_n582), .B2(new_n603), .ZN(new_n604));
  OAI21_X1  g418(.A(KEYINPUT89), .B1(new_n599), .B2(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(G475), .A2(G902), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT89), .ZN(new_n607));
  INV_X1    g421(.A(new_n359), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n608), .B1(new_n192), .B2(new_n600), .ZN(new_n609));
  AOI22_X1  g423(.A1(new_n576), .A2(new_n581), .B1(new_n609), .B2(new_n602), .ZN(new_n610));
  OAI211_X1 g424(.A(new_n596), .B(new_n607), .C1(new_n610), .C2(new_n591), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n605), .A2(new_n606), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(KEYINPUT20), .ZN(new_n613));
  NOR3_X1   g427(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n614), .B1(new_n599), .B2(new_n604), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n598), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n550), .A2(new_n560), .A3(new_n616), .ZN(new_n617));
  OAI21_X1  g431(.A(G210), .B1(G237), .B2(G902), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(KEYINPUT87), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n255), .A2(G125), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n622), .B1(new_n228), .B2(G125), .ZN(new_n623));
  INV_X1    g437(.A(G224), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n624), .A2(G953), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n623), .B(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(G110), .B(G122), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT85), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n240), .A2(KEYINPUT5), .ZN(new_n629));
  NOR3_X1   g443(.A1(new_n482), .A2(KEYINPUT5), .A3(G119), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n630), .A2(new_n235), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n249), .A2(new_n632), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n633), .B1(new_n421), .B2(new_n422), .ZN(new_n634));
  AND3_X1   g448(.A1(new_n415), .A2(new_n404), .A3(new_n406), .ZN(new_n635));
  AOI21_X1  g449(.A(KEYINPUT3), .B1(new_n408), .B2(G107), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n636), .A2(new_n409), .ZN(new_n637));
  OAI21_X1  g451(.A(G101), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n638), .A2(KEYINPUT4), .A3(new_n418), .ZN(new_n639));
  AND3_X1   g453(.A1(new_n639), .A2(new_n244), .A3(new_n432), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n628), .B1(new_n634), .B2(new_n640), .ZN(new_n641));
  AOI22_X1  g455(.A1(new_n247), .A2(new_n248), .B1(new_n631), .B2(new_n629), .ZN(new_n642));
  AND3_X1   g456(.A1(new_n410), .A2(KEYINPUT80), .A3(new_n418), .ZN(new_n643));
  AOI21_X1  g457(.A(KEYINPUT80), .B1(new_n410), .B2(new_n418), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n642), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n639), .A2(new_n244), .A3(new_n432), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n645), .A2(KEYINPUT85), .A3(new_n646), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n627), .B1(new_n641), .B2(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n645), .A2(new_n646), .A3(new_n627), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  OAI21_X1  g464(.A(KEYINPUT6), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n627), .ZN(new_n652));
  AND3_X1   g466(.A1(new_n645), .A2(KEYINPUT85), .A3(new_n646), .ZN(new_n653));
  AOI21_X1  g467(.A(KEYINPUT85), .B1(new_n645), .B2(new_n646), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n652), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT6), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n626), .B1(new_n651), .B2(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n627), .B(KEYINPUT8), .ZN(new_n659));
  OR2_X1    g473(.A1(new_n629), .A2(KEYINPUT86), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n629), .A2(KEYINPUT86), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n660), .A2(new_n631), .A3(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n419), .ZN(new_n663));
  AND3_X1   g477(.A1(new_n662), .A2(new_n663), .A3(new_n249), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n663), .A2(new_n642), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n659), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n625), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n623), .A2(KEYINPUT7), .A3(new_n667), .ZN(new_n668));
  AND2_X1   g482(.A1(new_n667), .A2(KEYINPUT7), .ZN(new_n669));
  OR2_X1    g483(.A1(new_n623), .A2(new_n669), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n666), .A2(new_n649), .A3(new_n668), .A4(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(new_n381), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n621), .B1(new_n658), .B2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n626), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n656), .B1(new_n655), .B2(new_n649), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n641), .A2(new_n647), .ZN(new_n676));
  AOI21_X1  g490(.A(KEYINPUT6), .B1(new_n676), .B2(new_n652), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n674), .B1(new_n675), .B2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n672), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n678), .A2(new_n679), .A3(new_n620), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n673), .A2(new_n680), .ZN(new_n681));
  OAI21_X1  g495(.A(G214), .B1(G237), .B2(G902), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NOR3_X1   g497(.A1(new_n478), .A2(new_n617), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n396), .A2(new_n684), .ZN(new_n685));
  XOR2_X1   g499(.A(KEYINPUT98), .B(G101), .Z(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(G3));
  AOI21_X1  g501(.A(G902), .B1(new_n330), .B2(new_n331), .ZN(new_n688));
  INV_X1    g502(.A(G472), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n294), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT99), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n460), .B1(new_n465), .B2(new_n466), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n402), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n441), .A2(new_n453), .ZN(new_n695));
  AOI21_X1  g509(.A(G902), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n471), .B1(new_n696), .B2(new_n397), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n476), .B1(new_n697), .B2(new_n470), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n691), .A2(new_n692), .A3(new_n395), .A4(new_n698), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n473), .A2(new_n395), .A3(new_n477), .ZN(new_n700));
  OAI21_X1  g514(.A(KEYINPUT99), .B1(new_n700), .B2(new_n690), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(new_n682), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n619), .B1(new_n658), .B2(new_n672), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n678), .A2(new_n679), .A3(new_n618), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n704), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n560), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n613), .A2(new_n615), .ZN(new_n709));
  INV_X1    g523(.A(new_n598), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n543), .A2(G902), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n539), .A2(KEYINPUT33), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT100), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n534), .A2(new_n716), .A3(new_n526), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n716), .B1(new_n534), .B2(new_n526), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n532), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(KEYINPUT33), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n713), .B1(new_n715), .B2(new_n721), .ZN(new_n722));
  XOR2_X1   g536(.A(KEYINPUT101), .B(G478), .Z(new_n723));
  NAND2_X1  g537(.A1(new_n540), .A2(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(new_n724), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n711), .B1(new_n722), .B2(new_n725), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n708), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n703), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(KEYINPUT102), .ZN(new_n729));
  XNOR2_X1  g543(.A(KEYINPUT34), .B(G104), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n729), .B(new_n730), .ZN(G6));
  NAND3_X1  g545(.A1(new_n605), .A2(new_n611), .A3(new_n614), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n598), .B1(new_n613), .B2(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  NOR3_X1   g548(.A1(new_n708), .A2(new_n550), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n703), .A2(new_n735), .ZN(new_n736));
  XOR2_X1   g550(.A(KEYINPUT35), .B(G107), .Z(new_n737));
  XNOR2_X1  g551(.A(new_n736), .B(new_n737), .ZN(G9));
  OAI21_X1  g552(.A(new_n379), .B1(KEYINPUT36), .B2(new_n374), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n374), .A2(KEYINPUT36), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n740), .B1(new_n377), .B2(new_n378), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n739), .A2(new_n741), .A3(new_n393), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n742), .B1(new_n382), .B2(new_n390), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n684), .A2(new_n691), .A3(new_n743), .ZN(new_n744));
  XOR2_X1   g558(.A(KEYINPUT37), .B(G110), .Z(new_n745));
  XNOR2_X1  g559(.A(new_n744), .B(new_n745), .ZN(G12));
  NOR3_X1   g560(.A1(new_n658), .A2(new_n672), .A3(new_n619), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n618), .B1(new_n678), .B2(new_n679), .ZN(new_n748));
  OAI211_X1 g562(.A(new_n743), .B(new_n682), .C1(new_n747), .C2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(G900), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n554), .B1(new_n557), .B2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(KEYINPUT103), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n548), .A2(new_n549), .A3(new_n733), .A4(new_n753), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n749), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n334), .A2(new_n698), .A3(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G128), .ZN(G30));
  XOR2_X1   g571(.A(new_n681), .B(KEYINPUT38), .Z(new_n758));
  NAND3_X1  g572(.A1(new_n548), .A2(new_n711), .A3(new_n549), .ZN(new_n759));
  NOR4_X1   g573(.A1(new_n758), .A2(new_n704), .A3(new_n743), .A4(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n752), .B(KEYINPUT39), .ZN(new_n761));
  OAI21_X1  g575(.A(KEYINPUT40), .B1(new_n478), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n327), .B1(new_n318), .B2(new_n319), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n274), .A2(new_n277), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(KEYINPUT104), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(new_n381), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n764), .A2(KEYINPUT104), .ZN(new_n767));
  OAI21_X1  g581(.A(G472), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n768), .A2(new_n296), .A3(new_n333), .ZN(new_n769));
  OR3_X1    g583(.A1(new_n478), .A2(KEYINPUT40), .A3(new_n761), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n760), .A2(new_n762), .A3(new_n769), .A4(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G143), .ZN(G45));
  OAI211_X1 g586(.A(new_n711), .B(new_n753), .C1(new_n722), .C2(new_n725), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n773), .A2(new_n749), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n334), .A2(new_n774), .A3(new_n698), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G146), .ZN(G48));
  AOI22_X1  g590(.A1(new_n693), .A2(new_n402), .B1(new_n441), .B2(new_n453), .ZN(new_n777));
  OAI21_X1  g591(.A(G469), .B1(new_n777), .B2(G902), .ZN(new_n778));
  AND3_X1   g592(.A1(new_n778), .A2(new_n477), .A3(new_n462), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n727), .A2(new_n334), .A3(new_n395), .A4(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(KEYINPUT41), .B(G113), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n780), .B(new_n781), .ZN(G15));
  NAND4_X1  g596(.A1(new_n735), .A2(new_n334), .A3(new_n395), .A4(new_n779), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G116), .ZN(G18));
  INV_X1    g598(.A(new_n743), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n617), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n778), .A2(new_n462), .A3(new_n477), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n682), .B1(new_n747), .B2(new_n748), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n786), .A2(new_n334), .A3(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G119), .ZN(G21));
  INV_X1    g605(.A(KEYINPUT107), .ZN(new_n792));
  AND3_X1   g606(.A1(new_n548), .A2(new_n711), .A3(new_n549), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n779), .A2(new_n560), .A3(new_n707), .A4(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n190), .B(KEYINPUT105), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n331), .A2(new_n280), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT106), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n321), .A2(new_n798), .ZN(new_n799));
  OAI211_X1 g613(.A(new_n320), .B(KEYINPUT106), .C1(new_n309), .C2(KEYINPUT28), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n265), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n796), .B1(new_n797), .B2(new_n801), .ZN(new_n802));
  OAI211_X1 g616(.A(new_n802), .B(new_n395), .C1(new_n689), .C2(new_n688), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n792), .B1(new_n794), .B2(new_n803), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n778), .A2(new_n462), .A3(new_n477), .A4(new_n560), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n805), .A2(new_n788), .A3(new_n759), .ZN(new_n806));
  AOI21_X1  g620(.A(KEYINPUT106), .B1(new_n312), .B2(new_n320), .ZN(new_n807));
  INV_X1    g621(.A(new_n800), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n327), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n809), .A2(new_n331), .A3(new_n280), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n381), .B1(new_n278), .B2(new_n293), .ZN(new_n811));
  AOI22_X1  g625(.A1(new_n810), .A2(new_n796), .B1(new_n811), .B2(G472), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n806), .A2(KEYINPUT107), .A3(new_n812), .A4(new_n395), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n804), .A2(new_n813), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(G122), .ZN(G24));
  INV_X1    g629(.A(KEYINPUT33), .ZN(new_n816));
  INV_X1    g630(.A(new_n719), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(new_n717), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n816), .B1(new_n818), .B2(new_n532), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n712), .B1(new_n819), .B2(new_n714), .ZN(new_n820));
  AOI211_X1 g634(.A(new_n752), .B(new_n616), .C1(new_n820), .C2(new_n724), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n812), .A2(new_n789), .A3(new_n743), .A4(new_n821), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n822), .B(G125), .ZN(G27));
  OAI21_X1  g637(.A(KEYINPUT108), .B1(new_n468), .B2(new_n469), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n401), .B1(new_n465), .B2(new_n466), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT84), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT108), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n827), .A2(new_n828), .A3(new_n460), .A4(new_n467), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n824), .A2(new_n829), .A3(G469), .A4(new_n464), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(new_n697), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n673), .A2(new_n477), .A3(new_n680), .A4(new_n682), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n831), .A2(new_n821), .A3(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT109), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n835), .B1(new_n332), .B2(KEYINPUT32), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n294), .A2(KEYINPUT109), .A3(new_n295), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n836), .A2(new_n837), .A3(new_n333), .A4(new_n326), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n834), .A2(new_n838), .A3(new_n395), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(KEYINPUT42), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n773), .A2(KEYINPUT42), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n832), .B1(new_n697), .B2(new_n830), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n334), .A2(new_n841), .A3(new_n395), .A4(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n844), .B(new_n219), .ZN(G33));
  XOR2_X1   g659(.A(new_n754), .B(KEYINPUT110), .Z(new_n846));
  NAND4_X1  g660(.A1(new_n846), .A2(new_n334), .A3(new_n395), .A4(new_n842), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(G134), .ZN(G36));
  NAND3_X1  g662(.A1(new_n673), .A2(new_n682), .A3(new_n680), .ZN(new_n849));
  INV_X1    g663(.A(new_n849), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n711), .B1(new_n820), .B2(new_n724), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n851), .B(KEYINPUT43), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n852), .A2(new_n690), .A3(new_n743), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT44), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n850), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT113), .ZN(new_n856));
  OR2_X1    g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n855), .A2(new_n856), .ZN(new_n858));
  AOI22_X1  g672(.A1(new_n857), .A2(new_n858), .B1(new_n854), .B2(new_n853), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n464), .B1(new_n468), .B2(new_n469), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT45), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n397), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n824), .A2(new_n829), .A3(KEYINPUT45), .A4(new_n464), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n471), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AOI22_X1  g678(.A1(new_n864), .A2(KEYINPUT46), .B1(new_n397), .B2(new_n696), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(KEYINPUT111), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n866), .B1(KEYINPUT46), .B2(new_n864), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n865), .A2(KEYINPUT111), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n477), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n869), .A2(new_n761), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT112), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n869), .A2(KEYINPUT112), .A3(new_n761), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n859), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n874), .B(G137), .ZN(G39));
  INV_X1    g689(.A(KEYINPUT47), .ZN(new_n876));
  OR2_X1    g690(.A1(new_n869), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n869), .A2(new_n876), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NOR4_X1   g693(.A1(new_n334), .A2(new_n395), .A3(new_n773), .A4(new_n849), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(G140), .ZN(G42));
  NAND2_X1  g696(.A1(new_n852), .A2(new_n554), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n778), .A2(new_n462), .ZN(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(new_n833), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n838), .A2(new_n395), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n889), .B(KEYINPUT48), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n883), .A2(new_n803), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(new_n789), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n395), .A2(new_n554), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n769), .A2(new_n886), .A3(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(new_n726), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n890), .A2(new_n551), .A3(new_n892), .A4(new_n896), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n812), .A2(new_n743), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n722), .A2(new_n711), .A3(new_n725), .ZN(new_n899));
  AOI22_X1  g713(.A1(new_n887), .A2(new_n898), .B1(new_n894), .B2(new_n899), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n758), .A2(new_n704), .A3(new_n779), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT119), .ZN(new_n902));
  AND3_X1   g716(.A1(new_n902), .A2(KEYINPUT50), .A3(new_n891), .ZN(new_n903));
  AOI21_X1  g717(.A(KEYINPUT50), .B1(new_n902), .B2(new_n891), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n900), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n885), .A2(new_n476), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n877), .A2(new_n878), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n891), .A2(new_n850), .ZN(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n905), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n897), .B1(new_n910), .B2(KEYINPUT51), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n911), .B1(KEYINPUT51), .B2(new_n910), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT52), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT115), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n752), .A2(new_n476), .ZN(new_n915));
  OAI211_X1 g729(.A(new_n742), .B(new_n915), .C1(new_n382), .C2(new_n390), .ZN(new_n916));
  INV_X1    g730(.A(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n914), .B1(new_n831), .B2(new_n917), .ZN(new_n918));
  AOI211_X1 g732(.A(KEYINPUT115), .B(new_n916), .C1(new_n830), .C2(new_n697), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n788), .A2(new_n759), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n769), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n756), .A2(new_n775), .A3(new_n822), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n913), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT116), .ZN(new_n926));
  INV_X1    g740(.A(new_n918), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n831), .A2(new_n914), .A3(new_n917), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n769), .A2(new_n921), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n913), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  AND3_X1   g745(.A1(new_n775), .A2(new_n756), .A3(new_n822), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n926), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g747(.A(KEYINPUT52), .B1(new_n920), .B2(new_n922), .ZN(new_n934));
  NOR3_X1   g748(.A1(new_n934), .A2(new_n924), .A3(KEYINPUT116), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n925), .B1(new_n933), .B2(new_n935), .ZN(new_n936));
  AOI211_X1 g750(.A(new_n598), .B(new_n752), .C1(new_n613), .C2(new_n732), .ZN(new_n937));
  AND3_X1   g751(.A1(new_n539), .A2(new_n546), .A3(new_n381), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n546), .B1(new_n539), .B2(new_n381), .ZN(new_n939));
  NOR3_X1   g753(.A1(new_n938), .A2(new_n939), .A3(new_n544), .ZN(new_n940));
  INV_X1    g754(.A(new_n549), .ZN(new_n941));
  OAI211_X1 g755(.A(new_n743), .B(new_n937), .C1(new_n940), .C2(new_n941), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n942), .A2(new_n849), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n334), .A2(new_n698), .A3(new_n943), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n812), .A2(new_n842), .A3(new_n743), .A4(new_n821), .ZN(new_n945));
  AND2_X1   g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n840), .A2(new_n946), .A3(new_n843), .A4(new_n847), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT53), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n726), .B1(new_n550), .B2(new_n711), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n683), .A2(new_n559), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n699), .A2(new_n701), .A3(new_n949), .A4(new_n950), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n951), .A2(new_n685), .A3(new_n744), .ZN(new_n952));
  NOR3_X1   g766(.A1(new_n947), .A2(new_n948), .A3(new_n952), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n814), .A2(new_n780), .A3(new_n783), .A4(new_n790), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(KEYINPUT118), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n780), .A2(new_n790), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT118), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n956), .A2(new_n957), .A3(new_n783), .A4(new_n814), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n936), .A2(new_n953), .A3(new_n955), .A4(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT54), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n931), .A2(new_n932), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n925), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n954), .A2(new_n952), .ZN(new_n963));
  AND4_X1   g777(.A1(new_n840), .A2(new_n946), .A3(new_n843), .A4(new_n847), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n962), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(new_n948), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n959), .A2(new_n960), .A3(new_n966), .ZN(new_n967));
  NOR3_X1   g781(.A1(new_n947), .A2(new_n954), .A3(new_n952), .ZN(new_n968));
  AOI21_X1  g782(.A(KEYINPUT53), .B1(new_n936), .B2(new_n968), .ZN(new_n969));
  OR3_X1    g783(.A1(new_n965), .A2(KEYINPUT117), .A3(new_n948), .ZN(new_n970));
  OAI21_X1  g784(.A(KEYINPUT117), .B1(new_n965), .B2(new_n948), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n969), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n967), .B1(new_n972), .B2(new_n960), .ZN(new_n973));
  OAI22_X1  g787(.A1(new_n912), .A2(new_n973), .B1(G952), .B2(G953), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n395), .A2(new_n477), .A3(new_n682), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n975), .B(KEYINPUT114), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n884), .B(KEYINPUT49), .Z(new_n977));
  NAND4_X1  g791(.A1(new_n976), .A2(new_n758), .A3(new_n851), .A4(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n974), .B1(new_n769), .B2(new_n978), .ZN(G75));
  NOR2_X1   g793(.A1(new_n675), .A2(new_n677), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n980), .B(new_n674), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n981), .B(KEYINPUT55), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n381), .B1(new_n959), .B2(new_n966), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n983), .A2(G210), .ZN(new_n984));
  INV_X1    g798(.A(KEYINPUT56), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n985), .A2(KEYINPUT120), .ZN(new_n986));
  OR2_X1    g800(.A1(new_n985), .A2(KEYINPUT120), .ZN(new_n987));
  AND4_X1   g801(.A1(new_n982), .A2(new_n984), .A3(new_n986), .A4(new_n987), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n982), .B1(new_n984), .B2(new_n985), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n399), .A2(G952), .ZN(new_n990));
  NOR3_X1   g804(.A1(new_n988), .A2(new_n989), .A3(new_n990), .ZN(G51));
  NAND3_X1  g805(.A1(new_n983), .A2(new_n863), .A3(new_n862), .ZN(new_n992));
  XOR2_X1   g806(.A(new_n992), .B(KEYINPUT121), .Z(new_n993));
  NAND2_X1  g807(.A1(new_n959), .A2(new_n966), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n994), .B(new_n960), .ZN(new_n995));
  XOR2_X1   g809(.A(new_n471), .B(KEYINPUT57), .Z(new_n996));
  OAI22_X1  g810(.A1(new_n995), .A2(new_n996), .B1(new_n461), .B2(new_n454), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n990), .B1(new_n993), .B2(new_n997), .ZN(G54));
  NAND3_X1  g812(.A1(new_n983), .A2(KEYINPUT58), .A3(G475), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n605), .A2(new_n611), .ZN(new_n1000));
  AND2_X1   g814(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n999), .A2(new_n1000), .ZN(new_n1002));
  NOR3_X1   g816(.A1(new_n1001), .A2(new_n1002), .A3(new_n990), .ZN(G60));
  NAND2_X1  g817(.A1(new_n715), .A2(new_n721), .ZN(new_n1004));
  XNOR2_X1  g818(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n1005));
  NAND2_X1  g819(.A1(G478), .A2(G902), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n1005), .B(new_n1006), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1004), .B1(new_n973), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g822(.A(new_n990), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1004), .A2(new_n1007), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n1009), .B1(new_n995), .B2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n1008), .A2(new_n1011), .ZN(G63));
  INV_X1    g826(.A(KEYINPUT61), .ZN(new_n1013));
  AND2_X1   g827(.A1(new_n739), .A2(new_n741), .ZN(new_n1014));
  NAND2_X1  g828(.A1(G217), .A2(G902), .ZN(new_n1015));
  XOR2_X1   g829(.A(new_n1015), .B(KEYINPUT60), .Z(new_n1016));
  AND4_X1   g830(.A1(KEYINPUT53), .A2(new_n951), .A3(new_n685), .A4(new_n744), .ZN(new_n1017));
  NAND4_X1  g831(.A1(new_n955), .A2(new_n964), .A3(new_n1017), .A4(new_n958), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n929), .A2(new_n930), .ZN(new_n1019));
  AOI21_X1  g833(.A(KEYINPUT52), .B1(new_n932), .B2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g834(.A(KEYINPUT116), .B1(new_n934), .B2(new_n924), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n931), .A2(new_n932), .A3(new_n926), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n1020), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g837(.A1(new_n1018), .A2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g838(.A(KEYINPUT53), .B1(new_n968), .B2(new_n962), .ZN(new_n1025));
  OAI211_X1 g839(.A(new_n1014), .B(new_n1016), .C1(new_n1024), .C2(new_n1025), .ZN(new_n1026));
  INV_X1    g840(.A(new_n1016), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n1027), .B1(new_n959), .B2(new_n966), .ZN(new_n1028));
  OAI211_X1 g842(.A(new_n1026), .B(new_n1009), .C1(new_n1028), .C2(new_n380), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n1013), .B1(new_n1029), .B2(KEYINPUT124), .ZN(new_n1030));
  AOI21_X1  g844(.A(KEYINPUT124), .B1(new_n1029), .B2(KEYINPUT123), .ZN(new_n1031));
  XNOR2_X1  g845(.A(new_n1030), .B(new_n1031), .ZN(G66));
  NOR3_X1   g846(.A1(new_n558), .A2(new_n624), .A3(new_n399), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n1033), .B1(new_n963), .B2(new_n399), .ZN(new_n1034));
  OAI21_X1  g848(.A(new_n980), .B1(G898), .B2(new_n399), .ZN(new_n1035));
  XNOR2_X1  g849(.A(new_n1034), .B(new_n1035), .ZN(G69));
  AOI21_X1  g850(.A(new_n399), .B1(G227), .B2(G900), .ZN(new_n1037));
  NAND4_X1  g851(.A1(new_n932), .A2(new_n840), .A3(new_n843), .A4(new_n847), .ZN(new_n1038));
  AOI21_X1  g852(.A(new_n1038), .B1(new_n879), .B2(new_n880), .ZN(new_n1039));
  OAI211_X1 g853(.A(new_n921), .B(new_n888), .C1(new_n872), .C2(new_n873), .ZN(new_n1040));
  NAND4_X1  g854(.A1(new_n1039), .A2(new_n1040), .A3(new_n874), .A4(new_n399), .ZN(new_n1041));
  XOR2_X1   g855(.A(new_n600), .B(KEYINPUT125), .Z(new_n1042));
  XNOR2_X1  g856(.A(new_n270), .B(new_n1042), .ZN(new_n1043));
  AOI21_X1  g857(.A(new_n1043), .B1(G900), .B2(G953), .ZN(new_n1044));
  NAND2_X1  g858(.A1(new_n1041), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g859(.A(new_n1045), .ZN(new_n1046));
  INV_X1    g860(.A(new_n1043), .ZN(new_n1047));
  NAND2_X1  g861(.A1(new_n771), .A2(new_n932), .ZN(new_n1048));
  XNOR2_X1  g862(.A(new_n1048), .B(KEYINPUT62), .ZN(new_n1049));
  NAND2_X1  g863(.A1(new_n949), .A2(new_n850), .ZN(new_n1050));
  NOR3_X1   g864(.A1(new_n1050), .A2(new_n478), .A3(new_n761), .ZN(new_n1051));
  AOI21_X1  g865(.A(new_n1049), .B1(new_n396), .B2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g866(.A1(new_n1052), .A2(new_n874), .A3(new_n881), .ZN(new_n1053));
  AOI21_X1  g867(.A(new_n1047), .B1(new_n1053), .B2(new_n399), .ZN(new_n1054));
  OAI21_X1  g868(.A(new_n1037), .B1(new_n1046), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g869(.A(new_n1037), .ZN(new_n1056));
  AND2_X1   g870(.A1(new_n1053), .A2(new_n399), .ZN(new_n1057));
  OAI211_X1 g871(.A(new_n1056), .B(new_n1045), .C1(new_n1057), .C2(new_n1047), .ZN(new_n1058));
  NAND2_X1  g872(.A1(new_n1055), .A2(new_n1058), .ZN(G72));
  NAND2_X1  g873(.A1(new_n276), .A2(new_n260), .ZN(new_n1060));
  NAND2_X1  g874(.A1(new_n1060), .A2(new_n265), .ZN(new_n1061));
  NAND4_X1  g875(.A1(new_n1052), .A2(new_n874), .A3(new_n881), .A4(new_n963), .ZN(new_n1062));
  XNOR2_X1  g876(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1063));
  NAND2_X1  g877(.A1(G472), .A2(G902), .ZN(new_n1064));
  XNOR2_X1  g878(.A(new_n1063), .B(new_n1064), .ZN(new_n1065));
  AOI21_X1  g879(.A(new_n1061), .B1(new_n1062), .B2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g880(.A1(new_n1060), .A2(new_n265), .ZN(new_n1067));
  XNOR2_X1  g881(.A(new_n1067), .B(KEYINPUT127), .ZN(new_n1068));
  NAND4_X1  g882(.A1(new_n1039), .A2(new_n1040), .A3(new_n874), .A4(new_n963), .ZN(new_n1069));
  AOI21_X1  g883(.A(new_n1068), .B1(new_n1069), .B2(new_n1065), .ZN(new_n1070));
  NAND2_X1  g884(.A1(new_n274), .A2(new_n277), .ZN(new_n1071));
  OAI21_X1  g885(.A(new_n1065), .B1(new_n1071), .B2(new_n315), .ZN(new_n1072));
  OAI21_X1  g886(.A(new_n1009), .B1(new_n972), .B2(new_n1072), .ZN(new_n1073));
  NOR3_X1   g887(.A1(new_n1066), .A2(new_n1070), .A3(new_n1073), .ZN(G57));
endmodule


