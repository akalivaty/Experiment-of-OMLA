//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 1 1 1 1 0 0 0 1 1 1 0 1 0 0 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 0 1 0 0 0 1 1 1 0 0 0 1 1 1 0 0 0 1 1 0 1 0 0 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:27 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n509, new_n510, new_n511,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n549, new_n550, new_n551,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n565, new_n566, new_n567, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n600, new_n601, new_n602,
    new_n603, new_n606, new_n608, new_n609, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n846, new_n847, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1242, new_n1243, new_n1244,
    new_n1245;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  OAI21_X1  g038(.A(G125), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n461), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  OAI211_X1 g041(.A(G137), .B(new_n461), .C1(new_n462), .C2(new_n463), .ZN(new_n467));
  AND2_X1   g042(.A1(new_n461), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G101), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n466), .A2(new_n470), .ZN(G160));
  OR2_X1    g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(G2105), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G136), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n461), .B1(new_n472), .B2(new_n473), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n461), .A2(G112), .ZN(new_n478));
  OAI21_X1  g053(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n475), .B(new_n477), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  XNOR2_X1  g055(.A(new_n480), .B(KEYINPUT65), .ZN(G162));
  OAI211_X1 g056(.A(G126), .B(G2105), .C1(new_n462), .C2(new_n463), .ZN(new_n482));
  INV_X1    g057(.A(G114), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(G138), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n487), .A2(G2105), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n488), .B1(new_n462), .B2(new_n463), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(KEYINPUT4), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n488), .B(new_n491), .C1(new_n463), .C2(new_n462), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n486), .B1(new_n490), .B2(new_n492), .ZN(G164));
  INV_X1    g068(.A(KEYINPUT5), .ZN(new_n494));
  INV_X1    g069(.A(G543), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(KEYINPUT5), .A2(G543), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AOI22_X1  g073(.A1(new_n498), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n499));
  INV_X1    g074(.A(G651), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  XNOR2_X1  g076(.A(KEYINPUT6), .B(G651), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(G88), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(G543), .ZN(new_n505));
  INV_X1    g080(.A(G50), .ZN(new_n506));
  OAI22_X1  g081(.A1(new_n503), .A2(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n501), .A2(new_n507), .ZN(G166));
  AND2_X1   g083(.A1(new_n496), .A2(new_n497), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n502), .A2(G89), .ZN(new_n510));
  NAND2_X1  g085(.A1(G63), .A2(G651), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g087(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n513));
  XNOR2_X1  g088(.A(new_n513), .B(KEYINPUT7), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n502), .A2(G51), .A3(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n512), .A2(new_n516), .ZN(G168));
  NAND2_X1  g092(.A1(G77), .A2(G543), .ZN(new_n518));
  INV_X1    g093(.A(G64), .ZN(new_n519));
  OAI211_X1 g094(.A(KEYINPUT66), .B(new_n518), .C1(new_n509), .C2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT66), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n519), .B1(new_n496), .B2(new_n497), .ZN(new_n522));
  INV_X1    g097(.A(new_n518), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n520), .A2(G651), .A3(new_n524), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n498), .A2(new_n502), .ZN(new_n526));
  AND2_X1   g101(.A1(KEYINPUT6), .A2(G651), .ZN(new_n527));
  NOR2_X1   g102(.A1(KEYINPUT6), .A2(G651), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n529), .A2(new_n495), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n526), .A2(G90), .B1(new_n530), .B2(G52), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n525), .A2(new_n531), .ZN(G301));
  INV_X1    g107(.A(G301), .ZN(G171));
  AOI22_X1  g108(.A1(new_n526), .A2(G81), .B1(new_n530), .B2(G43), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n498), .A2(G56), .ZN(new_n535));
  NAND2_X1  g110(.A1(G68), .A2(G543), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G651), .ZN(new_n538));
  AOI21_X1  g113(.A(KEYINPUT67), .B1(new_n534), .B2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(G81), .ZN(new_n540));
  INV_X1    g115(.A(G43), .ZN(new_n541));
  OAI22_X1  g116(.A1(new_n503), .A2(new_n540), .B1(new_n505), .B2(new_n541), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n500), .B1(new_n535), .B2(new_n536), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT67), .ZN(new_n544));
  NOR3_X1   g119(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n539), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  NAND4_X1  g122(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g123(.A1(G1), .A2(G3), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT68), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND4_X1  g126(.A1(G319), .A2(G483), .A3(G661), .A4(new_n551), .ZN(G188));
  OAI211_X1 g127(.A(G53), .B(G543), .C1(new_n527), .C2(new_n528), .ZN(new_n553));
  NOR2_X1   g128(.A1(KEYINPUT69), .A2(KEYINPUT9), .ZN(new_n554));
  NAND2_X1  g129(.A1(KEYINPUT69), .A2(KEYINPUT9), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n553), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  NAND4_X1  g132(.A1(new_n502), .A2(G53), .A3(G543), .A4(new_n555), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n526), .A2(G91), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n498), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n561));
  OAI211_X1 g136(.A(new_n559), .B(new_n560), .C1(new_n500), .C2(new_n561), .ZN(G299));
  OR2_X1    g137(.A1(new_n512), .A2(new_n516), .ZN(G286));
  OR2_X1    g138(.A1(new_n501), .A2(new_n507), .ZN(G303));
  OAI21_X1  g139(.A(G651), .B1(new_n498), .B2(G74), .ZN(new_n565));
  INV_X1    g140(.A(G49), .ZN(new_n566));
  INV_X1    g141(.A(G87), .ZN(new_n567));
  OAI221_X1 g142(.A(new_n565), .B1(new_n505), .B2(new_n566), .C1(new_n567), .C2(new_n503), .ZN(G288));
  NAND3_X1  g143(.A1(new_n502), .A2(G48), .A3(G543), .ZN(new_n569));
  INV_X1    g144(.A(G86), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n503), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n498), .A2(G61), .ZN(new_n572));
  NAND2_X1  g147(.A1(G73), .A2(G543), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n500), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(G305));
  AOI22_X1  g151(.A1(new_n498), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n577), .A2(new_n500), .ZN(new_n578));
  INV_X1    g153(.A(G85), .ZN(new_n579));
  INV_X1    g154(.A(G47), .ZN(new_n580));
  OAI22_X1  g155(.A1(new_n503), .A2(new_n579), .B1(new_n505), .B2(new_n580), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(G290));
  NAND2_X1  g158(.A1(G301), .A2(G868), .ZN(new_n584));
  INV_X1    g159(.A(G54), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n585), .B1(new_n505), .B2(KEYINPUT70), .ZN(new_n586));
  OR3_X1    g161(.A1(new_n529), .A2(KEYINPUT70), .A3(new_n495), .ZN(new_n587));
  NAND2_X1  g162(.A1(G79), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G66), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n509), .B2(new_n589), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n586), .A2(new_n587), .B1(new_n590), .B2(G651), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n526), .A2(KEYINPUT10), .A3(G92), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT10), .ZN(new_n593));
  INV_X1    g168(.A(G92), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n503), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  AND2_X1   g171(.A1(new_n591), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n584), .B1(new_n597), .B2(G868), .ZN(G284));
  OAI21_X1  g173(.A(new_n584), .B1(new_n597), .B2(G868), .ZN(G321));
  INV_X1    g174(.A(KEYINPUT71), .ZN(new_n600));
  INV_X1    g175(.A(G868), .ZN(new_n601));
  NOR2_X1   g176(.A1(G168), .A2(new_n601), .ZN(new_n602));
  AOI211_X1 g177(.A(new_n600), .B(new_n602), .C1(new_n601), .C2(G299), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n603), .B1(new_n600), .B2(new_n602), .ZN(G280));
  XNOR2_X1  g179(.A(G280), .B(KEYINPUT72), .ZN(G297));
  INV_X1    g180(.A(G559), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n597), .B1(new_n606), .B2(G860), .ZN(G148));
  NAND2_X1  g182(.A1(new_n597), .A2(new_n606), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(G868), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(G868), .B2(new_n546), .ZN(G323));
  XNOR2_X1  g185(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XNOR2_X1  g186(.A(KEYINPUT3), .B(G2104), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(new_n468), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT12), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT13), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(G2100), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n474), .A2(G135), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n476), .A2(G123), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n461), .A2(G111), .ZN(new_n619));
  OAI21_X1  g194(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n620));
  OAI211_X1 g195(.A(new_n617), .B(new_n618), .C1(new_n619), .C2(new_n620), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT73), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(G2096), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n616), .A2(new_n623), .ZN(G156));
  INV_X1    g199(.A(G14), .ZN(new_n625));
  XOR2_X1   g200(.A(KEYINPUT15), .B(G2435), .Z(new_n626));
  XOR2_X1   g201(.A(KEYINPUT74), .B(G2438), .Z(new_n627));
  XOR2_X1   g202(.A(new_n626), .B(new_n627), .Z(new_n628));
  INV_X1    g203(.A(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2427), .B(G2430), .ZN(new_n630));
  INV_X1    g205(.A(new_n630), .ZN(new_n631));
  OAI21_X1  g206(.A(KEYINPUT14), .B1(new_n629), .B2(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT75), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n629), .A2(new_n631), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(G2443), .B(G2446), .Z(new_n636));
  NAND2_X1  g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G1341), .B(G1348), .ZN(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(new_n639));
  INV_X1    g214(.A(new_n636), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n633), .A2(new_n634), .A3(new_n640), .ZN(new_n641));
  AND3_X1   g216(.A1(new_n637), .A2(new_n639), .A3(new_n641), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n639), .B1(new_n637), .B2(new_n641), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2451), .B(G2454), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT16), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n625), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  INV_X1    g222(.A(new_n646), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n648), .B1(new_n642), .B2(new_n643), .ZN(new_n649));
  AND2_X1   g224(.A1(new_n647), .A2(new_n649), .ZN(G401));
  INV_X1    g225(.A(KEYINPUT18), .ZN(new_n651));
  XOR2_X1   g226(.A(G2084), .B(G2090), .Z(new_n652));
  XNOR2_X1  g227(.A(G2067), .B(G2678), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n654), .A2(KEYINPUT17), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n652), .A2(new_n653), .ZN(new_n656));
  OAI21_X1  g231(.A(new_n651), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2100), .ZN(new_n658));
  XOR2_X1   g233(.A(G2072), .B(G2078), .Z(new_n659));
  AOI21_X1  g234(.A(new_n659), .B1(new_n654), .B2(KEYINPUT18), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G2096), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n658), .B(new_n661), .ZN(G227));
  XOR2_X1   g237(.A(G1971), .B(G1976), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT19), .ZN(new_n664));
  XOR2_X1   g239(.A(G1956), .B(G2474), .Z(new_n665));
  XOR2_X1   g240(.A(G1961), .B(G1966), .Z(new_n666));
  AND2_X1   g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT20), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n665), .A2(new_n666), .ZN(new_n670));
  NOR3_X1   g245(.A1(new_n664), .A2(new_n667), .A3(new_n670), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n671), .B1(new_n664), .B2(new_n670), .ZN(new_n672));
  AND2_X1   g247(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G1991), .B(G1996), .Z(new_n676));
  NAND2_X1  g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n673), .A2(new_n674), .ZN(new_n678));
  INV_X1    g253(.A(new_n676), .ZN(new_n679));
  OR2_X1    g254(.A1(new_n673), .A2(new_n674), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n678), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1981), .B(G1986), .ZN(new_n682));
  AND3_X1   g257(.A1(new_n677), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n682), .B1(new_n677), .B2(new_n681), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(G229));
  INV_X1    g260(.A(KEYINPUT93), .ZN(new_n686));
  NAND2_X1  g261(.A1(G162), .A2(G29), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n687), .B1(G29), .B2(G35), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT29), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n686), .B1(new_n690), .B2(G2090), .ZN(new_n691));
  INV_X1    g266(.A(G16), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(G19), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n693), .B1(new_n546), .B2(new_n692), .ZN(new_n694));
  XOR2_X1   g269(.A(KEYINPUT85), .B(G1341), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n692), .A2(G4), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n697), .B1(new_n597), .B2(new_n692), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(G1348), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n692), .A2(G20), .ZN(new_n700));
  XOR2_X1   g275(.A(new_n700), .B(KEYINPUT23), .Z(new_n701));
  AOI21_X1  g276(.A(new_n701), .B1(G299), .B2(G16), .ZN(new_n702));
  XOR2_X1   g277(.A(KEYINPUT94), .B(G1956), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT87), .B(KEYINPUT28), .ZN(new_n705));
  INV_X1    g280(.A(G29), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G26), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n705), .B(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n474), .A2(G140), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n476), .A2(G128), .ZN(new_n710));
  OR2_X1    g285(.A1(new_n461), .A2(G116), .ZN(new_n711));
  INV_X1    g286(.A(G104), .ZN(new_n712));
  AOI22_X1  g287(.A1(new_n711), .A2(KEYINPUT86), .B1(new_n712), .B2(new_n461), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n712), .A2(new_n461), .A3(KEYINPUT86), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G2104), .ZN(new_n715));
  OAI211_X1 g290(.A(new_n709), .B(new_n710), .C1(new_n713), .C2(new_n715), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n708), .B1(new_n716), .B2(G29), .ZN(new_n717));
  INV_X1    g292(.A(G2067), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  NOR4_X1   g294(.A1(new_n696), .A2(new_n699), .A3(new_n704), .A4(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n690), .A2(G2090), .ZN(new_n721));
  INV_X1    g296(.A(G2090), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n689), .A2(KEYINPUT93), .A3(new_n722), .ZN(new_n723));
  NAND4_X1  g298(.A1(new_n691), .A2(new_n720), .A3(new_n721), .A4(new_n723), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT31), .B(G11), .ZN(new_n725));
  INV_X1    g300(.A(KEYINPUT30), .ZN(new_n726));
  AND2_X1   g301(.A1(new_n726), .A2(G28), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n706), .B1(new_n726), .B2(G28), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n621), .A2(new_n706), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT90), .ZN(new_n730));
  OAI221_X1 g305(.A(new_n725), .B1(new_n727), .B2(new_n728), .C1(new_n729), .C2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n692), .A2(G21), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(G168), .B2(new_n692), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(G1966), .ZN(new_n734));
  AOI211_X1 g309(.A(new_n731), .B(new_n734), .C1(new_n730), .C2(new_n729), .ZN(new_n735));
  NOR2_X1   g310(.A1(G5), .A2(G16), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT91), .Z(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G301), .B2(new_n692), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(G1961), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n706), .A2(G33), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n474), .A2(G139), .ZN(new_n741));
  AOI22_X1  g316(.A1(new_n612), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n741), .B1(new_n742), .B2(new_n461), .ZN(new_n743));
  NAND2_X1  g318(.A1(G103), .A2(G2104), .ZN(new_n744));
  OAI21_X1  g319(.A(KEYINPUT88), .B1(new_n744), .B2(G2105), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT88), .ZN(new_n746));
  NAND4_X1  g321(.A1(new_n746), .A2(new_n461), .A3(G103), .A4(G2104), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT25), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n745), .A2(new_n747), .A3(KEYINPUT25), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n743), .A2(new_n752), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n740), .B1(new_n753), .B2(new_n706), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(G2072), .Z(new_n755));
  NAND3_X1  g330(.A1(new_n735), .A2(new_n739), .A3(new_n755), .ZN(new_n756));
  AOI22_X1  g331(.A1(new_n474), .A2(G141), .B1(G105), .B2(new_n468), .ZN(new_n757));
  NAND3_X1  g332(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT26), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND4_X1  g335(.A1(KEYINPUT26), .A2(G117), .A3(G2104), .A4(G2105), .ZN(new_n761));
  AOI22_X1  g336(.A1(new_n476), .A2(G129), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n757), .A2(new_n762), .ZN(new_n763));
  MUX2_X1   g338(.A(G32), .B(new_n763), .S(G29), .Z(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT27), .ZN(new_n765));
  INV_X1    g340(.A(G1996), .ZN(new_n766));
  OR2_X1    g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n765), .A2(new_n766), .ZN(new_n768));
  NAND2_X1  g343(.A1(G164), .A2(G29), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G27), .B2(G29), .ZN(new_n770));
  INV_X1    g345(.A(G2078), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(G2084), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT89), .B(KEYINPUT24), .ZN(new_n774));
  INV_X1    g349(.A(new_n774), .ZN(new_n775));
  AOI21_X1  g350(.A(G29), .B1(new_n775), .B2(G34), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G34), .B2(new_n775), .ZN(new_n777));
  OAI21_X1  g352(.A(G29), .B1(new_n466), .B2(new_n470), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n772), .B1(new_n773), .B2(new_n780), .ZN(new_n781));
  AOI22_X1  g356(.A1(new_n770), .A2(new_n771), .B1(G2084), .B2(new_n779), .ZN(new_n782));
  NAND4_X1  g357(.A1(new_n767), .A2(new_n768), .A3(new_n781), .A4(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n756), .A2(new_n783), .ZN(new_n784));
  OR2_X1    g359(.A1(new_n784), .A2(KEYINPUT92), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n784), .A2(KEYINPUT92), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n724), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT84), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n692), .A2(G23), .ZN(new_n789));
  INV_X1    g364(.A(KEYINPUT80), .ZN(new_n790));
  XNOR2_X1  g365(.A(G288), .B(new_n790), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n789), .B1(new_n791), .B2(new_n692), .ZN(new_n792));
  XOR2_X1   g367(.A(KEYINPUT33), .B(G1976), .Z(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT81), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n792), .B(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(G6), .A2(G16), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(new_n575), .B2(G16), .ZN(new_n797));
  XOR2_X1   g372(.A(KEYINPUT32), .B(G1981), .Z(new_n798));
  XOR2_X1   g373(.A(new_n797), .B(new_n798), .Z(new_n799));
  NAND2_X1  g374(.A1(new_n692), .A2(G22), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G166), .B2(new_n692), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT82), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n799), .B1(G1971), .B2(new_n803), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n803), .A2(G1971), .ZN(new_n805));
  AND3_X1   g380(.A1(new_n795), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(KEYINPUT34), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n788), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n692), .A2(G24), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(new_n582), .B2(new_n692), .ZN(new_n810));
  XOR2_X1   g385(.A(new_n810), .B(KEYINPUT79), .Z(new_n811));
  INV_X1    g386(.A(G1986), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT78), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n706), .A2(G25), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n461), .A2(G107), .ZN(new_n816));
  OAI21_X1  g391(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  AOI22_X1  g393(.A1(new_n476), .A2(G119), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT76), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n820), .B1(new_n474), .B2(G131), .ZN(new_n821));
  OAI211_X1 g396(.A(G131), .B(new_n461), .C1(new_n462), .C2(new_n463), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n822), .A2(KEYINPUT76), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n819), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT77), .ZN(new_n825));
  INV_X1    g400(.A(new_n825), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n815), .B1(new_n826), .B2(new_n706), .ZN(new_n827));
  XOR2_X1   g402(.A(KEYINPUT35), .B(G1991), .Z(new_n828));
  AND2_X1   g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n827), .A2(new_n828), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n814), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  AND2_X1   g406(.A1(new_n813), .A2(new_n831), .ZN(new_n832));
  NAND4_X1  g407(.A1(new_n795), .A2(new_n804), .A3(new_n807), .A4(new_n805), .ZN(new_n833));
  OR2_X1    g408(.A1(new_n827), .A2(new_n828), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n827), .A2(new_n828), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n834), .A2(KEYINPUT78), .A3(new_n835), .ZN(new_n836));
  NAND4_X1  g411(.A1(new_n832), .A2(KEYINPUT83), .A3(new_n833), .A4(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT83), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n813), .A2(new_n831), .A3(new_n836), .ZN(new_n839));
  INV_X1    g414(.A(new_n833), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n838), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n808), .B1(new_n837), .B2(new_n841), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n787), .B1(new_n842), .B2(KEYINPUT36), .ZN(new_n843));
  AND2_X1   g418(.A1(new_n842), .A2(KEYINPUT36), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n843), .A2(new_n844), .ZN(G311));
  OR2_X1    g420(.A1(new_n842), .A2(KEYINPUT36), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n842), .A2(KEYINPUT36), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n846), .A2(new_n847), .A3(new_n787), .ZN(G150));
  AOI22_X1  g423(.A1(new_n498), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n849), .A2(new_n500), .ZN(new_n850));
  INV_X1    g425(.A(G93), .ZN(new_n851));
  INV_X1    g426(.A(G55), .ZN(new_n852));
  OAI22_X1  g427(.A1(new_n503), .A2(new_n851), .B1(new_n505), .B2(new_n852), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(G860), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n856), .B(KEYINPUT37), .Z(new_n857));
  OAI21_X1  g432(.A(new_n855), .B1(new_n539), .B2(new_n545), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n854), .A2(new_n538), .A3(new_n534), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT38), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n597), .A2(G559), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n861), .B(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT39), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(G860), .B1(new_n865), .B2(KEYINPUT95), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n866), .B1(KEYINPUT95), .B2(new_n865), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n863), .A2(new_n864), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT96), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n857), .B1(new_n867), .B2(new_n869), .ZN(G145));
  INV_X1    g445(.A(KEYINPUT40), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n621), .B(G160), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(G162), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT100), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n490), .A2(new_n492), .ZN(new_n875));
  AND2_X1   g450(.A1(new_n482), .A2(new_n485), .ZN(new_n876));
  AND4_X1   g451(.A1(new_n875), .A2(new_n876), .A3(new_n757), .A4(new_n762), .ZN(new_n877));
  AOI22_X1  g452(.A1(new_n875), .A2(new_n876), .B1(new_n757), .B2(new_n762), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n753), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT97), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n716), .B(new_n880), .ZN(new_n881));
  AND2_X1   g456(.A1(new_n612), .A2(G127), .ZN(new_n882));
  AND2_X1   g457(.A1(G115), .A2(G2104), .ZN(new_n883));
  OAI21_X1  g458(.A(G2105), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND4_X1  g459(.A1(new_n884), .A2(new_n741), .A3(new_n751), .A4(new_n750), .ZN(new_n885));
  INV_X1    g460(.A(new_n492), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n491), .B1(new_n612), .B2(new_n488), .ZN(new_n887));
  OAI211_X1 g462(.A(new_n482), .B(new_n485), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n888), .A2(new_n763), .ZN(new_n889));
  NAND4_X1  g464(.A1(new_n875), .A2(new_n876), .A3(new_n757), .A4(new_n762), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n885), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  AND3_X1   g466(.A1(new_n879), .A2(new_n881), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n881), .B1(new_n879), .B2(new_n891), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  OR3_X1    g469(.A1(new_n461), .A2(KEYINPUT98), .A3(G118), .ZN(new_n895));
  OAI21_X1  g470(.A(KEYINPUT98), .B1(new_n461), .B2(G118), .ZN(new_n896));
  OR2_X1    g471(.A1(G106), .A2(G2105), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n895), .A2(G2104), .A3(new_n896), .A4(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n476), .A2(G130), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n474), .A2(G142), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT99), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n824), .A2(new_n902), .ZN(new_n903));
  OAI211_X1 g478(.A(new_n819), .B(KEYINPUT99), .C1(new_n821), .C2(new_n823), .ZN(new_n904));
  AND3_X1   g479(.A1(new_n903), .A2(new_n904), .A3(new_n614), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n614), .B1(new_n903), .B2(new_n904), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n901), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n903), .A2(new_n904), .ZN(new_n908));
  INV_X1    g483(.A(new_n614), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n901), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n903), .A2(new_n904), .A3(new_n614), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n907), .A2(new_n913), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n874), .B1(new_n894), .B2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n881), .ZN(new_n916));
  NOR3_X1   g491(.A1(new_n877), .A2(new_n878), .A3(new_n753), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n885), .B1(new_n889), .B2(new_n890), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n916), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n879), .A2(new_n881), .A3(new_n891), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n921), .A2(KEYINPUT100), .A3(new_n913), .A4(new_n907), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT101), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n915), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n894), .A2(new_n914), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n923), .B1(new_n915), .B2(new_n922), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n873), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT103), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT102), .ZN(new_n930));
  AOI22_X1  g505(.A1(new_n921), .A2(new_n930), .B1(new_n913), .B2(new_n907), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n894), .A2(KEYINPUT102), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n873), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n915), .A2(new_n922), .ZN(new_n934));
  AOI21_X1  g509(.A(G37), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n928), .A2(new_n929), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n929), .B1(new_n928), .B2(new_n935), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n871), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n928), .A2(new_n935), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(KEYINPUT103), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n928), .A2(new_n929), .A3(new_n935), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n940), .A2(KEYINPUT40), .A3(new_n941), .ZN(new_n942));
  AND2_X1   g517(.A1(new_n938), .A2(new_n942), .ZN(G395));
  XOR2_X1   g518(.A(new_n860), .B(new_n608), .Z(new_n944));
  INV_X1    g519(.A(new_n559), .ZN(new_n945));
  INV_X1    g520(.A(G91), .ZN(new_n946));
  OAI22_X1  g521(.A1(new_n561), .A2(new_n500), .B1(new_n946), .B2(new_n503), .ZN(new_n947));
  OR3_X1    g522(.A1(new_n945), .A2(new_n947), .A3(KEYINPUT104), .ZN(new_n948));
  NAND2_X1  g523(.A1(G299), .A2(KEYINPUT104), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n948), .A2(new_n597), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n591), .A2(new_n596), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n951), .A2(KEYINPUT104), .A3(G299), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  OR2_X1    g529(.A1(new_n944), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT41), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n953), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n950), .A2(KEYINPUT41), .A3(new_n952), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n944), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n955), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(KEYINPUT42), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n791), .B(new_n575), .ZN(new_n963));
  XNOR2_X1  g538(.A(G166), .B(new_n582), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n791), .B(G305), .ZN(new_n966));
  INV_X1    g541(.A(new_n964), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n965), .A2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  AND2_X1   g545(.A1(new_n970), .A2(KEYINPUT105), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT42), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n955), .A2(new_n972), .A3(new_n960), .ZN(new_n973));
  AND3_X1   g548(.A1(new_n962), .A2(new_n971), .A3(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n971), .B1(new_n962), .B2(new_n973), .ZN(new_n975));
  OAI21_X1  g550(.A(G868), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n976), .B1(G868), .B2(new_n854), .ZN(G295));
  OAI21_X1  g552(.A(new_n976), .B1(G868), .B2(new_n854), .ZN(G331));
  NAND2_X1  g553(.A1(G301), .A2(G286), .ZN(new_n979));
  NAND3_X1  g554(.A1(G168), .A2(new_n525), .A3(new_n531), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n858), .A2(new_n859), .A3(new_n979), .A4(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n534), .A2(KEYINPUT67), .A3(new_n538), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n544), .B1(new_n542), .B2(new_n543), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n854), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NOR4_X1   g559(.A1(new_n542), .A2(new_n850), .A3(new_n853), .A4(new_n543), .ZN(new_n985));
  INV_X1    g560(.A(new_n980), .ZN(new_n986));
  AOI21_X1  g561(.A(G168), .B1(new_n525), .B2(new_n531), .ZN(new_n987));
  OAI22_X1  g562(.A1(new_n984), .A2(new_n985), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(KEYINPUT106), .B1(new_n981), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT106), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n979), .A2(new_n980), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n990), .B1(new_n860), .B2(new_n991), .ZN(new_n992));
  OAI211_X1 g567(.A(new_n958), .B(new_n957), .C1(new_n989), .C2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT107), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n954), .A2(new_n994), .A3(new_n988), .A4(new_n981), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n981), .A2(new_n988), .ZN(new_n996));
  OAI21_X1  g571(.A(KEYINPUT107), .B1(new_n996), .B2(new_n953), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n993), .A2(new_n969), .A3(new_n995), .A4(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(G37), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  AND2_X1   g575(.A1(new_n995), .A2(new_n997), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n969), .B1(new_n1001), .B2(new_n993), .ZN(new_n1002));
  OR3_X1    g577(.A1(new_n1000), .A2(new_n1002), .A3(KEYINPUT43), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n959), .B1(new_n988), .B2(new_n981), .ZN(new_n1004));
  NOR3_X1   g579(.A1(new_n989), .A2(new_n992), .A3(new_n953), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n970), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  AND3_X1   g581(.A1(new_n1006), .A2(new_n999), .A3(new_n998), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT43), .ZN(new_n1008));
  OAI211_X1 g583(.A(new_n1003), .B(KEYINPUT44), .C1(new_n1007), .C2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g584(.A(KEYINPUT43), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n1006), .A2(new_n998), .A3(new_n1008), .A4(new_n999), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT44), .ZN(new_n1013));
  AOI21_X1  g588(.A(KEYINPUT108), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT108), .ZN(new_n1015));
  AOI211_X1 g590(.A(new_n1015), .B(KEYINPUT44), .C1(new_n1010), .C2(new_n1011), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1009), .B1(new_n1014), .B2(new_n1016), .ZN(G397));
  NAND2_X1  g592(.A1(new_n582), .A2(new_n812), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(KEYINPUT110), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n582), .A2(new_n812), .ZN(new_n1020));
  XNOR2_X1  g595(.A(new_n1019), .B(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(G1384), .B1(new_n875), .B2(new_n876), .ZN(new_n1022));
  AND2_X1   g597(.A1(new_n1022), .A2(KEYINPUT109), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT45), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1024), .B1(new_n1022), .B2(KEYINPUT109), .ZN(new_n1025));
  INV_X1    g600(.A(G40), .ZN(new_n1026));
  NOR3_X1   g601(.A1(new_n466), .A2(new_n470), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1027), .ZN(new_n1028));
  NOR3_X1   g603(.A1(new_n1023), .A2(new_n1025), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1021), .A2(new_n1030), .ZN(new_n1031));
  XNOR2_X1  g606(.A(new_n1031), .B(KEYINPUT111), .ZN(new_n1032));
  XNOR2_X1  g607(.A(new_n763), .B(new_n766), .ZN(new_n1033));
  XNOR2_X1  g608(.A(new_n716), .B(new_n718), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1035), .ZN(new_n1036));
  XNOR2_X1  g611(.A(new_n824), .B(new_n828), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1030), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1032), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT62), .ZN(new_n1040));
  INV_X1    g615(.A(G1966), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1024), .A2(G1384), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1027), .B1(G164), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(G1384), .ZN(new_n1045));
  AOI21_X1  g620(.A(KEYINPUT45), .B1(new_n888), .B2(new_n1045), .ZN(new_n1046));
  OAI211_X1 g621(.A(KEYINPUT118), .B(new_n1041), .C1(new_n1044), .C2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g622(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT50), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n888), .A2(new_n1049), .A3(new_n1045), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1048), .A2(new_n1050), .A3(new_n773), .A4(new_n1027), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1047), .A2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1024), .B1(G164), .B2(G1384), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n888), .A2(new_n1042), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1053), .A2(new_n1027), .A3(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(KEYINPUT118), .B1(new_n1055), .B2(new_n1041), .ZN(new_n1056));
  OAI21_X1  g631(.A(G286), .B1(new_n1052), .B2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1041), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT118), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1060), .A2(G168), .A3(new_n1051), .A4(new_n1047), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1057), .A2(G8), .A3(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(KEYINPUT51), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT124), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT51), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1061), .A2(new_n1065), .A3(G8), .ZN(new_n1066));
  AND3_X1   g641(.A1(new_n1063), .A2(new_n1064), .A3(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1064), .B1(new_n1063), .B2(new_n1066), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1040), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(G8), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1052), .A2(new_n1056), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1070), .B1(new_n1071), .B2(G168), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1065), .B1(new_n1072), .B2(new_n1057), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1066), .ZN(new_n1074));
  OAI21_X1  g649(.A(KEYINPUT124), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1063), .A2(new_n1064), .A3(new_n1066), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1075), .A2(KEYINPUT62), .A3(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(G288), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(new_n790), .ZN(new_n1079));
  NAND2_X1  g654(.A1(G288), .A2(KEYINPUT80), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1079), .A2(G1976), .A3(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(G1976), .ZN(new_n1082));
  AOI21_X1  g657(.A(KEYINPUT52), .B1(G288), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1022), .A2(new_n1027), .ZN(new_n1084));
  AOI21_X1  g659(.A(KEYINPUT115), .B1(new_n1084), .B2(G8), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT115), .ZN(new_n1086));
  AOI211_X1 g661(.A(new_n1086), .B(new_n1070), .C1(new_n1022), .C2(new_n1027), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1081), .B(new_n1083), .C1(new_n1085), .C2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(G1981), .B1(new_n571), .B2(new_n574), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n526), .A2(G86), .ZN(new_n1090));
  INV_X1    g665(.A(G61), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1091), .B1(new_n496), .B2(new_n497), .ZN(new_n1092));
  INV_X1    g667(.A(new_n573), .ZN(new_n1093));
  OAI21_X1  g668(.A(G651), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  XOR2_X1   g669(.A(KEYINPUT116), .B(G1981), .Z(new_n1095));
  NAND4_X1  g670(.A1(new_n1090), .A2(new_n1094), .A3(new_n569), .A4(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(KEYINPUT117), .B1(new_n1089), .B2(new_n1096), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1097), .A2(KEYINPUT49), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT49), .ZN(new_n1099));
  AOI211_X1 g674(.A(KEYINPUT117), .B(new_n1099), .C1(new_n1089), .C2(new_n1096), .ZN(new_n1100));
  OAI22_X1  g675(.A1(new_n1098), .A2(new_n1100), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1085), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1087), .ZN(new_n1103));
  AOI22_X1  g678(.A1(new_n1102), .A2(new_n1103), .B1(G1976), .B2(new_n791), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT52), .ZN(new_n1105));
  OAI211_X1 g680(.A(new_n1088), .B(new_n1101), .C1(new_n1104), .C2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT55), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1107), .A2(KEYINPUT112), .ZN(new_n1108));
  XNOR2_X1  g683(.A(new_n1108), .B(KEYINPUT113), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1070), .B1(KEYINPUT112), .B2(new_n1107), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1109), .B1(G303), .B2(new_n1110), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n1110), .B(new_n1109), .C1(new_n501), .C2(new_n507), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1112), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1048), .A2(new_n1027), .A3(new_n1050), .ZN(new_n1116));
  OAI22_X1  g691(.A1(new_n1115), .A2(G1971), .B1(new_n1116), .B2(G2090), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1114), .B1(new_n1117), .B2(G8), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1106), .A2(new_n1118), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1053), .A2(new_n771), .A3(new_n1027), .A4(new_n1054), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT125), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT53), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(G1961), .ZN(new_n1125));
  AOI22_X1  g700(.A1(new_n1120), .A2(new_n1124), .B1(new_n1116), .B2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1115), .A2(new_n771), .A3(new_n1123), .ZN(new_n1127));
  AOI21_X1  g702(.A(G301), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1116), .A2(G2090), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1044), .ZN(new_n1130));
  AOI21_X1  g705(.A(G1971), .B1(new_n1130), .B2(new_n1053), .ZN(new_n1131));
  OAI211_X1 g706(.A(new_n1114), .B(G8), .C1(new_n1129), .C2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT114), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1117), .A2(KEYINPUT114), .A3(G8), .A4(new_n1114), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  AND3_X1   g711(.A1(new_n1119), .A2(new_n1128), .A3(new_n1136), .ZN(new_n1137));
  AND3_X1   g712(.A1(new_n1069), .A2(new_n1077), .A3(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1139));
  AND3_X1   g714(.A1(new_n1101), .A2(new_n1082), .A3(new_n1078), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1096), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1139), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1142), .B1(new_n1136), .B2(new_n1106), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1105), .B1(new_n1139), .B2(new_n1081), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1101), .A2(new_n1088), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NOR3_X1   g721(.A1(new_n1071), .A2(new_n1070), .A3(G286), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1118), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1136), .A2(new_n1146), .A3(new_n1147), .A4(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT63), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1119), .A2(KEYINPUT63), .A3(new_n1136), .A4(new_n1147), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1143), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT54), .ZN(new_n1154));
  XOR2_X1   g729(.A(KEYINPUT126), .B(G2078), .Z(new_n1155));
  NOR2_X1   g730(.A1(new_n1155), .A2(new_n1122), .ZN(new_n1156));
  OAI211_X1 g731(.A(new_n1130), .B(new_n1156), .C1(new_n1023), .C2(new_n1025), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1116), .A2(new_n1125), .ZN(new_n1159));
  AND4_X1   g734(.A1(G301), .A2(new_n1157), .A3(new_n1158), .A4(new_n1159), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1154), .B1(new_n1160), .B2(new_n1128), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1157), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT127), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1157), .A2(new_n1158), .A3(KEYINPUT127), .A4(new_n1159), .ZN(new_n1165));
  AOI21_X1  g740(.A(G301), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1126), .A2(G301), .A3(new_n1127), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1167), .A2(KEYINPUT54), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1161), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1136), .A2(new_n1146), .A3(new_n1148), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT119), .ZN(new_n1172));
  AND3_X1   g747(.A1(new_n557), .A2(new_n1172), .A3(new_n558), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1172), .B1(new_n557), .B2(new_n558), .ZN(new_n1174));
  NOR3_X1   g749(.A1(new_n1173), .A2(new_n1174), .A3(KEYINPUT57), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n947), .A2(KEYINPUT120), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT120), .ZN(new_n1177));
  OAI221_X1 g752(.A(new_n1177), .B1(new_n503), .B2(new_n946), .C1(new_n561), .C2(new_n500), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1176), .A2(new_n1178), .ZN(new_n1179));
  AOI22_X1  g754(.A1(new_n1175), .A2(new_n1179), .B1(KEYINPUT57), .B2(G299), .ZN(new_n1180));
  INV_X1    g755(.A(G1956), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1116), .A2(new_n1181), .ZN(new_n1182));
  XNOR2_X1  g757(.A(KEYINPUT56), .B(G2072), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1130), .A2(new_n1053), .A3(new_n1183), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1180), .B1(new_n1182), .B2(new_n1184), .ZN(new_n1185));
  AND3_X1   g760(.A1(new_n1182), .A2(new_n1180), .A3(new_n1184), .ZN(new_n1186));
  INV_X1    g761(.A(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(G1348), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1116), .A2(new_n1188), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1022), .A2(new_n718), .A3(new_n1027), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n951), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1185), .B1(new_n1187), .B2(new_n1191), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT123), .ZN(new_n1193));
  OAI211_X1 g768(.A(new_n1193), .B(KEYINPUT61), .C1(new_n1186), .C2(new_n1185), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1182), .A2(new_n1184), .ZN(new_n1195));
  INV_X1    g770(.A(new_n1180), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1195), .A2(new_n1193), .A3(new_n1196), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT61), .ZN(new_n1198));
  NAND4_X1  g773(.A1(new_n1182), .A2(new_n1180), .A3(new_n1184), .A4(new_n1193), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n1197), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  AND2_X1   g775(.A1(new_n1194), .A2(new_n1200), .ZN(new_n1201));
  AND3_X1   g776(.A1(new_n1189), .A2(new_n951), .A3(new_n1190), .ZN(new_n1202));
  OAI21_X1  g777(.A(KEYINPUT60), .B1(new_n1202), .B2(new_n1191), .ZN(new_n1203));
  NOR2_X1   g778(.A1(new_n951), .A2(KEYINPUT60), .ZN(new_n1204));
  NAND3_X1  g779(.A1(new_n1189), .A2(new_n1190), .A3(new_n1204), .ZN(new_n1205));
  XOR2_X1   g780(.A(KEYINPUT58), .B(G1341), .Z(new_n1206));
  NAND2_X1  g781(.A1(new_n1084), .A2(new_n1206), .ZN(new_n1207));
  INV_X1    g782(.A(KEYINPUT121), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  NAND3_X1  g784(.A1(new_n1084), .A2(KEYINPUT121), .A3(new_n1206), .ZN(new_n1210));
  OAI211_X1 g785(.A(new_n1209), .B(new_n1210), .C1(G1996), .C2(new_n1055), .ZN(new_n1211));
  INV_X1    g786(.A(KEYINPUT122), .ZN(new_n1212));
  OR2_X1    g787(.A1(new_n1212), .A2(KEYINPUT59), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1212), .A2(KEYINPUT59), .ZN(new_n1214));
  AOI22_X1  g789(.A1(new_n1211), .A2(new_n546), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  OAI21_X1  g790(.A(new_n1210), .B1(new_n1055), .B2(G1996), .ZN(new_n1216));
  AOI21_X1  g791(.A(KEYINPUT121), .B1(new_n1084), .B2(new_n1206), .ZN(new_n1217));
  OAI211_X1 g792(.A(new_n546), .B(new_n1214), .C1(new_n1216), .C2(new_n1217), .ZN(new_n1218));
  INV_X1    g793(.A(new_n1218), .ZN(new_n1219));
  OAI211_X1 g794(.A(new_n1203), .B(new_n1205), .C1(new_n1215), .C2(new_n1219), .ZN(new_n1220));
  OAI21_X1  g795(.A(new_n1192), .B1(new_n1201), .B2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g796(.A1(new_n1171), .A2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g797(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1223));
  OAI21_X1  g798(.A(new_n1153), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  OAI21_X1  g799(.A(new_n1039), .B1(new_n1138), .B2(new_n1224), .ZN(new_n1225));
  NOR2_X1   g800(.A1(new_n1030), .A2(new_n1018), .ZN(new_n1226));
  AND2_X1   g801(.A1(new_n1226), .A2(KEYINPUT48), .ZN(new_n1227));
  NOR2_X1   g802(.A1(new_n1226), .A2(KEYINPUT48), .ZN(new_n1228));
  NOR3_X1   g803(.A1(new_n1227), .A2(new_n1228), .A3(new_n1038), .ZN(new_n1229));
  INV_X1    g804(.A(new_n1034), .ZN(new_n1230));
  OAI21_X1  g805(.A(new_n1029), .B1(new_n763), .B2(new_n1230), .ZN(new_n1231));
  NOR3_X1   g806(.A1(new_n1030), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1232));
  INV_X1    g807(.A(KEYINPUT46), .ZN(new_n1233));
  AOI21_X1  g808(.A(new_n1233), .B1(new_n1029), .B2(new_n766), .ZN(new_n1234));
  OAI21_X1  g809(.A(new_n1231), .B1(new_n1232), .B2(new_n1234), .ZN(new_n1235));
  XOR2_X1   g810(.A(new_n1235), .B(KEYINPUT47), .Z(new_n1236));
  NAND3_X1  g811(.A1(new_n1036), .A2(new_n826), .A3(new_n828), .ZN(new_n1237));
  OAI21_X1  g812(.A(new_n1237), .B1(G2067), .B2(new_n716), .ZN(new_n1238));
  AOI211_X1 g813(.A(new_n1229), .B(new_n1236), .C1(new_n1029), .C2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g814(.A1(new_n1225), .A2(new_n1239), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g815(.A1(new_n940), .A2(new_n941), .ZN(new_n1242));
  NOR2_X1   g816(.A1(G227), .A2(new_n459), .ZN(new_n1243));
  OAI21_X1  g817(.A(new_n1243), .B1(new_n683), .B2(new_n684), .ZN(new_n1244));
  AOI21_X1  g818(.A(new_n1244), .B1(new_n647), .B2(new_n649), .ZN(new_n1245));
  AND3_X1   g819(.A1(new_n1242), .A2(new_n1012), .A3(new_n1245), .ZN(G308));
  NAND3_X1  g820(.A1(new_n1242), .A2(new_n1012), .A3(new_n1245), .ZN(G225));
endmodule


