//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 0 0 1 1 1 0 0 0 1 0 0 0 0 1 1 0 1 0 0 1 1 1 1 1 0 0 1 0 0 0 0 0 0 0 0 1 0 0 1 1 0 1 0 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:23 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002;
  INV_X1    g000(.A(KEYINPUT30), .ZN(new_n187));
  XNOR2_X1  g001(.A(G143), .B(G146), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT0), .ZN(new_n189));
  INV_X1    g003(.A(G128), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n188), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  XOR2_X1   g005(.A(KEYINPUT0), .B(G128), .Z(new_n192));
  OAI21_X1  g006(.A(new_n191), .B1(new_n188), .B2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT64), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  OAI211_X1 g009(.A(new_n191), .B(KEYINPUT64), .C1(new_n188), .C2(new_n192), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT11), .ZN(new_n198));
  INV_X1    g012(.A(G134), .ZN(new_n199));
  NOR3_X1   g013(.A1(new_n198), .A2(new_n199), .A3(G137), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  AND2_X1   g015(.A1(KEYINPUT65), .A2(G134), .ZN(new_n202));
  NOR2_X1   g016(.A1(KEYINPUT65), .A2(G134), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G137), .ZN(new_n205));
  INV_X1    g019(.A(G137), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n206), .B1(new_n202), .B2(new_n203), .ZN(new_n207));
  AND3_X1   g021(.A1(new_n207), .A2(KEYINPUT66), .A3(new_n198), .ZN(new_n208));
  AOI21_X1  g022(.A(KEYINPUT66), .B1(new_n207), .B2(new_n198), .ZN(new_n209));
  OAI211_X1 g023(.A(new_n201), .B(new_n205), .C1(new_n208), .C2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G131), .ZN(new_n211));
  AOI21_X1  g025(.A(G131), .B1(new_n204), .B2(G137), .ZN(new_n212));
  OAI211_X1 g026(.A(new_n201), .B(new_n212), .C1(new_n208), .C2(new_n209), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n197), .B1(new_n211), .B2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT65), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(new_n199), .ZN(new_n216));
  NAND2_X1  g030(.A1(KEYINPUT65), .A2(G134), .ZN(new_n217));
  AOI21_X1  g031(.A(G137), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n206), .A2(G134), .ZN(new_n219));
  OAI21_X1  g033(.A(G131), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT67), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI211_X1 g036(.A(KEYINPUT67), .B(G131), .C1(new_n218), .C2(new_n219), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(G146), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G143), .ZN(new_n226));
  INV_X1    g040(.A(G143), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G146), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  OR3_X1    g043(.A1(new_n229), .A2(KEYINPUT1), .A3(new_n190), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n190), .B1(new_n226), .B2(KEYINPUT1), .ZN(new_n231));
  NOR3_X1   g045(.A1(new_n231), .A2(new_n188), .A3(KEYINPUT68), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT68), .ZN(new_n233));
  OAI21_X1  g047(.A(KEYINPUT1), .B1(new_n227), .B2(G146), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(G128), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n233), .B1(new_n235), .B2(new_n229), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n230), .B1(new_n232), .B2(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n224), .A2(new_n213), .A3(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n187), .B1(new_n214), .B2(new_n239), .ZN(new_n240));
  XNOR2_X1  g054(.A(G116), .B(G119), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(KEYINPUT69), .ZN(new_n243));
  XNOR2_X1  g057(.A(KEYINPUT2), .B(G113), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  XNOR2_X1  g059(.A(new_n243), .B(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n240), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(G131), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT66), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n250), .B1(new_n218), .B2(KEYINPUT11), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n207), .A2(KEYINPUT66), .A3(new_n198), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n200), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n249), .B1(new_n253), .B2(new_n205), .ZN(new_n254));
  INV_X1    g068(.A(new_n213), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n193), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n238), .A2(KEYINPUT70), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT70), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n224), .A2(new_n213), .A3(new_n258), .A4(new_n237), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n256), .A2(new_n257), .A3(KEYINPUT30), .A4(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT71), .ZN(new_n261));
  AND2_X1   g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n260), .A2(new_n261), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n248), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT31), .ZN(new_n265));
  INV_X1    g079(.A(new_n246), .ZN(new_n266));
  NAND4_X1  g080(.A1(new_n256), .A2(new_n257), .A3(new_n259), .A4(new_n266), .ZN(new_n267));
  XNOR2_X1  g081(.A(KEYINPUT26), .B(G101), .ZN(new_n268));
  INV_X1    g082(.A(G237), .ZN(new_n269));
  INV_X1    g083(.A(G953), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n269), .A2(new_n270), .A3(G210), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n268), .B(new_n271), .ZN(new_n272));
  XNOR2_X1  g086(.A(KEYINPUT72), .B(KEYINPUT27), .ZN(new_n273));
  XNOR2_X1  g087(.A(new_n272), .B(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n267), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n264), .A2(new_n265), .A3(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(KEYINPUT68), .B1(new_n231), .B2(new_n188), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n235), .A2(new_n233), .A3(new_n229), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AOI22_X1  g094(.A1(new_n222), .A2(new_n223), .B1(new_n280), .B2(new_n230), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n258), .B1(new_n281), .B2(new_n213), .ZN(new_n282));
  AND4_X1   g096(.A1(new_n258), .A2(new_n224), .A3(new_n213), .A4(new_n237), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n284), .A2(KEYINPUT71), .A3(KEYINPUT30), .A4(new_n256), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n260), .A2(new_n261), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n247), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(KEYINPUT31), .B1(new_n287), .B2(new_n275), .ZN(new_n288));
  INV_X1    g102(.A(new_n274), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT28), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n246), .B1(new_n214), .B2(new_n239), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n290), .B1(new_n267), .B2(new_n291), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n239), .A2(new_n246), .ZN(new_n293));
  AOI21_X1  g107(.A(KEYINPUT28), .B1(new_n293), .B2(new_n256), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n289), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n277), .A2(new_n288), .A3(new_n295), .ZN(new_n296));
  NOR2_X1   g110(.A1(G472), .A2(G902), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  XNOR2_X1  g112(.A(KEYINPUT73), .B(KEYINPUT32), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n296), .A2(KEYINPUT32), .A3(new_n297), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n264), .A2(new_n267), .A3(new_n289), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n274), .B1(new_n292), .B2(new_n294), .ZN(new_n304));
  AOI21_X1  g118(.A(KEYINPUT29), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G902), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n256), .A2(new_n257), .A3(new_n259), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(new_n246), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n290), .B1(new_n308), .B2(new_n267), .ZN(new_n309));
  OR2_X1    g123(.A1(new_n309), .A2(new_n294), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n274), .A2(KEYINPUT29), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n306), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  OAI21_X1  g126(.A(G472), .B1(new_n305), .B2(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n301), .A2(new_n302), .A3(new_n313), .ZN(new_n314));
  XNOR2_X1  g128(.A(G125), .B(G140), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT16), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT16), .ZN(new_n317));
  INV_X1    g131(.A(G140), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n317), .A2(new_n318), .A3(G125), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(new_n225), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n318), .A2(G125), .ZN(new_n322));
  INV_X1    g136(.A(G125), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G140), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  OAI211_X1 g139(.A(G146), .B(new_n319), .C1(new_n325), .C2(new_n317), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n321), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G110), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n190), .A2(G119), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT23), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  OR2_X1    g145(.A1(new_n190), .A2(G119), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n190), .A2(KEYINPUT23), .A3(G119), .ZN(new_n333));
  AND3_X1   g147(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n332), .A2(new_n329), .ZN(new_n335));
  XNOR2_X1  g149(.A(KEYINPUT24), .B(G110), .ZN(new_n336));
  OAI221_X1 g150(.A(new_n327), .B1(new_n328), .B2(new_n334), .C1(new_n335), .C2(new_n336), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n325), .A2(G146), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n334), .A2(new_n328), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n335), .A2(new_n336), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n338), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT74), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n326), .A2(new_n342), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n316), .A2(KEYINPUT74), .A3(G146), .A4(new_n319), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n341), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n337), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n270), .A2(G221), .A3(G234), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n347), .B(KEYINPUT75), .ZN(new_n348));
  XNOR2_X1  g162(.A(KEYINPUT22), .B(G137), .ZN(new_n349));
  XNOR2_X1  g163(.A(new_n348), .B(new_n349), .ZN(new_n350));
  OR2_X1    g164(.A1(new_n346), .A2(new_n350), .ZN(new_n351));
  XOR2_X1   g165(.A(new_n350), .B(KEYINPUT76), .Z(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(new_n346), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n351), .A2(new_n306), .A3(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT25), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n354), .B(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(G217), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n357), .B1(G234), .B2(new_n306), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n358), .A2(G902), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n351), .A2(new_n353), .A3(new_n360), .ZN(new_n361));
  AND2_X1   g175(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n314), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(KEYINPUT77), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT77), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n314), .A2(new_n365), .A3(new_n362), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  XNOR2_X1  g181(.A(KEYINPUT9), .B(G234), .ZN(new_n368));
  NOR3_X1   g182(.A1(new_n368), .A2(new_n357), .A3(G953), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT94), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n370), .B1(new_n190), .B2(G143), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n227), .A2(KEYINPUT94), .A3(G128), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n190), .A2(G143), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n373), .A2(new_n204), .A3(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(G122), .ZN(new_n377));
  OAI21_X1  g191(.A(KEYINPUT93), .B1(new_n377), .B2(G116), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT93), .ZN(new_n379));
  INV_X1    g193(.A(G116), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n379), .A2(new_n380), .A3(G122), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n377), .A2(G116), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  OR2_X1    g198(.A1(KEYINPUT78), .A2(G107), .ZN(new_n385));
  NAND2_X1  g199(.A1(KEYINPUT78), .A2(G107), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  AND2_X1   g202(.A1(KEYINPUT78), .A2(G107), .ZN(new_n389));
  NOR2_X1   g203(.A1(KEYINPUT78), .A2(G107), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n382), .A2(new_n391), .A3(new_n383), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n376), .B1(new_n388), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT13), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n374), .B1(new_n373), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n373), .A2(new_n394), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT95), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n373), .A2(KEYINPUT95), .A3(new_n394), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n395), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n393), .B1(new_n400), .B2(new_n199), .ZN(new_n401));
  INV_X1    g215(.A(G107), .ZN(new_n402));
  OR2_X1    g216(.A1(new_n382), .A2(KEYINPUT14), .ZN(new_n403));
  AOI22_X1  g217(.A1(new_n382), .A2(KEYINPUT14), .B1(G116), .B2(new_n377), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n402), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n392), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n373), .A2(new_n374), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n408), .B1(new_n203), .B2(new_n202), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n407), .B1(new_n409), .B2(new_n375), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n406), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n369), .B1(new_n401), .B2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n401), .A2(new_n411), .A3(new_n369), .ZN(new_n414));
  AOI21_X1  g228(.A(G902), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(G478), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n416), .A2(KEYINPUT15), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n415), .A2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(new_n414), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n306), .B1(new_n420), .B2(new_n412), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(new_n417), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n419), .A2(KEYINPUT96), .A3(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(KEYINPUT96), .B1(new_n419), .B2(new_n422), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT91), .ZN(new_n427));
  NAND2_X1  g241(.A1(KEYINPUT18), .A2(G131), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n269), .A2(new_n270), .A3(G214), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(new_n227), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n269), .A2(new_n270), .A3(G143), .A4(G214), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n428), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n325), .A2(G146), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n315), .A2(new_n225), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT87), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n433), .A2(new_n434), .A3(KEYINPUT87), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n432), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n430), .A2(new_n431), .A3(new_n428), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT88), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n440), .B(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n439), .A2(new_n442), .ZN(new_n443));
  XOR2_X1   g257(.A(G113), .B(G122), .Z(new_n444));
  XOR2_X1   g258(.A(KEYINPUT90), .B(G104), .Z(new_n445));
  XOR2_X1   g259(.A(new_n444), .B(new_n445), .Z(new_n446));
  NAND2_X1  g260(.A1(new_n430), .A2(new_n431), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(G131), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT17), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n430), .A2(new_n249), .A3(new_n431), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n448), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n447), .A2(KEYINPUT17), .A3(G131), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n451), .A2(new_n321), .A3(new_n326), .A4(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n443), .A2(new_n446), .A3(new_n453), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n315), .A2(KEYINPUT19), .ZN(new_n455));
  AND3_X1   g269(.A1(new_n322), .A2(new_n324), .A3(KEYINPUT19), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n225), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n343), .A2(new_n457), .A3(new_n344), .ZN(new_n458));
  AOI22_X1  g272(.A1(new_n458), .A2(KEYINPUT89), .B1(new_n448), .B2(new_n450), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT89), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n343), .A2(new_n457), .A3(new_n460), .A4(new_n344), .ZN(new_n461));
  AOI22_X1  g275(.A1(new_n459), .A2(new_n461), .B1(new_n442), .B2(new_n439), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n454), .B1(new_n462), .B2(new_n446), .ZN(new_n463));
  NOR2_X1   g277(.A1(G475), .A2(G902), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n427), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT20), .ZN(new_n466));
  AND3_X1   g280(.A1(new_n443), .A2(new_n446), .A3(new_n453), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n446), .B1(new_n443), .B2(new_n453), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n306), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  XNOR2_X1  g283(.A(KEYINPUT92), .B(G475), .ZN(new_n470));
  AOI22_X1  g284(.A1(new_n465), .A2(new_n466), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n459), .A2(new_n461), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(new_n443), .ZN(new_n473));
  INV_X1    g287(.A(new_n446), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n467), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n464), .ZN(new_n476));
  OAI21_X1  g290(.A(KEYINPUT91), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n463), .A2(new_n427), .A3(new_n464), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n477), .A2(KEYINPUT20), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n471), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(G234), .A2(G237), .ZN(new_n481));
  AND3_X1   g295(.A1(new_n481), .A2(G952), .A3(new_n270), .ZN(new_n482));
  AND3_X1   g296(.A1(new_n481), .A2(G902), .A3(G953), .ZN(new_n483));
  XNOR2_X1  g297(.A(KEYINPUT21), .B(G898), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NOR3_X1   g299(.A1(new_n426), .A2(new_n480), .A3(new_n485), .ZN(new_n486));
  OAI21_X1  g300(.A(G221), .B1(new_n368), .B2(G902), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(G469), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n489), .A2(new_n306), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n211), .A2(new_n213), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n385), .A2(G104), .A3(new_n386), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n402), .A2(G104), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(KEYINPUT3), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n402), .A2(G104), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(KEYINPUT3), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  OAI21_X1  g312(.A(G101), .B1(new_n495), .B2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(G101), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n493), .B1(new_n391), .B2(G104), .ZN(new_n501));
  OAI211_X1 g315(.A(new_n500), .B(new_n497), .C1(new_n501), .C2(KEYINPUT3), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n499), .A2(new_n502), .A3(KEYINPUT4), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT4), .ZN(new_n504));
  OAI211_X1 g318(.A(new_n504), .B(G101), .C1(new_n495), .C2(new_n498), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n503), .A2(new_n193), .A3(new_n505), .ZN(new_n506));
  AND2_X1   g320(.A1(new_n234), .A2(KEYINPUT80), .ZN(new_n507));
  OAI21_X1  g321(.A(G128), .B1(new_n234), .B2(KEYINPUT80), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n229), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n230), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n496), .B(KEYINPUT79), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n391), .A2(G104), .ZN(new_n512));
  OAI21_X1  g326(.A(G101), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n510), .A2(new_n502), .A3(new_n513), .ZN(new_n514));
  XNOR2_X1  g328(.A(KEYINPUT81), .B(KEYINPUT10), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n506), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n237), .A2(KEYINPUT10), .ZN(new_n518));
  NOR3_X1   g332(.A1(new_n495), .A2(G101), .A3(new_n498), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT79), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n496), .B(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(G104), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n387), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n500), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  OAI21_X1  g338(.A(KEYINPUT82), .B1(new_n519), .B2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT82), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n502), .A2(new_n526), .A3(new_n513), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n518), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n491), .B1(new_n517), .B2(new_n528), .ZN(new_n529));
  NOR3_X1   g343(.A1(new_n517), .A2(new_n491), .A3(new_n528), .ZN(new_n530));
  XNOR2_X1  g344(.A(G110), .B(G140), .ZN(new_n531));
  AND2_X1   g345(.A1(new_n270), .A2(G227), .ZN(new_n532));
  XNOR2_X1  g346(.A(new_n531), .B(new_n532), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  NOR3_X1   g348(.A1(new_n519), .A2(new_n524), .A3(KEYINPUT82), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n526), .B1(new_n502), .B2(new_n513), .ZN(new_n536));
  OAI211_X1 g350(.A(KEYINPUT10), .B(new_n237), .C1(new_n535), .C2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n491), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n537), .A2(new_n538), .A3(new_n506), .A4(new_n516), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n519), .A2(new_n524), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n514), .B1(new_n540), .B2(new_n237), .ZN(new_n541));
  AND3_X1   g355(.A1(new_n541), .A2(KEYINPUT12), .A3(new_n491), .ZN(new_n542));
  AOI21_X1  g356(.A(KEYINPUT12), .B1(new_n541), .B2(new_n491), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n539), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  AOI22_X1  g358(.A1(new_n529), .A2(new_n534), .B1(new_n544), .B2(new_n533), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n490), .B1(new_n545), .B2(G469), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n542), .A2(new_n543), .ZN(new_n547));
  NOR3_X1   g361(.A1(new_n547), .A2(new_n530), .A3(new_n533), .ZN(new_n548));
  INV_X1    g362(.A(new_n533), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n549), .B1(new_n529), .B2(new_n539), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n489), .B(new_n306), .C1(new_n548), .C2(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n488), .B1(new_n546), .B2(new_n551), .ZN(new_n552));
  OAI21_X1  g366(.A(G210), .B1(G237), .B2(G902), .ZN(new_n553));
  XOR2_X1   g367(.A(new_n553), .B(KEYINPUT86), .Z(new_n554));
  XNOR2_X1  g368(.A(G110), .B(G122), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT84), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n555), .B(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n503), .A2(new_n246), .A3(new_n505), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(G113), .ZN(new_n560));
  XOR2_X1   g374(.A(KEYINPUT83), .B(KEYINPUT5), .Z(new_n561));
  NOR2_X1   g375(.A1(new_n380), .A2(G119), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n563), .B1(new_n242), .B2(new_n561), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n245), .A2(new_n241), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n566), .B1(new_n525), .B2(new_n527), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n557), .B1(new_n559), .B2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n566), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n569), .B1(new_n535), .B2(new_n536), .ZN(new_n570));
  INV_X1    g384(.A(new_n557), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n570), .A2(new_n571), .A3(new_n558), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n568), .A2(KEYINPUT6), .A3(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT6), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n574), .B(new_n557), .C1(new_n559), .C2(new_n567), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n193), .A2(G125), .ZN(new_n576));
  INV_X1    g390(.A(new_n237), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n576), .B1(new_n577), .B2(G125), .ZN(new_n578));
  INV_X1    g392(.A(G224), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n579), .A2(G953), .ZN(new_n580));
  XOR2_X1   g394(.A(new_n578), .B(new_n580), .Z(new_n581));
  NAND3_X1  g395(.A1(new_n573), .A2(new_n575), .A3(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT7), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n578), .B1(new_n583), .B2(new_n580), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n580), .A2(new_n583), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n576), .B(new_n585), .C1(new_n577), .C2(G125), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n557), .B(KEYINPUT8), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT5), .ZN(new_n588));
  OAI21_X1  g402(.A(KEYINPUT85), .B1(new_n242), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(new_n563), .ZN(new_n590));
  NOR3_X1   g404(.A1(new_n242), .A2(KEYINPUT85), .A3(new_n588), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n565), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n587), .B1(new_n540), .B2(new_n592), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n569), .B1(new_n519), .B2(new_n524), .ZN(new_n594));
  AOI22_X1  g408(.A1(new_n584), .A2(new_n586), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(G902), .B1(new_n595), .B2(new_n572), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n554), .B1(new_n582), .B2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  OAI21_X1  g412(.A(G214), .B1(G237), .B2(G902), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n582), .A2(new_n554), .A3(new_n596), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  AND3_X1   g416(.A1(new_n486), .A2(new_n552), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n367), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(G101), .ZN(G3));
  INV_X1    g419(.A(G472), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n606), .B1(new_n296), .B2(new_n306), .ZN(new_n607));
  INV_X1    g421(.A(new_n297), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n267), .A2(new_n291), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(KEYINPUT28), .ZN(new_n610));
  INV_X1    g424(.A(new_n294), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n274), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n287), .A2(new_n275), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n612), .B1(new_n613), .B2(new_n265), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n608), .B1(new_n614), .B2(new_n288), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n607), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n616), .A2(new_n362), .A3(new_n552), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n413), .A2(new_n414), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n398), .A2(new_n399), .ZN(new_n619));
  INV_X1    g433(.A(new_n395), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(G134), .ZN(new_n622));
  AOI22_X1  g436(.A1(new_n622), .A2(new_n393), .B1(new_n406), .B2(new_n410), .ZN(new_n623));
  OAI21_X1  g437(.A(KEYINPUT97), .B1(new_n623), .B2(new_n369), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n618), .A2(new_n624), .A3(KEYINPUT33), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT33), .ZN(new_n626));
  OAI211_X1 g440(.A(new_n413), .B(new_n414), .C1(KEYINPUT97), .C2(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n625), .A2(G478), .A3(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n416), .A2(new_n306), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n629), .B1(new_n415), .B2(new_n416), .ZN(new_n630));
  AND2_X1   g444(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n480), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n485), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n598), .A2(new_n599), .A3(new_n600), .A4(new_n633), .ZN(new_n634));
  NOR3_X1   g448(.A1(new_n617), .A2(new_n632), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(KEYINPUT34), .B(G104), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G6));
  INV_X1    g451(.A(new_n425), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n638), .A2(new_n479), .A3(new_n471), .A4(new_n423), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n617), .A2(new_n634), .A3(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(KEYINPUT98), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT35), .B(G107), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G9));
  OR3_X1    g457(.A1(new_n352), .A2(new_n346), .A3(KEYINPUT36), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n346), .B1(new_n352), .B2(KEYINPUT36), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n644), .A2(new_n360), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(KEYINPUT99), .ZN(new_n647));
  OR2_X1    g461(.A1(new_n646), .A2(KEYINPUT99), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n359), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  AND3_X1   g463(.A1(new_n602), .A2(new_n649), .A3(new_n552), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n650), .A2(new_n486), .A3(new_n616), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(KEYINPUT100), .ZN(new_n652));
  XNOR2_X1  g466(.A(KEYINPUT37), .B(G110), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G12));
  INV_X1    g468(.A(G900), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n483), .A2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n482), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n639), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n650), .A2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n314), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(new_n190), .ZN(G30));
  NAND2_X1  g478(.A1(new_n598), .A2(new_n600), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(KEYINPUT38), .ZN(new_n666));
  INV_X1    g480(.A(new_n599), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n426), .A2(new_n480), .ZN(new_n668));
  NOR4_X1   g482(.A1(new_n666), .A2(new_n667), .A3(new_n649), .A4(new_n668), .ZN(new_n669));
  AND2_X1   g483(.A1(new_n264), .A2(new_n267), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n670), .A2(new_n289), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n308), .A2(new_n267), .A3(new_n289), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(new_n306), .ZN(new_n673));
  OAI21_X1  g487(.A(G472), .B1(new_n671), .B2(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n301), .A2(new_n674), .A3(new_n302), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n658), .B(KEYINPUT39), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n552), .A2(new_n676), .ZN(new_n677));
  OR2_X1    g491(.A1(new_n677), .A2(KEYINPUT40), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(KEYINPUT40), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n669), .A2(new_n675), .A3(new_n678), .A4(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G143), .ZN(G45));
  AND3_X1   g495(.A1(new_n480), .A2(new_n631), .A3(new_n658), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n650), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n683), .A2(new_n662), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(new_n225), .ZN(G48));
  NOR2_X1   g499(.A1(new_n548), .A2(new_n550), .ZN(new_n686));
  OAI21_X1  g500(.A(G469), .B1(new_n686), .B2(G902), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n687), .A2(new_n487), .A3(new_n551), .ZN(new_n688));
  NOR3_X1   g502(.A1(new_n688), .A2(new_n634), .A3(new_n632), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n314), .A2(new_n689), .A3(new_n362), .ZN(new_n690));
  XNOR2_X1  g504(.A(KEYINPUT41), .B(G113), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(G15));
  NOR3_X1   g506(.A1(new_n688), .A2(new_n634), .A3(new_n639), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n314), .A2(new_n693), .A3(new_n362), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G116), .ZN(G18));
  AND2_X1   g509(.A1(new_n486), .A2(new_n649), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n688), .A2(new_n601), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n696), .A2(new_n314), .A3(new_n697), .ZN(new_n698));
  XOR2_X1   g512(.A(KEYINPUT101), .B(G119), .Z(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(G21));
  OAI21_X1  g514(.A(new_n289), .B1(new_n309), .B2(new_n294), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n277), .A2(new_n288), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n297), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT102), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n702), .A2(KEYINPUT102), .A3(new_n297), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n296), .A2(new_n306), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(G472), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n707), .A2(new_n362), .A3(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(new_n688), .ZN(new_n711));
  INV_X1    g525(.A(new_n634), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT103), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n426), .A2(new_n713), .A3(new_n480), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n713), .B1(new_n426), .B2(new_n480), .ZN(new_n716));
  OAI211_X1 g530(.A(new_n711), .B(new_n712), .C1(new_n715), .C2(new_n716), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n710), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(new_n377), .ZN(G24));
  NAND2_X1  g533(.A1(new_n697), .A2(new_n682), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT104), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n607), .B1(new_n705), .B2(new_n706), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n722), .B1(new_n723), .B2(new_n649), .ZN(new_n724));
  AND3_X1   g538(.A1(new_n702), .A2(KEYINPUT102), .A3(new_n297), .ZN(new_n725));
  AOI21_X1  g539(.A(KEYINPUT102), .B1(new_n702), .B2(new_n297), .ZN(new_n726));
  OAI211_X1 g540(.A(new_n709), .B(new_n649), .C1(new_n725), .C2(new_n726), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n727), .A2(KEYINPUT104), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n721), .B1(new_n724), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(KEYINPUT105), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n727), .A2(KEYINPUT104), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n707), .A2(new_n722), .A3(new_n709), .A4(new_n649), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT105), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n733), .A2(new_n734), .A3(new_n721), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n730), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G125), .ZN(G27));
  AND3_X1   g551(.A1(new_n582), .A2(new_n554), .A3(new_n596), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n599), .B1(new_n738), .B2(new_n597), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT106), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  OAI211_X1 g555(.A(KEYINPUT106), .B(new_n599), .C1(new_n738), .C2(new_n597), .ZN(new_n742));
  AND3_X1   g556(.A1(new_n741), .A2(new_n552), .A3(new_n742), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n743), .A2(new_n314), .A3(new_n362), .A4(new_n682), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT42), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n741), .A2(new_n682), .A3(new_n552), .A4(new_n742), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n747), .A2(new_n745), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT108), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n749), .B1(new_n615), .B2(KEYINPUT32), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT32), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n298), .A2(KEYINPUT108), .A3(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT107), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n615), .A2(new_n753), .A3(KEYINPUT32), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n750), .A2(new_n752), .A3(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(new_n302), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n313), .B1(new_n756), .B2(new_n753), .ZN(new_n757));
  OAI211_X1 g571(.A(new_n748), .B(new_n362), .C1(new_n755), .C2(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n746), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G131), .ZN(G33));
  NAND4_X1  g574(.A1(new_n743), .A2(new_n314), .A3(new_n362), .A4(new_n660), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G134), .ZN(G36));
  NAND2_X1  g576(.A1(new_n741), .A2(new_n742), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n628), .A2(new_n630), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n480), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(KEYINPUT43), .ZN(new_n767));
  OAI211_X1 g581(.A(new_n767), .B(new_n649), .C1(new_n615), .C2(new_n607), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT44), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n764), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n770), .B1(new_n769), .B2(new_n768), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n545), .A2(KEYINPUT45), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(KEYINPUT109), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n545), .A2(KEYINPUT45), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n774), .A2(new_n489), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(new_n490), .ZN(new_n777));
  AOI21_X1  g591(.A(KEYINPUT46), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NOR3_X1   g592(.A1(new_n686), .A2(G469), .A3(G902), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n776), .A2(KEYINPUT46), .A3(new_n777), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n488), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n771), .A2(new_n676), .A3(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G137), .ZN(G39));
  INV_X1    g598(.A(new_n362), .ZN(new_n785));
  AND4_X1   g599(.A1(new_n662), .A2(new_n785), .A3(new_n682), .A4(new_n764), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n782), .A2(KEYINPUT47), .ZN(new_n787));
  INV_X1    g601(.A(new_n787), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n782), .A2(KEYINPUT47), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n786), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G140), .ZN(G42));
  NAND4_X1  g605(.A1(new_n362), .A2(new_n487), .A3(new_n599), .A4(new_n766), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n687), .A2(new_n551), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT49), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n792), .A2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(new_n675), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n793), .A2(new_n794), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n796), .A2(new_n797), .A3(new_n666), .A4(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n767), .A2(new_n482), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n800), .A2(new_n710), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n801), .A2(new_n667), .A3(new_n666), .A4(new_n711), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n802), .A2(KEYINPUT50), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n802), .A2(KEYINPUT50), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n763), .A2(new_n688), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n805), .A2(new_n482), .A3(new_n767), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n806), .B1(new_n732), .B2(new_n731), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n803), .A2(new_n804), .A3(new_n807), .ZN(new_n808));
  AND4_X1   g622(.A1(new_n362), .A2(new_n797), .A3(new_n482), .A4(new_n805), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n809), .A2(new_n479), .A3(new_n471), .A4(new_n765), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n810), .A2(KEYINPUT51), .ZN(new_n811));
  INV_X1    g625(.A(new_n789), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n793), .A2(new_n488), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n812), .A2(KEYINPUT115), .A3(new_n787), .A4(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n814), .A2(new_n764), .A3(new_n801), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n788), .A2(new_n789), .ZN(new_n816));
  AOI21_X1  g630(.A(KEYINPUT115), .B1(new_n816), .B2(new_n813), .ZN(new_n817));
  OAI211_X1 g631(.A(new_n808), .B(new_n811), .C1(new_n815), .C2(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n809), .A2(new_n480), .A3(new_n631), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n801), .A2(new_n697), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n819), .A2(G952), .A3(new_n270), .A4(new_n820), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n362), .B1(new_n755), .B2(new_n757), .ZN(new_n822));
  OR2_X1    g636(.A1(new_n822), .A2(new_n806), .ZN(new_n823));
  INV_X1    g637(.A(new_n823), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n824), .A2(KEYINPUT116), .A3(KEYINPUT48), .ZN(new_n825));
  XOR2_X1   g639(.A(KEYINPUT116), .B(KEYINPUT48), .Z(new_n826));
  AOI211_X1 g640(.A(new_n821), .B(new_n825), .C1(new_n824), .C2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n801), .A2(new_n764), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n828), .B1(new_n816), .B2(new_n813), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n808), .A2(new_n810), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n818), .B(new_n827), .C1(KEYINPUT51), .C2(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n419), .A2(new_n422), .ZN(new_n833));
  INV_X1    g647(.A(new_n833), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n632), .B1(new_n480), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(new_n712), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n651), .B1(new_n617), .B2(new_n836), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n837), .B1(new_n367), .B2(new_n603), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n480), .A2(new_n833), .A3(new_n659), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n741), .A2(new_n742), .A3(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT110), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n649), .A2(new_n552), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n842), .A2(new_n314), .A3(new_n843), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n840), .A2(new_n841), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n761), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n747), .B1(new_n731), .B2(new_n732), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n838), .A2(new_n848), .A3(KEYINPUT53), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n694), .B1(new_n710), .B2(new_n717), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n698), .A2(new_n690), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n852), .A2(new_n759), .A3(KEYINPUT113), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT113), .B1(new_n852), .B2(new_n759), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n849), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n662), .B1(new_n661), .B2(new_n683), .ZN(new_n856));
  INV_X1    g670(.A(new_n716), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n601), .B1(new_n857), .B2(new_n714), .ZN(new_n858));
  INV_X1    g672(.A(new_n552), .ZN(new_n859));
  XOR2_X1   g673(.A(new_n658), .B(KEYINPUT111), .Z(new_n860));
  NOR3_X1   g674(.A1(new_n859), .A2(new_n649), .A3(new_n860), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n858), .A2(new_n861), .A3(new_n675), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n856), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n734), .B1(new_n733), .B2(new_n721), .ZN(new_n864));
  AOI211_X1 g678(.A(KEYINPUT105), .B(new_n720), .C1(new_n731), .C2(new_n732), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n863), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT52), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OAI211_X1 g682(.A(KEYINPUT52), .B(new_n863), .C1(new_n864), .C2(new_n865), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n855), .A2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT54), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n838), .A2(new_n848), .A3(new_n759), .A4(new_n852), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n873), .B1(new_n868), .B2(new_n869), .ZN(new_n874));
  XNOR2_X1  g688(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  OAI211_X1 g690(.A(new_n871), .B(new_n872), .C1(new_n874), .C2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(new_n873), .ZN(new_n878));
  AOI21_X1  g692(.A(KEYINPUT52), .B1(new_n736), .B2(new_n863), .ZN(new_n879));
  INV_X1    g693(.A(new_n869), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n878), .B(new_n875), .C1(new_n879), .C2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT53), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n881), .B(KEYINPUT54), .C1(new_n882), .C2(new_n874), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n877), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(KEYINPUT114), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT114), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n877), .A2(new_n883), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n832), .B1(new_n885), .B2(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(G952), .A2(G953), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n799), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT117), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  OAI211_X1 g706(.A(KEYINPUT117), .B(new_n799), .C1(new_n888), .C2(new_n889), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(G75));
  NOR2_X1   g708(.A1(new_n270), .A2(G952), .ZN(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n871), .B1(new_n874), .B2(new_n876), .ZN(new_n897));
  INV_X1    g711(.A(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n898), .A2(new_n306), .ZN(new_n899));
  AOI21_X1  g713(.A(KEYINPUT56), .B1(new_n899), .B2(new_n554), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n573), .A2(new_n575), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(new_n581), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n902), .B(KEYINPUT55), .Z(new_n903));
  INV_X1    g717(.A(new_n903), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n896), .B1(new_n900), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n905), .B1(new_n900), .B2(new_n904), .ZN(G51));
  NAND2_X1  g720(.A1(new_n897), .A2(KEYINPUT54), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(new_n877), .ZN(new_n908));
  XNOR2_X1  g722(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(new_n490), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n911), .B1(new_n550), .B2(new_n548), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n899), .A2(new_n773), .A3(new_n775), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n895), .B1(new_n912), .B2(new_n913), .ZN(G54));
  NAND2_X1  g728(.A1(KEYINPUT58), .A2(G475), .ZN(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n897), .A2(G902), .A3(new_n916), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n917), .A2(new_n475), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n918), .A2(new_n895), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n917), .A2(KEYINPUT119), .A3(new_n475), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n917), .A2(new_n475), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT119), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n919), .A2(new_n920), .A3(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT120), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n919), .A2(KEYINPUT120), .A3(new_n920), .A4(new_n923), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(G60));
  NAND2_X1  g742(.A1(new_n625), .A2(new_n627), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n929), .B(KEYINPUT121), .Z(new_n930));
  XNOR2_X1  g744(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(new_n629), .Z(new_n932));
  AOI211_X1 g746(.A(new_n930), .B(new_n932), .C1(new_n907), .C2(new_n877), .ZN(new_n933));
  INV_X1    g747(.A(new_n932), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n885), .A2(new_n887), .A3(new_n934), .ZN(new_n935));
  AOI211_X1 g749(.A(new_n895), .B(new_n933), .C1(new_n930), .C2(new_n935), .ZN(G63));
  INV_X1    g750(.A(KEYINPUT61), .ZN(new_n937));
  NAND2_X1  g751(.A1(G217), .A2(G902), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT60), .ZN(new_n939));
  OAI21_X1  g753(.A(KEYINPUT123), .B1(new_n898), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n351), .A2(new_n353), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT123), .ZN(new_n942));
  INV_X1    g756(.A(new_n939), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n897), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n940), .A2(new_n941), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(new_n896), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n644), .A2(new_n645), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n947), .B1(new_n940), .B2(new_n944), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n937), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(new_n948), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n950), .A2(KEYINPUT61), .A3(new_n896), .A4(new_n945), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n949), .A2(new_n951), .ZN(G66));
  OAI21_X1  g766(.A(G953), .B1(new_n484), .B2(new_n579), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n838), .A2(new_n852), .ZN(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n953), .B1(new_n955), .B2(G953), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n901), .B1(G898), .B2(new_n270), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n956), .B(new_n957), .ZN(G69));
  INV_X1    g772(.A(KEYINPUT124), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n856), .B1(new_n730), .B2(new_n735), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(new_n680), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(KEYINPUT62), .ZN(new_n962));
  INV_X1    g776(.A(new_n677), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n367), .A2(new_n963), .A3(new_n764), .A4(new_n835), .ZN(new_n964));
  AND4_X1   g778(.A1(new_n783), .A2(new_n962), .A3(new_n790), .A4(new_n964), .ZN(new_n965));
  OR2_X1    g779(.A1(new_n961), .A2(KEYINPUT62), .ZN(new_n966));
  AOI21_X1  g780(.A(G953), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n240), .B1(new_n262), .B2(new_n263), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n455), .A2(new_n456), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n968), .B(new_n969), .Z(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n959), .B1(new_n967), .B2(new_n971), .ZN(new_n972));
  AND2_X1   g786(.A1(new_n790), .A2(new_n783), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n966), .A2(new_n973), .A3(new_n962), .A4(new_n964), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n974), .A2(new_n270), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n975), .A2(KEYINPUT124), .A3(new_n970), .ZN(new_n976));
  AND2_X1   g790(.A1(new_n972), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n970), .B1(G900), .B2(G953), .ZN(new_n978));
  INV_X1    g792(.A(new_n822), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n782), .A2(new_n676), .A3(new_n979), .A4(new_n858), .ZN(new_n980));
  AND3_X1   g794(.A1(new_n980), .A2(new_n759), .A3(new_n761), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n973), .A2(new_n960), .A3(new_n981), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n978), .B1(new_n982), .B2(G953), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT125), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n270), .B1(G227), .B2(G900), .ZN(new_n985));
  INV_X1    g799(.A(new_n985), .ZN(new_n986));
  OAI211_X1 g800(.A(new_n977), .B(new_n983), .C1(new_n984), .C2(new_n986), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n972), .A2(new_n984), .A3(new_n976), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n972), .A2(new_n976), .A3(new_n983), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n988), .A2(new_n989), .A3(new_n985), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n987), .A2(new_n990), .ZN(G72));
  XNOR2_X1  g805(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n992));
  NAND2_X1  g806(.A1(G472), .A2(G902), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n992), .B(new_n993), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n994), .B1(new_n982), .B2(new_n954), .ZN(new_n995));
  XOR2_X1   g809(.A(new_n303), .B(KEYINPUT127), .Z(new_n996));
  AOI21_X1  g810(.A(new_n895), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n881), .B1(new_n882), .B2(new_n874), .ZN(new_n998));
  INV_X1    g812(.A(new_n671), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n999), .A2(new_n303), .A3(new_n994), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n997), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n994), .B1(new_n974), .B2(new_n954), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n1001), .B1(new_n671), .B2(new_n1002), .ZN(G57));
endmodule


