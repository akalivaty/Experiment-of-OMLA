//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 0 0 1 0 0 0 1 0 1 1 0 0 1 1 1 1 0 0 0 1 1 1 1 0 1 1 1 0 0 0 1 1 1 1 0 1 0 0 0 1 1 0 0 0 0 0 1 1 0 0 0 0 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:54 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n564, new_n566, new_n567, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n616,
    new_n619, new_n621, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1186, new_n1187, new_n1188, new_n1190, new_n1191;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(KEYINPUT64), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  OAI21_X1  g038(.A(new_n462), .B1(new_n463), .B2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n465), .A2(KEYINPUT64), .A3(G2104), .ZN(new_n466));
  INV_X1    g041(.A(G137), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n469));
  NAND4_X1  g044(.A1(new_n464), .A2(new_n466), .A3(new_n468), .A4(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n463), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G101), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT65), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n470), .A2(KEYINPUT65), .A3(new_n472), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n465), .A2(G2104), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n469), .A2(new_n478), .A3(G125), .ZN(new_n479));
  NAND2_X1  g054(.A1(G113), .A2(G2104), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n477), .B1(G2105), .B2(new_n481), .ZN(G160));
  AND3_X1   g057(.A1(new_n464), .A2(new_n469), .A3(new_n466), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(G124), .ZN(new_n485));
  INV_X1    g060(.A(G2105), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n486), .A2(G112), .ZN(new_n487));
  OAI21_X1  g062(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n488));
  OAI22_X1  g063(.A1(new_n484), .A2(new_n485), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  AND2_X1   g064(.A1(new_n483), .A2(new_n486), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n489), .B1(G136), .B2(new_n490), .ZN(G162));
  INV_X1    g066(.A(KEYINPUT67), .ZN(new_n492));
  XNOR2_X1  g067(.A(KEYINPUT3), .B(G2104), .ZN(new_n493));
  INV_X1    g068(.A(G138), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n494), .A2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT66), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT66), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n499));
  AND3_X1   g074(.A1(new_n495), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n464), .A2(new_n466), .A3(new_n495), .A4(new_n469), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n493), .A2(new_n500), .B1(new_n501), .B2(KEYINPUT4), .ZN(new_n502));
  AND2_X1   g077(.A1(G126), .A2(G2105), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n464), .A2(new_n466), .A3(new_n469), .A4(new_n503), .ZN(new_n504));
  OR2_X1    g079(.A1(G102), .A2(G2105), .ZN(new_n505));
  OAI211_X1 g080(.A(new_n505), .B(G2104), .C1(G114), .C2(new_n486), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n492), .B1(new_n502), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n501), .A2(KEYINPUT4), .ZN(new_n509));
  NAND4_X1  g084(.A1(new_n493), .A2(new_n495), .A3(new_n497), .A4(new_n499), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n507), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n511), .A2(KEYINPUT67), .A3(new_n512), .ZN(new_n513));
  AND2_X1   g088(.A1(new_n508), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(G164));
  XNOR2_X1  g090(.A(KEYINPUT5), .B(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G62), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT68), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n517), .A2(new_n518), .B1(G75), .B2(G543), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n516), .A2(KEYINPUT68), .A3(G62), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G651), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT69), .ZN(new_n523));
  XNOR2_X1  g098(.A(KEYINPUT6), .B(G651), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n516), .A2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(G88), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n524), .A2(G543), .ZN(new_n527));
  INV_X1    g102(.A(G50), .ZN(new_n528));
  OAI22_X1  g103(.A1(new_n525), .A2(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n522), .A2(new_n523), .A3(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(G651), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n532), .B1(new_n519), .B2(new_n520), .ZN(new_n533));
  OAI21_X1  g108(.A(KEYINPUT69), .B1(new_n533), .B2(new_n529), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n531), .A2(new_n534), .ZN(G166));
  OR2_X1    g110(.A1(new_n527), .A2(KEYINPUT70), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n527), .A2(KEYINPUT70), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  AND2_X1   g113(.A1(new_n538), .A2(G51), .ZN(new_n539));
  NAND3_X1  g114(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT7), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n516), .A2(G63), .A3(G651), .ZN(new_n542));
  INV_X1    g117(.A(G89), .ZN(new_n543));
  OAI211_X1 g118(.A(new_n541), .B(new_n542), .C1(new_n525), .C2(new_n543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n539), .A2(new_n544), .ZN(G168));
  XOR2_X1   g120(.A(KEYINPUT71), .B(G52), .Z(new_n546));
  AOI21_X1  g121(.A(new_n546), .B1(new_n536), .B2(new_n537), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n516), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n548));
  INV_X1    g123(.A(G90), .ZN(new_n549));
  OAI22_X1  g124(.A1(new_n548), .A2(new_n532), .B1(new_n525), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n547), .A2(new_n550), .ZN(G171));
  INV_X1    g126(.A(new_n525), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n538), .A2(G43), .B1(G81), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(G68), .A2(G543), .ZN(new_n554));
  AND2_X1   g129(.A1(KEYINPUT5), .A2(G543), .ZN(new_n555));
  NOR2_X1   g130(.A1(KEYINPUT5), .A2(G543), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(G56), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n554), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  AOI21_X1  g134(.A(new_n532), .B1(new_n559), .B2(KEYINPUT72), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n560), .B1(KEYINPUT72), .B2(new_n559), .ZN(new_n561));
  AND2_X1   g136(.A1(new_n553), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G860), .ZN(G153));
  NAND4_X1  g138(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n564));
  XOR2_X1   g139(.A(new_n564), .B(KEYINPUT73), .Z(G176));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND4_X1  g142(.A1(G319), .A2(G483), .A3(G661), .A4(new_n567), .ZN(G188));
  AND2_X1   g143(.A1(new_n524), .A2(G543), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G53), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT9), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n570), .B(new_n571), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n516), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n573));
  INV_X1    g148(.A(G91), .ZN(new_n574));
  OAI22_X1  g149(.A1(new_n573), .A2(new_n532), .B1(new_n525), .B2(new_n574), .ZN(new_n575));
  OR2_X1    g150(.A1(new_n572), .A2(new_n575), .ZN(G299));
  INV_X1    g151(.A(G171), .ZN(G301));
  OR2_X1    g152(.A1(new_n539), .A2(new_n544), .ZN(G286));
  AND2_X1   g153(.A1(new_n531), .A2(new_n534), .ZN(G303));
  INV_X1    g154(.A(G74), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n532), .B1(new_n557), .B2(new_n580), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n581), .B1(G49), .B2(new_n569), .ZN(new_n582));
  AOI21_X1  g157(.A(KEYINPUT74), .B1(new_n552), .B2(G87), .ZN(new_n583));
  AND4_X1   g158(.A1(KEYINPUT74), .A2(new_n516), .A3(new_n524), .A4(G87), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n582), .B1(new_n583), .B2(new_n584), .ZN(G288));
  INV_X1    g160(.A(G61), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n557), .A2(new_n586), .ZN(new_n587));
  AND2_X1   g162(.A1(G73), .A2(G543), .ZN(new_n588));
  OAI21_X1  g163(.A(G651), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n516), .A2(new_n524), .A3(G86), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n524), .A2(G48), .A3(G543), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(G305));
  NAND2_X1  g167(.A1(new_n538), .A2(G47), .ZN(new_n593));
  NAND2_X1  g168(.A1(G72), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G60), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n557), .B2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT75), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n532), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n598), .B1(new_n597), .B2(new_n596), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n552), .A2(G85), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n593), .A2(new_n599), .A3(new_n600), .ZN(G290));
  NAND2_X1  g176(.A1(G301), .A2(G868), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n552), .A2(G92), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT10), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n603), .B(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n538), .A2(G54), .ZN(new_n606));
  NAND2_X1  g181(.A1(G79), .A2(G543), .ZN(new_n607));
  XNOR2_X1  g182(.A(KEYINPUT76), .B(G66), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n557), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(G651), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n605), .A2(new_n606), .A3(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n602), .B1(new_n612), .B2(G868), .ZN(G284));
  OAI21_X1  g188(.A(new_n602), .B1(new_n612), .B2(G868), .ZN(G321));
  INV_X1    g189(.A(G868), .ZN(new_n615));
  NAND2_X1  g190(.A1(G299), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(new_n615), .B2(G168), .ZN(G297));
  OAI21_X1  g192(.A(new_n616), .B1(new_n615), .B2(G168), .ZN(G280));
  INV_X1    g193(.A(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n612), .B1(new_n619), .B2(G860), .ZN(G148));
  OAI21_X1  g195(.A(KEYINPUT77), .B1(new_n562), .B2(G868), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n611), .A2(G559), .ZN(new_n622));
  NOR2_X1   g197(.A1(new_n622), .A2(new_n615), .ZN(new_n623));
  MUX2_X1   g198(.A(new_n621), .B(KEYINPUT77), .S(new_n623), .Z(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g200(.A1(new_n493), .A2(new_n471), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(KEYINPUT12), .Z(new_n627));
  INV_X1    g202(.A(G2100), .ZN(new_n628));
  OAI22_X1  g203(.A1(new_n627), .A2(KEYINPUT13), .B1(KEYINPUT78), .B2(new_n628), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n629), .B1(KEYINPUT13), .B2(new_n627), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n628), .A2(KEYINPUT78), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  INV_X1    g207(.A(G123), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n486), .A2(G111), .ZN(new_n634));
  OAI21_X1  g209(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n635));
  OAI22_X1  g210(.A1(new_n484), .A2(new_n633), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n636), .B1(G135), .B2(new_n490), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2096), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n632), .A2(new_n638), .ZN(G156));
  INV_X1    g214(.A(KEYINPUT14), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2427), .B(G2438), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2430), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT15), .B(G2435), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n640), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n644), .B1(new_n643), .B2(new_n642), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2451), .B(G2454), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT16), .ZN(new_n647));
  XOR2_X1   g222(.A(G1341), .B(G1348), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n645), .B(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(G2443), .B(G2446), .Z(new_n651));
  OAI21_X1  g226(.A(G14), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n652), .B1(new_n651), .B2(new_n650), .ZN(G401));
  XNOR2_X1  g228(.A(G2072), .B(G2078), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(KEYINPUT17), .Z(new_n655));
  XNOR2_X1  g230(.A(G2067), .B(G2678), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2084), .B(G2090), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT79), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n654), .A2(new_n656), .ZN(new_n661));
  NOR3_X1   g236(.A1(new_n658), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT80), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n660), .A2(new_n656), .A3(new_n654), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(KEYINPUT18), .Z(new_n665));
  NAND3_X1  g240(.A1(new_n655), .A2(new_n660), .A3(new_n657), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n663), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G2096), .B(G2100), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(G227));
  XOR2_X1   g244(.A(G1956), .B(G2474), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT81), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1961), .B(G1966), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1971), .B(G1976), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT19), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(KEYINPUT20), .Z(new_n678));
  NOR2_X1   g253(.A1(new_n671), .A2(new_n673), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n680), .A2(new_n676), .A3(new_n674), .ZN(new_n681));
  OAI211_X1 g256(.A(new_n678), .B(new_n681), .C1(new_n676), .C2(new_n680), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G1991), .B(G1996), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT82), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n684), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1981), .B(G1986), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n687), .A2(new_n689), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n690), .A2(new_n691), .ZN(G229));
  XOR2_X1   g267(.A(KEYINPUT83), .B(G29), .Z(new_n693));
  INV_X1    g268(.A(KEYINPUT24), .ZN(new_n694));
  OR2_X1    g269(.A1(new_n694), .A2(G34), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n694), .A2(G34), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n693), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(G160), .ZN(new_n698));
  INV_X1    g273(.A(G29), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n697), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(G2084), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n702), .B(KEYINPUT90), .Z(new_n703));
  INV_X1    g278(.A(G16), .ZN(new_n704));
  NOR2_X1   g279(.A1(G168), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(new_n704), .B2(G21), .ZN(new_n706));
  INV_X1    g281(.A(G1966), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT31), .B(G11), .ZN(new_n709));
  INV_X1    g284(.A(G28), .ZN(new_n710));
  AOI21_X1  g285(.A(G29), .B1(new_n710), .B2(KEYINPUT30), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(KEYINPUT92), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(KEYINPUT30), .B2(new_n710), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n711), .A2(KEYINPUT92), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n709), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(new_n693), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n715), .B1(new_n637), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n708), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n704), .A2(G5), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(G171), .B2(new_n704), .ZN(new_n720));
  OAI22_X1  g295(.A1(new_n706), .A2(new_n707), .B1(G1961), .B2(new_n720), .ZN(new_n721));
  AND2_X1   g296(.A1(new_n720), .A2(G1961), .ZN(new_n722));
  NOR3_X1   g297(.A1(new_n718), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n699), .A2(G32), .ZN(new_n724));
  AND2_X1   g299(.A1(new_n490), .A2(G141), .ZN(new_n725));
  NAND3_X1  g300(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT26), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n726), .A2(new_n727), .ZN(new_n729));
  AOI22_X1  g304(.A1(new_n728), .A2(new_n729), .B1(G105), .B2(new_n471), .ZN(new_n730));
  INV_X1    g305(.A(G129), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n730), .B1(new_n484), .B2(new_n731), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n725), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT91), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n724), .B1(new_n734), .B2(new_n699), .ZN(new_n735));
  XNOR2_X1  g310(.A(KEYINPUT27), .B(G1996), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n699), .A2(G33), .ZN(new_n738));
  AOI22_X1  g313(.A1(new_n493), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n739), .A2(new_n486), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT89), .ZN(new_n741));
  AND2_X1   g316(.A1(new_n490), .A2(G139), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n486), .A2(G103), .A3(G2104), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT25), .ZN(new_n744));
  NOR3_X1   g319(.A1(new_n741), .A2(new_n742), .A3(new_n744), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n738), .B1(new_n745), .B2(new_n699), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(G2072), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(new_n701), .B2(new_n700), .ZN(new_n748));
  AND4_X1   g323(.A1(new_n703), .A2(new_n723), .A3(new_n737), .A4(new_n748), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n716), .A2(G35), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(G162), .B2(new_n716), .ZN(new_n751));
  XNOR2_X1  g326(.A(KEYINPUT94), .B(KEYINPUT29), .ZN(new_n752));
  AND2_X1   g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n751), .A2(new_n752), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n755), .A2(G2090), .ZN(new_n756));
  XNOR2_X1  g331(.A(KEYINPUT95), .B(KEYINPUT23), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT96), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n704), .A2(G20), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n758), .B(new_n759), .Z(new_n760));
  NOR2_X1   g335(.A1(new_n572), .A2(new_n575), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n760), .B1(new_n761), .B2(new_n704), .ZN(new_n762));
  INV_X1    g337(.A(G1956), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  AND3_X1   g339(.A1(new_n756), .A2(KEYINPUT97), .A3(new_n764), .ZN(new_n765));
  AOI21_X1  g340(.A(KEYINPUT97), .B1(new_n756), .B2(new_n764), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n693), .A2(G27), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT93), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G164), .B2(new_n693), .ZN(new_n769));
  INV_X1    g344(.A(G2078), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(new_n755), .B2(G2090), .ZN(new_n772));
  NOR3_X1   g347(.A1(new_n765), .A2(new_n766), .A3(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(G128), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n486), .A2(G116), .ZN(new_n775));
  OAI21_X1  g350(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n776));
  OAI22_X1  g351(.A1(new_n484), .A2(new_n774), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(G140), .B2(new_n490), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n778), .A2(new_n699), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT86), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n693), .A2(G26), .ZN(new_n781));
  XOR2_X1   g356(.A(KEYINPUT87), .B(KEYINPUT28), .Z(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n780), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(G2067), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n704), .A2(G19), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(new_n562), .B2(new_n704), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(G1341), .Z(new_n788));
  NAND2_X1  g363(.A1(new_n704), .A2(G4), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(new_n612), .B2(new_n704), .ZN(new_n790));
  INV_X1    g365(.A(G1348), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n788), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n785), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n794), .A2(KEYINPUT88), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT88), .ZN(new_n796));
  NOR3_X1   g371(.A1(new_n785), .A2(new_n793), .A3(new_n796), .ZN(new_n797));
  OAI211_X1 g372(.A(new_n749), .B(new_n773), .C1(new_n795), .C2(new_n797), .ZN(new_n798));
  MUX2_X1   g373(.A(G6), .B(G305), .S(G16), .Z(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT32), .ZN(new_n800));
  INV_X1    g375(.A(G1981), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n704), .A2(G22), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G166), .B2(new_n704), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n804), .A2(G1971), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n804), .A2(G1971), .ZN(new_n806));
  MUX2_X1   g381(.A(G23), .B(G288), .S(G16), .Z(new_n807));
  XNOR2_X1  g382(.A(KEYINPUT33), .B(G1976), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n802), .A2(new_n805), .A3(new_n806), .A4(new_n809), .ZN(new_n810));
  OR2_X1    g385(.A1(new_n810), .A2(KEYINPUT34), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n810), .A2(KEYINPUT34), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n693), .A2(G25), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT84), .ZN(new_n814));
  OAI21_X1  g389(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n815));
  INV_X1    g390(.A(G107), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n815), .B1(new_n816), .B2(G2105), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT85), .ZN(new_n818));
  INV_X1    g393(.A(G119), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n818), .B1(new_n484), .B2(new_n819), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n820), .B1(G131), .B2(new_n490), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n814), .B1(new_n821), .B2(new_n693), .ZN(new_n822));
  XOR2_X1   g397(.A(KEYINPUT35), .B(G1991), .Z(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NOR2_X1   g399(.A1(G16), .A2(G24), .ZN(new_n825));
  INV_X1    g400(.A(G290), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n825), .B1(new_n826), .B2(G16), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(G1986), .Z(new_n828));
  NAND4_X1  g403(.A1(new_n811), .A2(new_n812), .A3(new_n824), .A4(new_n828), .ZN(new_n829));
  OR2_X1    g404(.A1(new_n829), .A2(KEYINPUT36), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(KEYINPUT36), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n798), .B1(new_n830), .B2(new_n831), .ZN(G311));
  XNOR2_X1  g407(.A(G311), .B(KEYINPUT98), .ZN(G150));
  AOI22_X1  g408(.A1(new_n516), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n834));
  INV_X1    g409(.A(G93), .ZN(new_n835));
  OAI22_X1  g410(.A1(new_n834), .A2(new_n532), .B1(new_n525), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n836), .B1(new_n538), .B2(G55), .ZN(new_n837));
  INV_X1    g412(.A(G860), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT37), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n837), .A2(KEYINPUT99), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n553), .A2(new_n561), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n837), .A2(KEYINPUT99), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n562), .A2(KEYINPUT99), .A3(new_n837), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT38), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n612), .A2(G559), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n847), .B(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT39), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n851), .B(KEYINPUT100), .Z(new_n852));
  OAI21_X1  g427(.A(new_n838), .B1(new_n849), .B2(new_n850), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n840), .B1(new_n852), .B2(new_n853), .ZN(G145));
  NAND3_X1  g429(.A1(new_n504), .A2(new_n506), .A3(KEYINPUT102), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  AOI21_X1  g431(.A(KEYINPUT102), .B1(new_n504), .B2(new_n506), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n511), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n778), .B(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n490), .A2(G142), .ZN(new_n860));
  INV_X1    g435(.A(G130), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n486), .A2(G118), .ZN(new_n862));
  OAI21_X1  g437(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n863));
  OAI221_X1 g438(.A(new_n860), .B1(new_n861), .B2(new_n484), .C1(new_n862), .C2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n859), .B(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n821), .B(new_n627), .ZN(new_n866));
  OR2_X1    g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n865), .A2(new_n866), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n734), .ZN(new_n870));
  AND2_X1   g445(.A1(new_n870), .A2(new_n745), .ZN(new_n871));
  INV_X1    g446(.A(new_n733), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n745), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n869), .A2(new_n874), .ZN(new_n875));
  OAI211_X1 g450(.A(new_n867), .B(new_n868), .C1(new_n871), .C2(new_n873), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n637), .B(KEYINPUT101), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(new_n698), .ZN(new_n879));
  XOR2_X1   g454(.A(new_n879), .B(G162), .Z(new_n880));
  AOI21_X1  g455(.A(G37), .B1(new_n877), .B2(new_n880), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n877), .A2(new_n880), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n882), .A2(KEYINPUT103), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT103), .ZN(new_n884));
  NOR3_X1   g459(.A1(new_n877), .A2(new_n880), .A3(new_n884), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n881), .B1(new_n883), .B2(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g462(.A1(new_n611), .A2(new_n761), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT104), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n612), .A2(G299), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n611), .A2(new_n761), .A3(KEYINPUT104), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  OR2_X1    g468(.A1(new_n893), .A2(KEYINPUT41), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(KEYINPUT41), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n846), .B(new_n622), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n898), .B1(new_n893), .B2(new_n897), .ZN(new_n899));
  NAND2_X1  g474(.A1(G303), .A2(G290), .ZN(new_n900));
  NAND2_X1  g475(.A1(G166), .A2(new_n826), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(G288), .B(G305), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n902), .B(new_n903), .ZN(new_n904));
  AND2_X1   g479(.A1(new_n904), .A2(KEYINPUT42), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n904), .A2(KEYINPUT42), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n899), .A2(new_n907), .ZN(new_n908));
  OAI221_X1 g483(.A(new_n898), .B1(new_n893), .B2(new_n897), .C1(new_n905), .C2(new_n906), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n908), .A2(new_n909), .A3(G868), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT105), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n911), .B1(new_n837), .B2(G868), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n908), .A2(new_n909), .A3(KEYINPUT105), .A4(G868), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n916), .B(KEYINPUT106), .ZN(G295));
  INV_X1    g492(.A(new_n916), .ZN(G331));
  INV_X1    g493(.A(KEYINPUT44), .ZN(new_n919));
  NAND2_X1  g494(.A1(G286), .A2(G301), .ZN(new_n920));
  NAND2_X1  g495(.A1(G168), .A2(G171), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n846), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT107), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n844), .A2(new_n845), .A3(new_n920), .A4(new_n921), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n846), .A2(new_n922), .A3(KEYINPUT107), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n894), .A2(new_n926), .A3(new_n895), .A4(new_n927), .ZN(new_n928));
  AND2_X1   g503(.A1(new_n923), .A2(new_n925), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(new_n893), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n903), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n902), .B(new_n932), .ZN(new_n933));
  OAI21_X1  g508(.A(KEYINPUT109), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT109), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n928), .A2(new_n935), .A3(new_n904), .A4(new_n930), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n926), .A2(new_n927), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(new_n893), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n939), .B1(new_n896), .B2(new_n929), .ZN(new_n940));
  AOI21_X1  g515(.A(G37), .B1(new_n940), .B2(new_n933), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n937), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(KEYINPUT43), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT43), .ZN(new_n944));
  AOI21_X1  g519(.A(G37), .B1(new_n931), .B2(new_n933), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n945), .A2(KEYINPUT108), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT108), .ZN(new_n947));
  AOI211_X1 g522(.A(new_n947), .B(G37), .C1(new_n931), .C2(new_n933), .ZN(new_n948));
  OAI211_X1 g523(.A(new_n944), .B(new_n937), .C1(new_n946), .C2(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n919), .B1(new_n943), .B2(new_n949), .ZN(new_n950));
  AND3_X1   g525(.A1(new_n937), .A2(new_n944), .A3(new_n941), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n937), .B1(new_n946), .B2(new_n948), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n951), .B1(KEYINPUT43), .B2(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n950), .B1(new_n919), .B2(new_n953), .ZN(G397));
  INV_X1    g529(.A(G40), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n955), .B1(new_n481), .B2(G2105), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n475), .A2(new_n956), .A3(new_n476), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT111), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n475), .A2(new_n956), .A3(KEYINPUT111), .A4(new_n476), .ZN(new_n960));
  AND2_X1   g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT102), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n507), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(new_n855), .ZN(new_n964));
  AOI21_X1  g539(.A(G1384), .B1(new_n964), .B2(new_n511), .ZN(new_n965));
  XNOR2_X1  g540(.A(KEYINPUT110), .B(KEYINPUT45), .ZN(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n961), .A2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  XOR2_X1   g545(.A(new_n821), .B(new_n823), .Z(new_n971));
  XNOR2_X1  g546(.A(new_n971), .B(KEYINPUT112), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n778), .B(G2067), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n872), .A2(G1996), .ZN(new_n974));
  OAI211_X1 g549(.A(new_n973), .B(new_n974), .C1(new_n870), .C2(G1996), .ZN(new_n975));
  OR2_X1    g550(.A1(new_n972), .A2(new_n975), .ZN(new_n976));
  XNOR2_X1  g551(.A(G290), .B(G1986), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n970), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n959), .A2(new_n960), .ZN(new_n979));
  INV_X1    g554(.A(G1384), .ZN(new_n980));
  AOI21_X1  g555(.A(KEYINPUT45), .B1(new_n858), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT115), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT45), .ZN(new_n983));
  AOI22_X1  g558(.A1(new_n963), .A2(new_n855), .B1(new_n509), .B2(new_n510), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n983), .B1(new_n984), .B2(G1384), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT115), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n985), .A2(new_n986), .A3(new_n959), .A4(new_n960), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n514), .A2(new_n980), .A3(new_n967), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT53), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n989), .A2(G2078), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n982), .A2(new_n987), .A3(new_n988), .A4(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(G1961), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n508), .A2(new_n980), .A3(new_n513), .ZN(new_n993));
  AND2_X1   g568(.A1(new_n993), .A2(KEYINPUT50), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n858), .A2(new_n980), .ZN(new_n995));
  OAI211_X1 g570(.A(new_n959), .B(new_n960), .C1(new_n995), .C2(KEYINPUT50), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n992), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n991), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n993), .A2(new_n966), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n858), .A2(KEYINPUT45), .A3(new_n980), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n961), .A2(new_n999), .A3(new_n770), .A4(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(new_n989), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(KEYINPUT121), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT121), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1001), .A2(new_n1004), .A3(new_n989), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n998), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(KEYINPUT122), .B1(new_n1006), .B2(G301), .ZN(new_n1007));
  AND3_X1   g582(.A1(new_n1001), .A2(new_n1004), .A3(new_n989), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1004), .B1(new_n1001), .B2(new_n989), .ZN(new_n1009));
  OAI211_X1 g584(.A(new_n997), .B(new_n991), .C1(new_n1008), .C2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT122), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1010), .A2(new_n1011), .A3(G171), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n770), .A2(KEYINPUT53), .ZN(new_n1013));
  NOR3_X1   g588(.A1(new_n968), .A2(new_n957), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n993), .A2(KEYINPUT50), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT50), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n965), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n961), .A2(new_n1015), .A3(new_n1017), .ZN(new_n1018));
  AOI22_X1  g593(.A1(new_n1000), .A2(new_n1014), .B1(new_n1018), .B2(new_n992), .ZN(new_n1019));
  OAI211_X1 g594(.A(new_n1019), .B(G301), .C1(new_n1008), .C2(new_n1009), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1007), .A2(new_n1012), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT54), .ZN(new_n1022));
  AND2_X1   g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n982), .A2(new_n987), .A3(new_n988), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(new_n707), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n994), .A2(new_n996), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(new_n701), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1025), .A2(G168), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(G8), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1029), .A2(KEYINPUT120), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(KEYINPUT51), .ZN(new_n1032));
  AOI22_X1  g607(.A1(new_n1024), .A2(new_n707), .B1(new_n1026), .B2(new_n701), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1033), .A2(new_n1029), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(G286), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT51), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1028), .A2(new_n1036), .A3(new_n1030), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1032), .A2(new_n1035), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT123), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n531), .A2(G8), .A3(new_n534), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT55), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n531), .A2(new_n534), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(G2090), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n961), .A2(new_n1015), .A3(new_n1045), .A4(new_n1017), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  AND3_X1   g622(.A1(new_n1000), .A2(new_n959), .A3(new_n960), .ZN(new_n1048));
  AOI21_X1  g623(.A(G1971), .B1(new_n1048), .B2(new_n999), .ZN(new_n1049));
  OAI211_X1 g624(.A(G8), .B(new_n1044), .C1(new_n1047), .C2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n965), .A2(new_n959), .A3(new_n960), .ZN(new_n1051));
  OR2_X1    g626(.A1(new_n583), .A2(new_n584), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1052), .A2(G1976), .A3(new_n582), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1051), .A2(G8), .A3(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(KEYINPUT52), .ZN(new_n1055));
  INV_X1    g630(.A(G1976), .ZN(new_n1056));
  AOI21_X1  g631(.A(KEYINPUT52), .B1(G288), .B2(new_n1056), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1051), .A2(new_n1053), .A3(new_n1057), .A4(G8), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n589), .A2(new_n801), .A3(new_n590), .A4(new_n591), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n588), .B1(new_n516), .B2(G61), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1060), .A2(new_n532), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n590), .A2(new_n591), .ZN(new_n1062));
  OAI21_X1  g637(.A(G1981), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  OR2_X1    g638(.A1(KEYINPUT113), .A2(KEYINPUT49), .ZN(new_n1064));
  AND3_X1   g639(.A1(new_n1059), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1064), .B1(new_n1059), .B2(new_n1063), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1067), .A2(new_n1051), .A3(G8), .ZN(new_n1068));
  AND3_X1   g643(.A1(new_n1055), .A2(new_n1058), .A3(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1050), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT114), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n514), .A2(new_n1071), .A3(new_n1016), .A4(new_n980), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1016), .B1(new_n858), .B2(new_n980), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n979), .A2(new_n1073), .ZN(new_n1074));
  OAI21_X1  g649(.A(KEYINPUT114), .B1(new_n993), .B2(KEYINPUT50), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1072), .A2(new_n1074), .A3(new_n1045), .A4(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(G1971), .ZN(new_n1077));
  INV_X1    g652(.A(new_n999), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1000), .A2(new_n959), .A3(new_n960), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1077), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1076), .A2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1044), .B1(new_n1081), .B2(G8), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1039), .B1(new_n1070), .B2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1019), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1022), .B1(new_n1084), .B2(G171), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1006), .A2(G301), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1081), .A2(G8), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1044), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1055), .A2(new_n1058), .A3(new_n1068), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1029), .B1(new_n1080), .B2(new_n1046), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1091), .B1(new_n1092), .B2(new_n1044), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1090), .A2(new_n1093), .A3(KEYINPUT123), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1038), .A2(new_n1083), .A3(new_n1087), .A4(new_n1094), .ZN(new_n1095));
  OAI21_X1  g670(.A(KEYINPUT124), .B1(new_n1023), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1030), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1098), .B1(new_n1033), .B2(G168), .ZN(new_n1099));
  AOI22_X1  g674(.A1(new_n1099), .A2(new_n1036), .B1(new_n1034), .B2(G286), .ZN(new_n1100));
  AOI22_X1  g675(.A1(new_n1100), .A2(new_n1032), .B1(new_n1086), .B2(new_n1085), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT124), .ZN(new_n1102));
  AND2_X1   g677(.A1(new_n1083), .A2(new_n1094), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1097), .A2(new_n1101), .A3(new_n1102), .A4(new_n1103), .ZN(new_n1104));
  XNOR2_X1  g679(.A(G299), .B(KEYINPUT117), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT57), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1106), .B1(new_n575), .B2(KEYINPUT116), .ZN(new_n1107));
  XNOR2_X1  g682(.A(new_n1105), .B(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1072), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1110));
  XNOR2_X1  g685(.A(KEYINPUT56), .B(G2072), .ZN(new_n1111));
  AOI22_X1  g686(.A1(new_n1109), .A2(new_n763), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1108), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(G2067), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1051), .ZN(new_n1115));
  AOI22_X1  g690(.A1(new_n1018), .A2(new_n791), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1116), .A2(new_n611), .ZN(new_n1117));
  XOR2_X1   g692(.A(new_n1117), .B(KEYINPUT118), .Z(new_n1118));
  NOR2_X1   g693(.A1(new_n1108), .A2(new_n1112), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1113), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  AOI211_X1 g695(.A(KEYINPUT119), .B(KEYINPUT61), .C1(new_n1108), .C2(new_n1112), .ZN(new_n1121));
  AND3_X1   g696(.A1(new_n1108), .A2(KEYINPUT61), .A3(new_n1112), .ZN(new_n1122));
  NOR3_X1   g697(.A1(new_n1121), .A2(new_n1119), .A3(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1048), .A2(new_n999), .ZN(new_n1124));
  XNOR2_X1  g699(.A(KEYINPUT58), .B(G1341), .ZN(new_n1125));
  OAI22_X1  g700(.A1(new_n1124), .A2(G1996), .B1(new_n1115), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(new_n562), .ZN(new_n1127));
  XNOR2_X1  g702(.A(new_n1127), .B(KEYINPUT59), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT60), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1116), .A2(new_n1129), .A3(new_n612), .ZN(new_n1130));
  XNOR2_X1  g705(.A(new_n1116), .B(new_n612), .ZN(new_n1131));
  OAI211_X1 g706(.A(new_n1128), .B(new_n1130), .C1(new_n1129), .C2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1120), .B1(new_n1123), .B2(new_n1132), .ZN(new_n1133));
  AND3_X1   g708(.A1(new_n1096), .A2(new_n1104), .A3(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1068), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1052), .A2(new_n1056), .A3(new_n582), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1059), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1137), .A2(G8), .A3(new_n1051), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1138), .B1(new_n1050), .B2(new_n1091), .ZN(new_n1139));
  NOR3_X1   g714(.A1(new_n1033), .A2(new_n1029), .A3(G286), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1140), .A2(new_n1090), .A3(new_n1093), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT63), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1092), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1142), .B1(new_n1144), .B2(new_n1089), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1145), .A2(new_n1140), .A3(new_n1093), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1139), .B1(new_n1143), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT62), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1032), .A2(new_n1148), .A3(new_n1035), .A4(new_n1037), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT125), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1007), .A2(new_n1012), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1103), .A2(new_n1149), .A3(new_n1150), .A4(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1099), .A2(new_n1036), .ZN(new_n1154));
  OAI21_X1  g729(.A(KEYINPUT62), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT126), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1038), .A2(KEYINPUT126), .A3(KEYINPUT62), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1152), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  NOR3_X1   g734(.A1(new_n1006), .A2(KEYINPUT122), .A3(G301), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1011), .B1(new_n1010), .B2(G171), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1083), .A2(new_n1094), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1150), .B1(new_n1164), .B2(new_n1149), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1147), .B1(new_n1159), .B2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n978), .B1(new_n1134), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n821), .A2(new_n823), .ZN(new_n1168));
  OR2_X1    g743(.A1(new_n975), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n778), .A2(new_n1114), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n969), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT48), .ZN(new_n1172));
  OR3_X1    g747(.A1(new_n969), .A2(G1986), .A3(G290), .ZN(new_n1173));
  AOI22_X1  g748(.A1(new_n976), .A2(new_n970), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  OR2_X1    g749(.A1(new_n1173), .A2(new_n1172), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1171), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n969), .B1(new_n973), .B2(new_n733), .ZN(new_n1177));
  OR3_X1    g752(.A1(new_n969), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1178));
  OAI21_X1  g753(.A(KEYINPUT46), .B1(new_n969), .B2(G1996), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1177), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  XOR2_X1   g755(.A(new_n1180), .B(KEYINPUT47), .Z(new_n1181));
  NAND2_X1  g756(.A1(new_n1176), .A2(new_n1181), .ZN(new_n1182));
  XNOR2_X1  g757(.A(new_n1182), .B(KEYINPUT127), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1167), .A2(new_n1183), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g759(.A(G229), .ZN(new_n1186));
  NOR3_X1   g760(.A1(G227), .A2(new_n460), .A3(G401), .ZN(new_n1187));
  NAND3_X1  g761(.A1(new_n886), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1188));
  NOR2_X1   g762(.A1(new_n1188), .A2(new_n953), .ZN(G308));
  AND2_X1   g763(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1190));
  AND2_X1   g764(.A1(new_n952), .A2(KEYINPUT43), .ZN(new_n1191));
  OAI211_X1 g765(.A(new_n1190), .B(new_n886), .C1(new_n1191), .C2(new_n951), .ZN(G225));
endmodule


