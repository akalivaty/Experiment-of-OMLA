//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 1 0 1 0 1 1 0 0 1 1 1 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 1 1 0 1 1 1 0 1 0 1 1 0 0 1 0 1 0 1 1 1 0 0 0 1 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:01 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n716, new_n717, new_n718, new_n719, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n768, new_n769, new_n770, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT31), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT69), .ZN(new_n189));
  INV_X1    g003(.A(G116), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n190), .A2(G119), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT68), .ZN(new_n192));
  INV_X1    g006(.A(G119), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n192), .B1(new_n193), .B2(G116), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n190), .A2(KEYINPUT68), .A3(G119), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n191), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  XNOR2_X1  g010(.A(KEYINPUT2), .B(G113), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n189), .B1(new_n196), .B2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n193), .A2(G116), .ZN(new_n200));
  AND3_X1   g014(.A1(new_n190), .A2(KEYINPUT68), .A3(G119), .ZN(new_n201));
  AOI21_X1  g015(.A(KEYINPUT68), .B1(new_n190), .B2(G119), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n200), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(new_n197), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n199), .A2(new_n204), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n203), .A2(new_n189), .A3(new_n197), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G137), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n208), .B1(KEYINPUT11), .B2(G134), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT11), .ZN(new_n210));
  INV_X1    g024(.A(G134), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT65), .ZN(new_n213));
  XNOR2_X1  g027(.A(KEYINPUT64), .B(G137), .ZN(new_n214));
  AND2_X1   g028(.A1(KEYINPUT11), .A2(G134), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n208), .A2(KEYINPUT64), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT64), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G137), .ZN(new_n219));
  AND4_X1   g033(.A1(new_n213), .A2(new_n217), .A3(new_n219), .A4(new_n215), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n212), .B1(new_n216), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G131), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT66), .ZN(new_n223));
  INV_X1    g037(.A(G131), .ZN(new_n224));
  OAI211_X1 g038(.A(new_n224), .B(new_n212), .C1(new_n216), .C2(new_n220), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n222), .A2(new_n223), .A3(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n221), .A2(KEYINPUT66), .A3(G131), .ZN(new_n227));
  XNOR2_X1  g041(.A(G143), .B(G146), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n228), .A2(KEYINPUT0), .A3(G128), .ZN(new_n229));
  XNOR2_X1  g043(.A(KEYINPUT0), .B(G128), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n229), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n226), .A2(new_n227), .A3(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G128), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n234), .A2(KEYINPUT1), .ZN(new_n235));
  INV_X1    g049(.A(G143), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G146), .ZN(new_n237));
  INV_X1    g051(.A(G146), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G143), .ZN(new_n239));
  OAI22_X1  g053(.A1(new_n235), .A2(new_n237), .B1(new_n239), .B2(G128), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(KEYINPUT67), .B1(new_n228), .B2(new_n235), .ZN(new_n242));
  AND4_X1   g056(.A1(KEYINPUT67), .A2(new_n235), .A3(new_n239), .A4(new_n237), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n241), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  OAI21_X1  g058(.A(G131), .B1(new_n211), .B2(new_n208), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n245), .B1(new_n214), .B2(new_n211), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n225), .A2(new_n244), .A3(new_n247), .ZN(new_n248));
  AOI21_X1  g062(.A(KEYINPUT30), .B1(new_n233), .B2(new_n248), .ZN(new_n249));
  AND3_X1   g063(.A1(new_n226), .A2(new_n227), .A3(new_n232), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n248), .A2(KEYINPUT70), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n235), .A2(new_n239), .A3(new_n237), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT67), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n228), .A2(KEYINPUT67), .A3(new_n235), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n246), .B1(new_n256), .B2(new_n241), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT70), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n257), .A2(new_n258), .A3(new_n225), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n251), .A2(KEYINPUT30), .A3(new_n259), .ZN(new_n260));
  OAI21_X1  g074(.A(KEYINPUT71), .B1(new_n250), .B2(new_n260), .ZN(new_n261));
  AND4_X1   g075(.A1(new_n258), .A2(new_n225), .A3(new_n244), .A4(new_n247), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n258), .B1(new_n257), .B2(new_n225), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT71), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n264), .A2(new_n265), .A3(new_n233), .A4(KEYINPUT30), .ZN(new_n266));
  AOI211_X1 g080(.A(new_n207), .B(new_n249), .C1(new_n261), .C2(new_n266), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n233), .A2(new_n207), .A3(new_n251), .A4(new_n259), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT73), .ZN(new_n269));
  INV_X1    g083(.A(G953), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(KEYINPUT73), .A2(G953), .ZN(new_n272));
  AND2_X1   g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  XNOR2_X1  g087(.A(KEYINPUT72), .B(G237), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n273), .A2(G210), .A3(new_n274), .ZN(new_n275));
  OR2_X1    g089(.A1(new_n275), .A2(KEYINPUT27), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(KEYINPUT27), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g092(.A(KEYINPUT26), .B(G101), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n276), .A2(new_n277), .A3(new_n279), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n268), .A2(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n188), .B1(new_n267), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n261), .A2(new_n266), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n249), .A2(new_n207), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n285), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n289), .A2(KEYINPUT31), .A3(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT28), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n233), .A2(new_n248), .ZN(new_n293));
  INV_X1    g107(.A(new_n207), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n292), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n293), .A2(new_n294), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n264), .A2(KEYINPUT28), .A3(new_n233), .A4(new_n207), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT74), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n283), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n281), .A2(KEYINPUT74), .A3(new_n282), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  AOI22_X1  g117(.A1(new_n286), .A2(new_n291), .B1(new_n298), .B2(new_n303), .ZN(new_n304));
  NOR2_X1   g118(.A1(G472), .A2(G902), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n187), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(KEYINPUT75), .ZN(new_n308));
  INV_X1    g122(.A(G472), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT29), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n295), .A2(new_n296), .A3(new_n297), .A4(new_n302), .ZN(new_n311));
  INV_X1    g125(.A(new_n268), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n312), .B1(new_n287), .B2(new_n288), .ZN(new_n313));
  OAI211_X1 g127(.A(new_n310), .B(new_n311), .C1(new_n313), .C2(new_n284), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n251), .A2(new_n259), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n294), .B1(new_n250), .B2(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n292), .B1(new_n316), .B2(new_n268), .ZN(new_n317));
  INV_X1    g131(.A(new_n295), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n283), .A2(new_n310), .ZN(new_n320));
  AOI21_X1  g134(.A(G902), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n309), .B1(new_n314), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n286), .A2(new_n291), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n298), .A2(new_n303), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n306), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n322), .B1(new_n325), .B2(KEYINPUT32), .ZN(new_n326));
  AOI21_X1  g140(.A(KEYINPUT31), .B1(new_n289), .B2(new_n290), .ZN(new_n327));
  AOI211_X1 g141(.A(new_n188), .B(new_n285), .C1(new_n287), .C2(new_n288), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n324), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(KEYINPUT32), .B1(new_n329), .B2(new_n305), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT75), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n308), .A2(new_n326), .A3(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(G234), .ZN(new_n334));
  OAI21_X1  g148(.A(G217), .B1(new_n334), .B2(G902), .ZN(new_n335));
  XNOR2_X1  g149(.A(new_n335), .B(KEYINPUT76), .ZN(new_n336));
  INV_X1    g150(.A(G221), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n337), .A2(new_n334), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n273), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(KEYINPUT77), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT77), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n273), .A2(new_n341), .A3(new_n338), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  XNOR2_X1  g157(.A(KEYINPUT22), .B(G137), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n340), .A2(new_n342), .A3(new_n344), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT23), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n349), .B1(new_n193), .B2(G128), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n234), .A2(KEYINPUT23), .A3(G119), .ZN(new_n351));
  OAI211_X1 g165(.A(new_n350), .B(new_n351), .C1(G119), .C2(new_n234), .ZN(new_n352));
  XNOR2_X1  g166(.A(G119), .B(G128), .ZN(new_n353));
  XOR2_X1   g167(.A(KEYINPUT24), .B(G110), .Z(new_n354));
  OAI22_X1  g168(.A1(new_n352), .A2(G110), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  XNOR2_X1  g169(.A(G125), .B(G140), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(KEYINPUT16), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT16), .ZN(new_n358));
  INV_X1    g172(.A(G140), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n358), .A2(new_n359), .A3(G125), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n357), .A2(G146), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n359), .A2(G125), .ZN(new_n362));
  INV_X1    g176(.A(G125), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(G140), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n355), .B(new_n361), .C1(G146), .C2(new_n365), .ZN(new_n366));
  AOI22_X1  g180(.A1(new_n352), .A2(G110), .B1(new_n353), .B2(new_n354), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n360), .B1(new_n365), .B2(new_n358), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n368), .A2(new_n238), .ZN(new_n369));
  AOI21_X1  g183(.A(G146), .B1(new_n357), .B2(new_n360), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n367), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n366), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n348), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(G902), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n346), .A2(new_n366), .A3(new_n371), .A4(new_n347), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n373), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT25), .ZN(new_n377));
  AND2_X1   g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n376), .A2(new_n377), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n336), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  AND2_X1   g194(.A1(new_n373), .A2(new_n375), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n336), .A2(G902), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n382), .B(KEYINPUT78), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n380), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(G104), .ZN(new_n387));
  OAI21_X1  g201(.A(KEYINPUT3), .B1(new_n387), .B2(G107), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT3), .ZN(new_n389));
  INV_X1    g203(.A(G107), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n389), .A2(new_n390), .A3(G104), .ZN(new_n391));
  INV_X1    g205(.A(G101), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n387), .A2(G107), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n388), .A2(new_n391), .A3(new_n392), .A4(new_n393), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n387), .A2(G107), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n390), .A2(G104), .ZN(new_n396));
  OAI21_X1  g210(.A(G101), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n394), .A2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n244), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n240), .B1(new_n254), .B2(new_n255), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(new_n398), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n226), .A2(new_n403), .A3(new_n227), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT12), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n226), .A2(new_n403), .A3(KEYINPUT12), .A4(new_n227), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n388), .A2(new_n391), .A3(new_n393), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT4), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n409), .A2(new_n410), .A3(G101), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n409), .A2(G101), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n412), .A2(KEYINPUT4), .A3(new_n394), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n232), .A2(new_n411), .A3(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT10), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n415), .B1(new_n401), .B2(new_n398), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n244), .A2(KEYINPUT10), .A3(new_n399), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n414), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n226), .A2(new_n227), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n408), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n273), .A2(G227), .ZN(new_n423));
  XOR2_X1   g237(.A(G110), .B(G140), .Z(new_n424));
  XNOR2_X1  g238(.A(new_n423), .B(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(KEYINPUT79), .B1(new_n419), .B2(new_n420), .ZN(new_n426));
  AND2_X1   g240(.A1(new_n226), .A2(new_n227), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT79), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n427), .A2(new_n428), .A3(new_n418), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n425), .B1(new_n419), .B2(new_n420), .ZN(new_n431));
  AOI22_X1  g245(.A1(new_n422), .A2(new_n425), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(G469), .B1(new_n432), .B2(G902), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n408), .A2(new_n431), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n427), .A2(new_n418), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n435), .B1(new_n429), .B2(new_n426), .ZN(new_n436));
  INV_X1    g250(.A(new_n425), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n434), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(G469), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n438), .A2(new_n439), .A3(new_n374), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n433), .A2(new_n440), .ZN(new_n441));
  OAI21_X1  g255(.A(G214), .B1(G237), .B2(G902), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(G210), .B1(G237), .B2(G902), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n205), .A2(new_n206), .A3(new_n411), .A4(new_n413), .ZN(new_n446));
  OAI211_X1 g260(.A(KEYINPUT5), .B(new_n200), .C1(new_n201), .C2(new_n202), .ZN(new_n447));
  INV_X1    g261(.A(G113), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT5), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n448), .B1(new_n191), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n196), .A2(new_n198), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n399), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n446), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g268(.A(G110), .B(G122), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n446), .A2(new_n453), .A3(new_n455), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT6), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n459), .A2(KEYINPUT80), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n457), .A2(new_n458), .A3(new_n460), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n454), .B(new_n456), .C1(KEYINPUT80), .C2(new_n459), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n229), .B(G125), .C1(new_n228), .C2(new_n230), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n463), .B1(new_n401), .B2(G125), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n270), .A2(G224), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n464), .B(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n461), .A2(new_n462), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n465), .A2(KEYINPUT7), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n464), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n468), .ZN(new_n470));
  OAI211_X1 g284(.A(new_n463), .B(new_n470), .C1(new_n401), .C2(G125), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT82), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT81), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n394), .A2(new_n397), .A3(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n451), .A2(new_n475), .A3(new_n452), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n455), .B(KEYINPUT8), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n475), .B1(new_n451), .B2(new_n452), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n473), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n451), .A2(new_n452), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n481), .A2(new_n474), .A3(new_n399), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n482), .A2(KEYINPUT82), .A3(new_n477), .A4(new_n476), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n472), .A2(new_n480), .A3(new_n483), .A4(new_n458), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT83), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n484), .A2(new_n485), .A3(new_n374), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n467), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n485), .B1(new_n484), .B2(new_n374), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n445), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n484), .A2(new_n374), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(KEYINPUT83), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n491), .A2(new_n444), .A3(new_n467), .A4(new_n486), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n443), .B1(new_n489), .B2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(G952), .ZN(new_n494));
  AOI211_X1 g308(.A(G953), .B(new_n494), .C1(G234), .C2(G237), .ZN(new_n495));
  AOI211_X1 g309(.A(new_n374), .B(new_n273), .C1(G234), .C2(G237), .ZN(new_n496));
  XNOR2_X1  g310(.A(KEYINPUT21), .B(G898), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  XNOR2_X1  g313(.A(KEYINPUT9), .B(G234), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n337), .B1(new_n501), .B2(new_n374), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n441), .A2(new_n493), .A3(new_n499), .A4(new_n503), .ZN(new_n504));
  XNOR2_X1  g318(.A(G113), .B(G122), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n505), .B(new_n387), .ZN(new_n506));
  AND2_X1   g320(.A1(KEYINPUT72), .A2(G237), .ZN(new_n507));
  NOR2_X1   g321(.A1(KEYINPUT72), .A2(G237), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n271), .B(new_n272), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(G214), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n236), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n273), .A2(G143), .A3(G214), .A4(new_n274), .ZN(new_n512));
  AND3_X1   g326(.A1(new_n511), .A2(new_n512), .A3(new_n224), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n224), .B1(new_n511), .B2(new_n512), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(KEYINPUT85), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT85), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n517), .B1(new_n513), .B2(new_n514), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n356), .B(KEYINPUT19), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n369), .B1(new_n238), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n516), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(KEYINPUT18), .A2(G131), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n511), .A2(new_n512), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT84), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n511), .A2(new_n512), .A3(KEYINPUT84), .A4(new_n522), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n356), .B(new_n238), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n506), .B1(new_n521), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT88), .ZN(new_n532));
  AND3_X1   g346(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT17), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT86), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n535), .B1(new_n369), .B2(new_n370), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n368), .A2(new_n238), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n537), .A2(KEYINPUT86), .A3(new_n361), .ZN(new_n538));
  AOI22_X1  g352(.A1(new_n515), .A2(new_n534), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT87), .ZN(new_n540));
  AND4_X1   g354(.A1(new_n540), .A2(new_n524), .A3(KEYINPUT17), .A4(G131), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n540), .B1(new_n514), .B2(KEYINPUT17), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n533), .B1(new_n539), .B2(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n532), .B1(new_n544), .B2(new_n506), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n524), .A2(G131), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n511), .A2(new_n512), .A3(new_n224), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n546), .A2(new_n534), .A3(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n524), .A2(KEYINPUT17), .A3(G131), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(KEYINPUT87), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n536), .A2(new_n538), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n514), .A2(new_n540), .A3(KEYINPUT17), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n548), .A2(new_n550), .A3(new_n551), .A4(new_n552), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n553), .A2(new_n532), .A3(new_n506), .A4(new_n529), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n531), .B1(new_n545), .B2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT20), .ZN(new_n557));
  NOR2_X1   g371(.A1(G475), .A2(G902), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n553), .A2(new_n506), .A3(new_n529), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(KEYINPUT88), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n530), .B1(new_n561), .B2(new_n554), .ZN(new_n562));
  INV_X1    g376(.A(new_n558), .ZN(new_n563));
  OAI21_X1  g377(.A(KEYINPUT20), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n559), .A2(new_n564), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n544), .A2(new_n506), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n566), .B1(new_n554), .B2(new_n561), .ZN(new_n567));
  OAI21_X1  g381(.A(G475), .B1(new_n567), .B2(G902), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n501), .A2(G217), .A3(new_n270), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  XNOR2_X1  g384(.A(G128), .B(G143), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(new_n211), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n572), .B(KEYINPUT89), .ZN(new_n573));
  XOR2_X1   g387(.A(G116), .B(G122), .Z(new_n574));
  XNOR2_X1  g388(.A(new_n574), .B(G107), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n571), .A2(KEYINPUT13), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n236), .A2(G128), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n576), .B(G134), .C1(KEYINPUT13), .C2(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n573), .A2(new_n575), .A3(new_n578), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n571), .B(new_n211), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n190), .A2(KEYINPUT14), .A3(G122), .ZN(new_n581));
  OAI211_X1 g395(.A(G107), .B(new_n581), .C1(new_n574), .C2(KEYINPUT14), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n580), .B(new_n582), .C1(G107), .C2(new_n574), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n570), .B1(new_n579), .B2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n579), .A2(new_n583), .A3(new_n570), .ZN(new_n586));
  AOI21_X1  g400(.A(G902), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT15), .ZN(new_n588));
  AND2_X1   g402(.A1(new_n588), .A2(KEYINPUT90), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n588), .A2(KEYINPUT90), .ZN(new_n590));
  OAI21_X1  g404(.A(G478), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  XOR2_X1   g405(.A(new_n587), .B(new_n591), .Z(new_n592));
  NAND3_X1  g406(.A1(new_n565), .A2(new_n568), .A3(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n504), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n333), .A2(new_n386), .A3(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n595), .B(G101), .ZN(G3));
  AOI21_X1  g410(.A(new_n309), .B1(new_n329), .B2(new_n374), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n597), .A2(new_n325), .ZN(new_n598));
  AND3_X1   g412(.A1(new_n438), .A2(new_n439), .A3(new_n374), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n422), .A2(new_n425), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n430), .A2(new_n431), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n600), .A2(G469), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(G469), .A2(G902), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n503), .B1(new_n599), .B2(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n605), .A2(new_n385), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n598), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT91), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n489), .A2(new_n492), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n608), .B1(new_n609), .B2(new_n442), .ZN(new_n610));
  AOI211_X1 g424(.A(KEYINPUT91), .B(new_n443), .C1(new_n489), .C2(new_n492), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n557), .B1(new_n556), .B2(new_n558), .ZN(new_n613));
  NOR3_X1   g427(.A1(new_n562), .A2(KEYINPUT20), .A3(new_n563), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n568), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT92), .ZN(new_n616));
  INV_X1    g430(.A(new_n586), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n616), .B1(new_n617), .B2(new_n584), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT33), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OAI211_X1 g434(.A(new_n616), .B(KEYINPUT33), .C1(new_n617), .C2(new_n584), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n620), .A2(G478), .A3(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(G478), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n623), .A2(new_n374), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n624), .B1(new_n587), .B2(new_n623), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(KEYINPUT93), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT93), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n622), .A2(new_n628), .A3(new_n625), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n615), .A2(new_n631), .ZN(new_n632));
  NOR4_X1   g446(.A1(new_n607), .A2(new_n498), .A3(new_n612), .A4(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(new_n387), .ZN(new_n634));
  XNOR2_X1  g448(.A(KEYINPUT94), .B(KEYINPUT34), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G6));
  INV_X1    g450(.A(new_n592), .ZN(new_n637));
  AND2_X1   g451(.A1(new_n568), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n559), .A2(KEYINPUT95), .A3(new_n564), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  AOI21_X1  g454(.A(KEYINPUT95), .B1(new_n559), .B2(new_n564), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n638), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NOR3_X1   g456(.A1(new_n642), .A2(new_n612), .A3(new_n498), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n643), .A2(new_n598), .A3(new_n606), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT35), .B(G107), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G9));
  NOR2_X1   g460(.A1(new_n348), .A2(KEYINPUT36), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(new_n372), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n383), .ZN(new_n649));
  AND2_X1   g463(.A1(new_n380), .A2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n594), .A2(new_n598), .A3(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT37), .B(G110), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G12));
  INV_X1    g468(.A(G900), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n495), .B1(new_n496), .B2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  OAI211_X1 g471(.A(new_n638), .B(new_n657), .C1(new_n640), .C2(new_n641), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(KEYINPUT96), .ZN(new_n659));
  INV_X1    g473(.A(new_n641), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n639), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT96), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n661), .A2(new_n662), .A3(new_n638), .A4(new_n657), .ZN(new_n663));
  AND2_X1   g477(.A1(new_n659), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n605), .A2(new_n650), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n665), .B1(new_n610), .B2(new_n611), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n329), .A2(new_n305), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n331), .B1(new_n667), .B2(new_n187), .ZN(new_n668));
  AOI211_X1 g482(.A(KEYINPUT75), .B(KEYINPUT32), .C1(new_n329), .C2(new_n305), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n666), .B1(new_n670), .B2(new_n326), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT97), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n664), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  NOR3_X1   g487(.A1(new_n612), .A2(new_n605), .A3(new_n650), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n333), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n659), .A2(new_n663), .ZN(new_n676));
  OAI21_X1  g490(.A(KEYINPUT97), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n673), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G128), .ZN(G30));
  INV_X1    g493(.A(KEYINPUT100), .ZN(new_n680));
  AND2_X1   g494(.A1(new_n316), .A2(new_n268), .ZN(new_n681));
  OAI22_X1  g495(.A1(new_n267), .A2(new_n285), .B1(new_n302), .B2(new_n681), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n309), .B1(new_n682), .B2(new_n374), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n683), .B1(new_n325), .B2(KEYINPUT32), .ZN(new_n684));
  AND3_X1   g498(.A1(new_n670), .A2(new_n680), .A3(new_n684), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n680), .B1(new_n670), .B2(new_n684), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(KEYINPUT101), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n615), .A2(new_n637), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  XOR2_X1   g504(.A(KEYINPUT98), .B(KEYINPUT38), .Z(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(KEYINPUT99), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n609), .B(new_n692), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n690), .A2(new_n442), .A3(new_n650), .A4(new_n693), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n502), .B1(new_n433), .B2(new_n440), .ZN(new_n695));
  XOR2_X1   g509(.A(new_n656), .B(KEYINPUT39), .Z(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(KEYINPUT40), .ZN(new_n698));
  OR3_X1    g512(.A1(new_n688), .A2(new_n694), .A3(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G143), .ZN(G45));
  NAND3_X1  g514(.A1(new_n615), .A2(new_n631), .A3(new_n657), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n675), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(new_n238), .ZN(G48));
  NAND2_X1  g517(.A1(KEYINPUT102), .A2(G469), .ZN(new_n704));
  AND3_X1   g518(.A1(new_n438), .A2(new_n374), .A3(new_n704), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n704), .B1(new_n438), .B2(new_n374), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n503), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n708), .A2(new_n385), .ZN(new_n709));
  NOR3_X1   g523(.A1(new_n612), .A2(new_n632), .A3(new_n498), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n333), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(KEYINPUT41), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G113), .ZN(G15));
  NAND3_X1  g527(.A1(new_n643), .A2(new_n333), .A3(new_n709), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G116), .ZN(G18));
  NOR2_X1   g529(.A1(new_n650), .A2(new_n498), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n716), .A2(new_n565), .A3(new_n568), .A4(new_n592), .ZN(new_n717));
  NOR3_X1   g531(.A1(new_n612), .A2(new_n708), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n333), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G119), .ZN(G21));
  INV_X1    g534(.A(new_n706), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n438), .A2(new_n374), .A3(new_n704), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n721), .A2(new_n499), .A3(new_n503), .A4(new_n722), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n612), .A2(new_n689), .A3(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(new_n317), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT103), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n725), .A2(new_n726), .A3(new_n295), .ZN(new_n727));
  OAI21_X1  g541(.A(KEYINPUT103), .B1(new_n317), .B2(new_n318), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n727), .A2(new_n728), .A3(new_n303), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n306), .B1(new_n323), .B2(new_n729), .ZN(new_n730));
  NOR3_X1   g544(.A1(new_n597), .A2(new_n730), .A3(new_n385), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n724), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G122), .ZN(G24));
  NOR3_X1   g547(.A1(new_n597), .A2(new_n730), .A3(new_n650), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n612), .A2(new_n708), .ZN(new_n735));
  INV_X1    g549(.A(new_n701), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n734), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(KEYINPUT104), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT104), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n734), .A2(new_n735), .A3(new_n739), .A4(new_n736), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G125), .ZN(G27));
  INV_X1    g556(.A(KEYINPUT42), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n489), .A2(new_n442), .A3(new_n492), .ZN(new_n744));
  INV_X1    g558(.A(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n695), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n701), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n333), .A2(new_n386), .A3(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT105), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n329), .A2(KEYINPUT32), .A3(new_n305), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n311), .A2(new_n310), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n289), .A2(new_n268), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n751), .B1(new_n283), .B2(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n725), .A2(new_n295), .A3(new_n320), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(new_n374), .ZN(new_n755));
  OAI21_X1  g569(.A(G472), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n750), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n386), .B1(new_n757), .B2(new_n330), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n605), .A2(new_n744), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n630), .B1(new_n565), .B2(new_n568), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n759), .A2(KEYINPUT42), .A3(new_n760), .A4(new_n657), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n749), .B1(new_n758), .B2(new_n761), .ZN(new_n762));
  NOR3_X1   g576(.A1(new_n701), .A2(new_n746), .A3(new_n743), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n307), .A2(new_n750), .A3(new_n756), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n763), .A2(KEYINPUT105), .A3(new_n386), .A4(new_n764), .ZN(new_n765));
  AOI22_X1  g579(.A1(new_n743), .A2(new_n748), .B1(new_n762), .B2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(new_n224), .ZN(G33));
  NAND3_X1  g581(.A1(new_n333), .A2(new_n386), .A3(new_n759), .ZN(new_n768));
  INV_X1    g582(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(new_n664), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G134), .ZN(G36));
  INV_X1    g585(.A(new_n615), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(new_n631), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(KEYINPUT43), .ZN(new_n774));
  NOR3_X1   g588(.A1(new_n774), .A2(new_n598), .A3(new_n650), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n744), .B1(new_n775), .B2(KEYINPUT44), .ZN(new_n776));
  OR2_X1    g590(.A1(new_n432), .A2(KEYINPUT45), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n432), .A2(KEYINPUT45), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n777), .A2(G469), .A3(new_n778), .ZN(new_n779));
  AOI21_X1  g593(.A(KEYINPUT46), .B1(new_n779), .B2(new_n603), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n780), .A2(new_n599), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n779), .A2(KEYINPUT46), .A3(new_n603), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n502), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n783), .A2(new_n696), .ZN(new_n784));
  OAI211_X1 g598(.A(new_n776), .B(new_n784), .C1(KEYINPUT44), .C2(new_n775), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G137), .ZN(G39));
  XNOR2_X1  g600(.A(new_n783), .B(KEYINPUT47), .ZN(new_n787));
  NOR3_X1   g601(.A1(new_n668), .A2(new_n669), .A3(new_n757), .ZN(new_n788));
  NOR3_X1   g602(.A1(new_n701), .A2(new_n386), .A3(new_n744), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n787), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(KEYINPUT106), .B(G140), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n790), .B(new_n791), .ZN(G42));
  NOR4_X1   g606(.A1(new_n773), .A2(new_n385), .A3(new_n443), .A4(new_n502), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  OR2_X1    g608(.A1(new_n794), .A2(KEYINPUT107), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(KEYINPUT107), .ZN(new_n796));
  XOR2_X1   g610(.A(new_n707), .B(KEYINPUT49), .Z(new_n797));
  NOR2_X1   g611(.A1(new_n797), .A2(new_n693), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n688), .A2(new_n795), .A3(new_n796), .A4(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(new_n495), .ZN(new_n800));
  NOR4_X1   g614(.A1(new_n774), .A2(new_n800), .A3(new_n708), .A4(new_n744), .ZN(new_n801));
  INV_X1    g615(.A(new_n758), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(KEYINPUT48), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n774), .A2(new_n800), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n805), .A2(new_n731), .ZN(new_n806));
  AOI211_X1 g620(.A(new_n494), .B(G953), .C1(new_n806), .C2(new_n735), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n804), .A2(new_n807), .ZN(new_n808));
  NOR4_X1   g622(.A1(new_n708), .A2(new_n385), .A3(new_n800), .A4(new_n744), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n688), .A2(new_n809), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n808), .B1(new_n760), .B2(new_n810), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n693), .A2(new_n708), .A3(new_n442), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n806), .A2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT50), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n813), .B(new_n814), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n806), .A2(KEYINPUT114), .A3(new_n745), .ZN(new_n816));
  AOI21_X1  g630(.A(KEYINPUT114), .B1(new_n806), .B2(new_n745), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n705), .A2(new_n706), .A3(new_n503), .ZN(new_n818));
  OAI22_X1  g632(.A1(new_n816), .A2(new_n817), .B1(new_n787), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n801), .A2(new_n734), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n815), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n688), .A2(new_n772), .A3(new_n630), .A4(new_n809), .ZN(new_n822));
  OR2_X1    g636(.A1(new_n822), .A2(KEYINPUT115), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(KEYINPUT115), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n821), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n811), .B1(new_n825), .B2(KEYINPUT51), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(KEYINPUT51), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(KEYINPUT116), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT116), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n825), .A2(new_n829), .A3(KEYINPUT51), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n826), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n612), .A2(new_n689), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n605), .A2(new_n651), .A3(new_n656), .ZN(new_n833));
  OAI211_X1 g647(.A(new_n832), .B(new_n833), .C1(new_n685), .C2(new_n686), .ZN(new_n834));
  AOI22_X1  g648(.A1(new_n738), .A2(new_n740), .B1(new_n671), .B2(new_n736), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n678), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT52), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n678), .A2(new_n834), .A3(new_n835), .A4(KEYINPUT52), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  AND4_X1   g654(.A1(new_n568), .A2(new_n745), .A3(new_n592), .A4(new_n657), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n333), .A2(new_n661), .A3(new_n665), .A4(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n734), .A2(new_n736), .A3(new_n759), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n842), .B(new_n843), .C1(new_n768), .C2(new_n676), .ZN(new_n844));
  AOI22_X1  g658(.A1(new_n333), .A2(new_n718), .B1(new_n724), .B2(new_n731), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n845), .A2(new_n714), .A3(new_n711), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n766), .A2(new_n844), .A3(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n609), .A2(new_n499), .A3(new_n442), .ZN(new_n848));
  INV_X1    g662(.A(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n598), .A2(new_n849), .A3(new_n760), .A4(new_n606), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n595), .A2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT108), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n595), .A2(KEYINPUT108), .A3(new_n850), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n615), .A2(new_n848), .A3(new_n592), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n598), .A2(new_n855), .A3(new_n606), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n652), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n857), .A2(KEYINPUT109), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT109), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n652), .A2(new_n856), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n853), .A2(new_n854), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g676(.A(KEYINPUT110), .B1(new_n847), .B2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n841), .A2(new_n665), .A3(new_n661), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n843), .B1(new_n788), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n865), .B1(new_n769), .B2(new_n664), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n845), .A2(new_n711), .A3(new_n714), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n748), .A2(new_n743), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n762), .A2(new_n765), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n866), .A2(new_n867), .A3(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n853), .A2(new_n854), .A3(new_n861), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT110), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n871), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n840), .B1(new_n863), .B2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT53), .ZN(new_n876));
  AOI21_X1  g690(.A(KEYINPUT111), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n877), .B1(new_n876), .B2(new_n875), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n847), .A2(new_n862), .A3(KEYINPUT110), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n873), .B1(new_n871), .B2(new_n872), .ZN(new_n880));
  AOI22_X1  g694(.A1(new_n879), .A2(new_n880), .B1(new_n838), .B2(new_n839), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n881), .A2(KEYINPUT111), .A3(KEYINPUT53), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n878), .A2(KEYINPUT54), .A3(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT112), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n884), .B1(new_n881), .B2(KEYINPUT53), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n875), .A2(KEYINPUT112), .A3(new_n876), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n867), .A2(new_n870), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(KEYINPUT113), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n872), .A2(new_n876), .A3(new_n844), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n888), .A2(new_n840), .A3(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n885), .A2(new_n886), .A3(new_n890), .ZN(new_n891));
  OR2_X1    g705(.A1(new_n891), .A2(KEYINPUT54), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n831), .A2(new_n883), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n494), .A2(new_n270), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n894), .B(KEYINPUT117), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n799), .B1(new_n893), .B2(new_n895), .ZN(G75));
  AND2_X1   g710(.A1(new_n891), .A2(G902), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(G210), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT56), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n461), .A2(new_n462), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(new_n466), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT55), .ZN(new_n902));
  AND3_X1   g716(.A1(new_n898), .A2(new_n899), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n902), .B1(new_n898), .B2(new_n899), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n273), .A2(G952), .ZN(new_n905));
  NOR3_X1   g719(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(G51));
  XOR2_X1   g720(.A(new_n891), .B(KEYINPUT54), .Z(new_n907));
  XNOR2_X1  g721(.A(new_n603), .B(KEYINPUT57), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n438), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n897), .A2(G469), .A3(new_n778), .A4(new_n777), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n905), .B1(new_n909), .B2(new_n910), .ZN(G54));
  NAND4_X1  g725(.A1(new_n891), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT118), .ZN(new_n913));
  AND3_X1   g727(.A1(new_n912), .A2(new_n913), .A3(new_n562), .ZN(new_n914));
  INV_X1    g728(.A(new_n905), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n915), .B1(new_n912), .B2(new_n562), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n913), .B1(new_n912), .B2(new_n562), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n914), .A2(new_n916), .A3(new_n917), .ZN(G60));
  NAND2_X1  g732(.A1(new_n620), .A2(new_n621), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n624), .B(KEYINPUT59), .Z(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n915), .B1(new_n907), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n892), .A2(new_n883), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n919), .B1(new_n923), .B2(new_n920), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n922), .A2(new_n924), .ZN(G63));
  NAND2_X1  g739(.A1(G217), .A2(G902), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(KEYINPUT119), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT60), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n891), .A2(new_n648), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(KEYINPUT120), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT120), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n891), .A2(new_n931), .A3(new_n648), .A4(new_n928), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n891), .A2(new_n928), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n381), .B(KEYINPUT121), .Z(new_n935));
  AOI21_X1  g749(.A(new_n905), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n933), .A2(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT61), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n933), .A2(KEYINPUT61), .A3(new_n936), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(G66));
  INV_X1    g755(.A(new_n497), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n270), .B1(new_n942), .B2(G224), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n872), .A2(new_n846), .ZN(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n943), .B1(new_n945), .B2(new_n273), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n900), .B1(G898), .B2(new_n273), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(KEYINPUT122), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n946), .B(new_n948), .ZN(G69));
  AOI21_X1  g763(.A(new_n249), .B1(new_n261), .B2(new_n266), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(new_n519), .ZN(new_n951));
  INV_X1    g765(.A(new_n273), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(G900), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n784), .A2(new_n832), .A3(new_n802), .ZN(new_n954));
  AND3_X1   g768(.A1(new_n785), .A2(new_n790), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n678), .A2(new_n835), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT123), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n956), .B(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n870), .A2(new_n770), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(KEYINPUT124), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n955), .A2(new_n958), .A3(new_n960), .ZN(new_n961));
  OAI211_X1 g775(.A(new_n951), .B(new_n953), .C1(new_n961), .C2(new_n952), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n699), .A2(new_n958), .ZN(new_n963));
  OR2_X1    g777(.A1(new_n963), .A2(KEYINPUT62), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n760), .B1(new_n772), .B2(new_n637), .ZN(new_n965));
  NOR3_X1   g779(.A1(new_n965), .A2(new_n697), .A3(new_n744), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n966), .A2(new_n333), .A3(new_n386), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n785), .A2(new_n790), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n968), .B1(new_n963), .B2(KEYINPUT62), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n952), .B1(new_n964), .B2(new_n969), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n962), .B1(new_n970), .B2(new_n951), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n273), .B1(G227), .B2(G900), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n971), .B(new_n972), .ZN(G72));
  XNOR2_X1  g787(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n309), .A2(new_n374), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n974), .B(new_n975), .Z(new_n976));
  NAND2_X1  g790(.A1(new_n752), .A2(new_n283), .ZN(new_n977));
  OR2_X1    g791(.A1(new_n977), .A2(KEYINPUT127), .ZN(new_n978));
  AOI22_X1  g792(.A1(new_n977), .A2(KEYINPUT127), .B1(new_n289), .B2(new_n290), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n976), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  AND3_X1   g794(.A1(new_n878), .A2(new_n882), .A3(new_n980), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n964), .A2(new_n944), .A3(new_n969), .ZN(new_n982));
  INV_X1    g796(.A(new_n976), .ZN(new_n983));
  AOI211_X1 g797(.A(new_n283), .B(new_n313), .C1(new_n982), .C2(new_n983), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n752), .A2(new_n284), .ZN(new_n985));
  INV_X1    g799(.A(new_n985), .ZN(new_n986));
  OR2_X1    g800(.A1(new_n961), .A2(new_n945), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n986), .B1(new_n987), .B2(new_n983), .ZN(new_n988));
  OR3_X1    g802(.A1(new_n988), .A2(KEYINPUT126), .A3(new_n905), .ZN(new_n989));
  OAI21_X1  g803(.A(KEYINPUT126), .B1(new_n988), .B2(new_n905), .ZN(new_n990));
  AOI211_X1 g804(.A(new_n981), .B(new_n984), .C1(new_n989), .C2(new_n990), .ZN(G57));
endmodule


