//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 0 1 0 0 0 0 0 1 0 0 1 0 0 1 1 1 0 1 0 1 1 1 0 0 0 1 1 1 0 1 0 0 0 0 1 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n738, new_n739, new_n740, new_n742, new_n743,
    new_n744, new_n745, new_n747, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n860, new_n861, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n870, new_n871,
    new_n872, new_n873, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n912, new_n913, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971;
  INV_X1    g000(.A(KEYINPUT86), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT34), .ZN(new_n203));
  NOR2_X1   g002(.A1(G127gat), .A2(G134gat), .ZN(new_n204));
  XOR2_X1   g003(.A(KEYINPUT67), .B(G127gat), .Z(new_n205));
  AOI21_X1  g004(.A(new_n204), .B1(new_n205), .B2(G134gat), .ZN(new_n206));
  INV_X1    g005(.A(G113gat), .ZN(new_n207));
  INV_X1    g006(.A(G120gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT1), .ZN(new_n210));
  NAND2_X1  g009(.A1(G113gat), .A2(G120gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  AND2_X1   g011(.A1(new_n207), .A2(KEYINPUT68), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n207), .A2(KEYINPUT68), .ZN(new_n214));
  OAI21_X1  g013(.A(G120gat), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n210), .B1(G113gat), .B2(G120gat), .ZN(new_n216));
  INV_X1    g015(.A(new_n204), .ZN(new_n217));
  NAND2_X1  g016(.A1(G127gat), .A2(G134gat), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  AOI22_X1  g018(.A1(new_n206), .A2(new_n212), .B1(new_n215), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(G169gat), .A2(G176gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(KEYINPUT23), .ZN(new_n222));
  INV_X1    g021(.A(G169gat), .ZN(new_n223));
  INV_X1    g022(.A(G176gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n222), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT25), .ZN(new_n227));
  NOR2_X1   g026(.A1(G169gat), .A2(G176gat), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n227), .B1(new_n228), .B2(KEYINPUT23), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n226), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT24), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n231), .A2(G183gat), .A3(G190gat), .ZN(new_n232));
  XNOR2_X1  g031(.A(G183gat), .B(G190gat), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n232), .B1(new_n233), .B2(new_n231), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT65), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n230), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  OAI211_X1 g035(.A(KEYINPUT65), .B(new_n232), .C1(new_n233), .C2(new_n231), .ZN(new_n237));
  NAND2_X1  g036(.A1(G183gat), .A2(G190gat), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n238), .A2(KEYINPUT24), .ZN(new_n239));
  INV_X1    g038(.A(G183gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(G190gat), .ZN(new_n241));
  INV_X1    g040(.A(G190gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(G183gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n239), .B1(new_n244), .B2(KEYINPUT24), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n223), .A2(new_n224), .A3(KEYINPUT23), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT64), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n228), .A2(KEYINPUT64), .A3(KEYINPUT23), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n245), .A2(new_n250), .A3(new_n226), .ZN(new_n251));
  AOI22_X1  g050(.A1(new_n236), .A2(new_n237), .B1(new_n251), .B2(new_n227), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT26), .ZN(new_n253));
  AND3_X1   g052(.A1(new_n225), .A2(new_n253), .A3(new_n221), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n238), .B1(new_n225), .B2(new_n253), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT27), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n256), .A2(G183gat), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n240), .A2(KEYINPUT27), .ZN(new_n258));
  OAI21_X1  g057(.A(KEYINPUT66), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n240), .A2(KEYINPUT27), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n256), .A2(G183gat), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT66), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n260), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT28), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n264), .A2(G190gat), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n259), .A2(new_n263), .A3(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n260), .A2(new_n261), .A3(new_n242), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(new_n264), .ZN(new_n268));
  AOI211_X1 g067(.A(new_n254), .B(new_n255), .C1(new_n266), .C2(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n220), .B1(new_n252), .B2(new_n269), .ZN(new_n270));
  OAI211_X1 g069(.A(new_n226), .B(new_n232), .C1(new_n233), .C2(new_n231), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n246), .A2(new_n247), .ZN(new_n272));
  AOI21_X1  g071(.A(KEYINPUT64), .B1(new_n228), .B2(KEYINPUT23), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n227), .B1(new_n271), .B2(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n231), .B1(new_n241), .B2(new_n243), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n235), .B1(new_n276), .B2(new_n239), .ZN(new_n277));
  AND2_X1   g076(.A1(new_n226), .A2(new_n229), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n277), .A2(new_n278), .A3(new_n237), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n275), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n219), .A2(new_n215), .ZN(new_n281));
  INV_X1    g080(.A(G134gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(KEYINPUT67), .B(G127gat), .ZN(new_n283));
  OAI211_X1 g082(.A(new_n212), .B(new_n217), .C1(new_n282), .C2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n281), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n266), .A2(new_n268), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n254), .A2(new_n255), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n280), .A2(new_n285), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n270), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(G227gat), .ZN(new_n291));
  INV_X1    g090(.A(G233gat), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n203), .B1(new_n290), .B2(new_n294), .ZN(new_n295));
  AOI211_X1 g094(.A(KEYINPUT34), .B(new_n293), .C1(new_n270), .C2(new_n289), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n270), .A2(new_n293), .A3(new_n289), .ZN(new_n298));
  XOR2_X1   g097(.A(G71gat), .B(G99gat), .Z(new_n299));
  XNOR2_X1  g098(.A(G15gat), .B(G43gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n299), .B(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(KEYINPUT33), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n298), .A2(KEYINPUT32), .A3(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT69), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND4_X1  g104(.A1(new_n298), .A2(KEYINPUT69), .A3(KEYINPUT32), .A4(new_n302), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n298), .A2(KEYINPUT32), .ZN(new_n308));
  INV_X1    g107(.A(new_n298), .ZN(new_n309));
  OAI211_X1 g108(.A(new_n308), .B(new_n301), .C1(new_n309), .C2(KEYINPUT33), .ZN(new_n310));
  AOI211_X1 g109(.A(KEYINPUT70), .B(new_n297), .C1(new_n307), .C2(new_n310), .ZN(new_n311));
  AND3_X1   g110(.A1(new_n307), .A2(new_n297), .A3(new_n310), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n297), .B1(new_n307), .B2(new_n310), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n311), .B1(new_n314), .B2(KEYINPUT70), .ZN(new_n315));
  INV_X1    g114(.A(G22gat), .ZN(new_n316));
  OR2_X1    g115(.A1(KEYINPUT76), .A2(G148gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(KEYINPUT76), .A2(G148gat), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n317), .A2(G141gat), .A3(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(G141gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(G148gat), .ZN(new_n321));
  OR3_X1    g120(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(G155gat), .A2(G162gat), .ZN(new_n323));
  AOI22_X1  g122(.A1(new_n319), .A2(new_n321), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(G155gat), .B(G162gat), .ZN(new_n325));
  INV_X1    g124(.A(G148gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(G141gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n321), .A2(new_n327), .ZN(new_n328));
  XNOR2_X1  g127(.A(KEYINPUT75), .B(KEYINPUT2), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n325), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n324), .A2(new_n330), .ZN(new_n331));
  XNOR2_X1  g130(.A(G197gat), .B(G204gat), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT22), .ZN(new_n333));
  INV_X1    g132(.A(G211gat), .ZN(new_n334));
  INV_X1    g133(.A(G218gat), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n333), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n332), .A2(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(G211gat), .B(G218gat), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n338), .A2(new_n332), .A3(new_n336), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT29), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT3), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n331), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n319), .A2(new_n321), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n322), .A2(new_n323), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n328), .A2(new_n329), .ZN(new_n350));
  INV_X1    g149(.A(new_n325), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n349), .A2(new_n345), .A3(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n342), .B1(new_n353), .B2(new_n343), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n316), .B1(new_n346), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n353), .A2(new_n343), .ZN(new_n356));
  INV_X1    g155(.A(new_n342), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n349), .A2(new_n352), .ZN(new_n359));
  AOI21_X1  g158(.A(KEYINPUT29), .B1(new_n340), .B2(new_n341), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n359), .B1(new_n360), .B2(KEYINPUT3), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n358), .A2(G22gat), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n355), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(G228gat), .A2(G233gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n355), .A2(new_n362), .A3(G228gat), .A4(G233gat), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n365), .A2(KEYINPUT79), .A3(new_n366), .ZN(new_n367));
  XNOR2_X1  g166(.A(G78gat), .B(G106gat), .ZN(new_n368));
  INV_X1    g167(.A(G50gat), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n368), .B(new_n369), .ZN(new_n370));
  XNOR2_X1  g169(.A(KEYINPUT78), .B(KEYINPUT31), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n370), .B(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n367), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT35), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n365), .A2(KEYINPUT79), .A3(new_n366), .A4(new_n372), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n374), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT6), .ZN(new_n378));
  XOR2_X1   g177(.A(G1gat), .B(G29gat), .Z(new_n379));
  XNOR2_X1  g178(.A(new_n379), .B(KEYINPUT0), .ZN(new_n380));
  XNOR2_X1  g179(.A(G57gat), .B(G85gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n380), .B(new_n381), .ZN(new_n382));
  NAND4_X1  g181(.A1(new_n349), .A2(new_n281), .A3(new_n352), .A4(new_n284), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT4), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n220), .A2(KEYINPUT4), .A3(new_n331), .ZN(new_n386));
  AND2_X1   g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT5), .ZN(new_n388));
  NAND2_X1  g187(.A1(G225gat), .A2(G233gat), .ZN(new_n389));
  OAI21_X1  g188(.A(KEYINPUT3), .B1(new_n324), .B2(new_n330), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n353), .A2(new_n390), .A3(new_n285), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n387), .A2(new_n388), .A3(new_n389), .A4(new_n391), .ZN(new_n392));
  NAND4_X1  g191(.A1(new_n391), .A2(new_n385), .A3(new_n386), .A4(new_n389), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n359), .A2(new_n285), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(new_n383), .ZN(new_n395));
  INV_X1    g194(.A(new_n389), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n393), .A2(KEYINPUT5), .A3(new_n397), .ZN(new_n398));
  AOI211_X1 g197(.A(new_n378), .B(new_n382), .C1(new_n392), .C2(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n392), .A2(new_n398), .A3(new_n382), .ZN(new_n400));
  AND2_X1   g199(.A1(new_n400), .A2(new_n378), .ZN(new_n401));
  INV_X1    g200(.A(new_n382), .ZN(new_n402));
  INV_X1    g201(.A(new_n398), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n393), .A2(KEYINPUT5), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n402), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n399), .B1(new_n401), .B2(new_n405), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n377), .A2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT74), .ZN(new_n408));
  AOI21_X1  g207(.A(KEYINPUT29), .B1(new_n280), .B2(new_n288), .ZN(new_n409));
  NAND2_X1  g208(.A1(G226gat), .A2(G233gat), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(KEYINPUT72), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT72), .ZN(new_n413));
  AOI22_X1  g212(.A1(new_n275), .A2(new_n279), .B1(new_n286), .B2(new_n287), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n413), .B(new_n410), .C1(new_n414), .C2(KEYINPUT29), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n410), .B1(new_n280), .B2(new_n288), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n416), .A2(new_n357), .ZN(new_n417));
  AND3_X1   g216(.A1(new_n412), .A2(new_n415), .A3(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT71), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n343), .B1(new_n252), .B2(new_n269), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n416), .B1(new_n420), .B2(new_n410), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n419), .B1(new_n421), .B2(new_n342), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n410), .B1(new_n414), .B2(KEYINPUT29), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n411), .B1(new_n252), .B2(new_n269), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n425), .A2(KEYINPUT71), .A3(new_n357), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n418), .B1(new_n422), .B2(new_n426), .ZN(new_n427));
  XOR2_X1   g226(.A(G8gat), .B(G36gat), .Z(new_n428));
  XNOR2_X1  g227(.A(new_n428), .B(KEYINPUT73), .ZN(new_n429));
  XNOR2_X1  g228(.A(G64gat), .B(G92gat), .ZN(new_n430));
  XOR2_X1   g229(.A(new_n429), .B(new_n430), .Z(new_n431));
  OAI21_X1  g230(.A(new_n408), .B1(new_n427), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n422), .A2(new_n426), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n412), .A2(new_n415), .A3(new_n417), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n431), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n435), .A2(KEYINPUT74), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n432), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT30), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n427), .A2(new_n439), .A3(new_n431), .ZN(new_n440));
  AOI21_X1  g239(.A(KEYINPUT71), .B1(new_n425), .B2(new_n357), .ZN(new_n441));
  AOI211_X1 g240(.A(new_n419), .B(new_n342), .C1(new_n423), .C2(new_n424), .ZN(new_n442));
  OAI211_X1 g241(.A(new_n434), .B(new_n431), .C1(new_n441), .C2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(KEYINPUT30), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n440), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n407), .A2(new_n438), .A3(new_n445), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n202), .B1(new_n315), .B2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT87), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n400), .A2(new_n378), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT77), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n400), .A2(KEYINPUT77), .A3(new_n378), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n451), .A2(new_n405), .A3(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n399), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n438), .A2(new_n455), .A3(new_n445), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n374), .A2(new_n376), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n307), .A2(new_n310), .ZN(new_n459));
  INV_X1    g258(.A(new_n297), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n307), .A2(new_n297), .A3(new_n310), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n458), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  OAI211_X1 g262(.A(new_n448), .B(KEYINPUT35), .C1(new_n456), .C2(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n461), .A2(KEYINPUT70), .A3(new_n462), .ZN(new_n465));
  INV_X1    g264(.A(new_n311), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AOI22_X1  g266(.A1(new_n432), .A2(new_n437), .B1(new_n440), .B2(new_n444), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n467), .A2(KEYINPUT86), .A3(new_n468), .A4(new_n407), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n447), .A2(new_n464), .A3(new_n469), .ZN(new_n470));
  NOR3_X1   g269(.A1(new_n312), .A2(new_n313), .A3(new_n457), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n471), .A2(new_n468), .A3(new_n455), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n448), .B1(new_n472), .B2(KEYINPUT35), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n395), .A2(new_n396), .ZN(new_n474));
  XNOR2_X1  g273(.A(new_n474), .B(KEYINPUT81), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n387), .A2(new_n391), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(new_n396), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n475), .A2(KEYINPUT39), .A3(new_n477), .ZN(new_n478));
  XNOR2_X1  g277(.A(KEYINPUT80), .B(KEYINPUT39), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n476), .A2(new_n396), .A3(new_n479), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n478), .A2(new_n382), .A3(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT82), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n482), .A2(KEYINPUT40), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n483), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n478), .A2(new_n382), .A3(new_n485), .A4(new_n480), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n484), .A2(new_n405), .A3(new_n486), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n458), .B1(new_n468), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n405), .A2(new_n378), .A3(new_n400), .ZN(new_n489));
  AND3_X1   g288(.A1(new_n489), .A2(new_n443), .A3(new_n454), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT84), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n441), .A2(new_n442), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT37), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n434), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n491), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n433), .A2(KEYINPUT84), .A3(new_n493), .A4(new_n434), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n495), .A2(new_n496), .A3(new_n436), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n412), .A2(new_n357), .A3(new_n424), .A4(new_n415), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n425), .A2(new_n342), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n498), .A2(new_n499), .A3(KEYINPUT37), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT83), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT38), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n498), .A2(new_n499), .A3(KEYINPUT83), .A4(KEYINPUT37), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n502), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n490), .B1(new_n497), .B2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT85), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n435), .A2(KEYINPUT37), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n508), .A2(new_n496), .A3(new_n495), .A4(new_n436), .ZN(new_n509));
  AOI22_X1  g308(.A1(new_n506), .A2(new_n507), .B1(KEYINPUT38), .B2(new_n509), .ZN(new_n510));
  OAI211_X1 g309(.A(KEYINPUT85), .B(new_n490), .C1(new_n497), .C2(new_n505), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n488), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT36), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n467), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n456), .A2(new_n457), .ZN(new_n515));
  OAI21_X1  g314(.A(KEYINPUT36), .B1(new_n312), .B2(new_n313), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  OAI22_X1  g316(.A1(new_n470), .A2(new_n473), .B1(new_n512), .B2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT18), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT91), .ZN(new_n521));
  XNOR2_X1  g320(.A(G15gat), .B(G22gat), .ZN(new_n522));
  OR2_X1    g321(.A1(new_n522), .A2(G1gat), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT89), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT16), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n522), .B1(new_n526), .B2(G1gat), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n523), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n525), .A2(new_n528), .A3(G8gat), .ZN(new_n529));
  INV_X1    g328(.A(G8gat), .ZN(new_n530));
  OAI211_X1 g329(.A(new_n523), .B(new_n527), .C1(new_n524), .C2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT90), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n532), .B(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT14), .ZN(new_n535));
  INV_X1    g334(.A(G29gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n538));
  AOI21_X1  g337(.A(G36gat), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(G36gat), .ZN(new_n540));
  NOR3_X1   g339(.A1(new_n535), .A2(new_n540), .A3(G29gat), .ZN(new_n541));
  OR3_X1    g340(.A1(new_n539), .A2(KEYINPUT15), .A3(new_n541), .ZN(new_n542));
  OAI21_X1  g341(.A(KEYINPUT15), .B1(new_n539), .B2(new_n541), .ZN(new_n543));
  XNOR2_X1  g342(.A(G43gat), .B(G50gat), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  OR2_X1    g344(.A1(new_n543), .A2(new_n544), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT88), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n545), .A2(new_n546), .A3(KEYINPUT88), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n521), .B1(new_n534), .B2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n551), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n532), .B(KEYINPUT90), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n553), .A2(new_n554), .A3(KEYINPUT91), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT17), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n551), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n547), .A2(KEYINPUT17), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n532), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n556), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(G229gat), .A2(G233gat), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n520), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n553), .A2(new_n554), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n567), .B1(new_n552), .B2(new_n555), .ZN(new_n568));
  XOR2_X1   g367(.A(new_n564), .B(KEYINPUT13), .Z(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  OR2_X1    g369(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n556), .A2(new_n562), .A3(KEYINPUT18), .A4(new_n564), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n566), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(G113gat), .B(G141gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(G197gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(KEYINPUT11), .B(G169gat), .ZN(new_n576));
  XOR2_X1   g375(.A(new_n575), .B(new_n576), .Z(new_n577));
  XOR2_X1   g376(.A(new_n577), .B(KEYINPUT12), .Z(new_n578));
  NAND2_X1  g377(.A1(new_n573), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n578), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n566), .A2(new_n571), .A3(new_n580), .A4(new_n572), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(G190gat), .B(G218gat), .ZN(new_n584));
  NAND2_X1  g383(.A1(G85gat), .A2(G92gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(KEYINPUT7), .ZN(new_n586));
  NAND2_X1  g385(.A1(G99gat), .A2(G106gat), .ZN(new_n587));
  INV_X1    g386(.A(G85gat), .ZN(new_n588));
  INV_X1    g387(.A(G92gat), .ZN(new_n589));
  AOI22_X1  g388(.A1(KEYINPUT8), .A2(new_n587), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n586), .A2(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(G99gat), .B(G106gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n591), .B(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n593), .B1(new_n558), .B2(new_n559), .ZN(new_n594));
  NAND2_X1  g393(.A1(G232gat), .A2(G233gat), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(KEYINPUT41), .ZN(new_n597));
  XOR2_X1   g396(.A(new_n591), .B(new_n592), .Z(new_n598));
  OAI21_X1  g397(.A(new_n597), .B1(new_n551), .B2(new_n598), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n584), .B1(new_n594), .B2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  OR2_X1    g400(.A1(new_n601), .A2(KEYINPUT94), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n596), .A2(KEYINPUT41), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(G134gat), .ZN(new_n604));
  INV_X1    g403(.A(G162gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n594), .ZN(new_n607));
  INV_X1    g406(.A(new_n584), .ZN(new_n608));
  INV_X1    g407(.A(new_n599), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n607), .A2(KEYINPUT93), .A3(new_n608), .A4(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT93), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n611), .A2(new_n612), .A3(new_n600), .ZN(new_n613));
  NAND4_X1  g412(.A1(new_n602), .A2(new_n606), .A3(new_n610), .A4(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n610), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n606), .B1(new_n601), .B2(KEYINPUT94), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT92), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n619), .A2(G57gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(G64gat), .ZN(new_n621));
  NAND2_X1  g420(.A1(G71gat), .A2(G78gat), .ZN(new_n622));
  OR2_X1    g421(.A1(G71gat), .A2(G78gat), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT9), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n622), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n621), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g425(.A(KEYINPUT9), .B1(G57gat), .B2(G64gat), .ZN(new_n627));
  AND2_X1   g426(.A1(G57gat), .A2(G64gat), .ZN(new_n628));
  OAI211_X1 g427(.A(new_n622), .B(new_n623), .C1(new_n627), .C2(new_n628), .ZN(new_n629));
  AND2_X1   g428(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n630), .A2(KEYINPUT21), .ZN(new_n631));
  AND2_X1   g430(.A1(G231gat), .A2(G233gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(G127gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n554), .B1(KEYINPUT21), .B2(new_n630), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(G155gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(G183gat), .B(G211gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n637), .B(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n618), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT97), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT95), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n591), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(new_n598), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT10), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n593), .A2(new_n630), .A3(new_n646), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n648), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n593), .A2(KEYINPUT10), .A3(new_n630), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(G230gat), .A2(G233gat), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n644), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n648), .A2(new_n650), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n657), .A2(G230gat), .A3(G233gat), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n653), .A2(new_n644), .A3(new_n654), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n656), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(G120gat), .B(G148gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(G176gat), .B(G204gat), .ZN(new_n662));
  XOR2_X1   g461(.A(new_n661), .B(new_n662), .Z(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n660), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT98), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT96), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n653), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n651), .A2(KEYINPUT96), .A3(new_n652), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n668), .A2(new_n654), .A3(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n670), .A2(new_n658), .A3(new_n663), .ZN(new_n671));
  AND3_X1   g470(.A1(new_n665), .A2(new_n666), .A3(new_n671), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n666), .B1(new_n665), .B2(new_n671), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n643), .A2(new_n674), .ZN(new_n675));
  NOR3_X1   g474(.A1(new_n519), .A2(new_n583), .A3(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n455), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(G1gat), .ZN(G1324gat));
  INV_X1    g478(.A(new_n468), .ZN(new_n680));
  XOR2_X1   g479(.A(KEYINPUT16), .B(G8gat), .Z(new_n681));
  AND3_X1   g480(.A1(new_n676), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n530), .B1(new_n676), .B2(new_n680), .ZN(new_n683));
  OAI21_X1  g482(.A(KEYINPUT42), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n684), .B1(KEYINPUT42), .B2(new_n682), .ZN(G1325gat));
  INV_X1    g484(.A(G15gat), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n676), .A2(new_n686), .A3(new_n467), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n514), .A2(new_n516), .ZN(new_n688));
  AND2_X1   g487(.A1(new_n676), .A2(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n687), .B1(new_n689), .B2(new_n686), .ZN(G1326gat));
  NAND2_X1  g489(.A1(new_n676), .A2(new_n457), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(KEYINPUT99), .ZN(new_n692));
  XOR2_X1   g491(.A(KEYINPUT43), .B(G22gat), .Z(new_n693));
  XNOR2_X1  g492(.A(new_n692), .B(new_n693), .ZN(G1327gat));
  NAND2_X1  g493(.A1(new_n518), .A2(new_n618), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n518), .A2(KEYINPUT44), .A3(new_n618), .ZN(new_n698));
  AND2_X1   g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n642), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n665), .A2(new_n671), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(KEYINPUT98), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n665), .A2(new_n666), .A3(new_n671), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n583), .A2(new_n700), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n699), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(G29gat), .B1(new_n706), .B2(new_n455), .ZN(new_n707));
  AND3_X1   g506(.A1(new_n518), .A2(new_n618), .A3(new_n705), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n708), .A2(new_n536), .A3(new_n677), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT45), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n707), .A2(new_n710), .ZN(G1328gat));
  NAND3_X1  g510(.A1(new_n708), .A2(new_n540), .A3(new_n680), .ZN(new_n712));
  XOR2_X1   g511(.A(new_n712), .B(KEYINPUT46), .Z(new_n713));
  OAI21_X1  g512(.A(G36gat), .B1(new_n706), .B2(new_n468), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(G1329gat));
  INV_X1    g514(.A(G43gat), .ZN(new_n716));
  INV_X1    g515(.A(new_n706), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(new_n688), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n716), .B1(new_n718), .B2(KEYINPUT100), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n719), .B1(KEYINPUT100), .B2(new_n718), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n708), .A2(new_n716), .A3(new_n467), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n720), .A2(KEYINPUT47), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n718), .A2(G43gat), .ZN(new_n723));
  AND2_X1   g522(.A1(new_n723), .A2(new_n721), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n722), .B1(KEYINPUT47), .B2(new_n724), .ZN(G1330gat));
  INV_X1    g524(.A(KEYINPUT48), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n717), .A2(new_n457), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(G50gat), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n726), .B1(new_n728), .B2(KEYINPUT102), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n457), .A2(new_n369), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(KEYINPUT101), .ZN(new_n731));
  AOI22_X1  g530(.A1(new_n727), .A2(G50gat), .B1(new_n708), .B2(new_n731), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n729), .B(new_n732), .ZN(G1331gat));
  AND4_X1   g532(.A1(new_n518), .A2(new_n583), .A3(new_n643), .A4(new_n704), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(new_n677), .ZN(new_n735));
  XNOR2_X1  g534(.A(KEYINPUT103), .B(G57gat), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n735), .B(new_n736), .ZN(G1332gat));
  NAND2_X1  g536(.A1(new_n734), .A2(new_n680), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n738), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n739));
  XOR2_X1   g538(.A(KEYINPUT49), .B(G64gat), .Z(new_n740));
  OAI21_X1  g539(.A(new_n739), .B1(new_n738), .B2(new_n740), .ZN(G1333gat));
  INV_X1    g540(.A(G71gat), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n734), .A2(new_n742), .A3(new_n467), .ZN(new_n743));
  AND2_X1   g542(.A1(new_n734), .A2(new_n688), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n743), .B1(new_n744), .B2(new_n742), .ZN(new_n745));
  XOR2_X1   g544(.A(new_n745), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g545(.A1(new_n734), .A2(new_n457), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g547(.A1(new_n700), .A2(new_n582), .A3(new_n674), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(KEYINPUT104), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n697), .A2(new_n698), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(KEYINPUT105), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT105), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n697), .A2(new_n753), .A3(new_n698), .A4(new_n750), .ZN(new_n754));
  AND2_X1   g553(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  OAI21_X1  g555(.A(G85gat), .B1(new_n756), .B2(new_n455), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n518), .A2(new_n583), .A3(new_n642), .A4(new_n618), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT51), .ZN(new_n759));
  OR2_X1    g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT106), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n758), .A2(new_n759), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n760), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n758), .A2(KEYINPUT106), .A3(new_n759), .ZN(new_n764));
  NOR3_X1   g563(.A1(new_n674), .A2(G85gat), .A3(new_n455), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n763), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n757), .A2(new_n766), .ZN(G1336gat));
  INV_X1    g566(.A(KEYINPUT52), .ZN(new_n768));
  NOR3_X1   g567(.A1(new_n674), .A2(G92gat), .A3(new_n468), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n763), .A2(new_n764), .A3(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT108), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n771), .B1(new_n751), .B2(new_n468), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(G92gat), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n751), .A2(new_n771), .A3(new_n468), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n768), .B(new_n770), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n589), .B1(new_n755), .B2(new_n680), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT107), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n760), .A2(new_n777), .A3(new_n762), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n758), .A2(KEYINPUT107), .A3(new_n759), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n776), .B1(new_n769), .B2(new_n780), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n775), .B1(new_n781), .B2(new_n768), .ZN(G1337gat));
  INV_X1    g581(.A(new_n688), .ZN(new_n783));
  OAI21_X1  g582(.A(G99gat), .B1(new_n756), .B2(new_n783), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n674), .A2(new_n315), .A3(G99gat), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n763), .A2(new_n764), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n784), .A2(new_n786), .ZN(G1338gat));
  NOR3_X1   g586(.A1(new_n674), .A2(G106gat), .A3(new_n458), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n763), .A2(new_n764), .A3(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT53), .ZN(new_n790));
  OAI21_X1  g589(.A(G106gat), .B1(new_n751), .B2(new_n458), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n789), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT110), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n752), .A2(new_n457), .A3(new_n754), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(G106gat), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT109), .ZN(new_n796));
  AOI22_X1  g595(.A1(new_n795), .A2(new_n796), .B1(new_n780), .B2(new_n788), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n794), .A2(KEYINPUT109), .A3(G106gat), .ZN(new_n798));
  AOI211_X1 g597(.A(new_n793), .B(new_n790), .C1(new_n797), .C2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n795), .A2(new_n796), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n780), .A2(new_n788), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n800), .A2(new_n798), .A3(new_n801), .ZN(new_n802));
  AOI21_X1  g601(.A(KEYINPUT110), .B1(new_n802), .B2(KEYINPUT53), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n792), .B1(new_n799), .B2(new_n803), .ZN(G1339gat));
  NOR2_X1   g603(.A1(new_n680), .A2(new_n455), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n675), .A2(new_n582), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT111), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n653), .A2(new_n654), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT54), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(new_n670), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(KEYINPUT112), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT112), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n811), .A2(new_n670), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(KEYINPUT54), .B1(new_n656), .B2(new_n659), .ZN(new_n817));
  OAI21_X1  g616(.A(KEYINPUT113), .B1(new_n817), .B2(new_n663), .ZN(new_n818));
  INV_X1    g617(.A(new_n659), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n810), .B1(new_n819), .B2(new_n655), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT113), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n820), .A2(new_n821), .A3(new_n664), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n816), .A2(new_n818), .A3(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT55), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n816), .A2(new_n818), .A3(KEYINPUT55), .A4(new_n822), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n825), .A2(new_n671), .A3(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT114), .ZN(new_n828));
  AOI22_X1  g627(.A1(new_n563), .A2(new_n565), .B1(new_n568), .B2(new_n570), .ZN(new_n829));
  INV_X1    g628(.A(new_n577), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n828), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n568), .A2(new_n570), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n564), .B1(new_n556), .B2(new_n562), .ZN(new_n833));
  OAI211_X1 g632(.A(KEYINPUT114), .B(new_n577), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  AND2_X1   g633(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n835), .A2(new_n618), .A3(new_n581), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n827), .A2(new_n836), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n825), .A2(new_n582), .A3(new_n671), .A4(new_n826), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT115), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n835), .A2(new_n704), .A3(new_n839), .A4(new_n581), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n831), .A2(new_n581), .A3(new_n834), .ZN(new_n841));
  OAI21_X1  g640(.A(KEYINPUT115), .B1(new_n674), .B2(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n838), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(new_n618), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n837), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT116), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n642), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  AOI211_X1 g646(.A(KEYINPUT116), .B(new_n837), .C1(new_n844), .C2(new_n843), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n808), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  AND3_X1   g648(.A1(new_n849), .A2(KEYINPUT117), .A3(new_n458), .ZN(new_n850));
  AOI21_X1  g649(.A(KEYINPUT117), .B1(new_n849), .B2(new_n458), .ZN(new_n851));
  OAI211_X1 g650(.A(new_n467), .B(new_n805), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  OAI21_X1  g651(.A(G113gat), .B1(new_n852), .B2(new_n583), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n849), .A2(new_n677), .ZN(new_n854));
  AND3_X1   g653(.A1(new_n854), .A2(new_n468), .A3(new_n471), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n583), .A2(new_n213), .A3(new_n214), .ZN(new_n856));
  XOR2_X1   g655(.A(new_n856), .B(KEYINPUT118), .Z(new_n857));
  NAND2_X1  g656(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n853), .A2(new_n858), .ZN(G1340gat));
  NOR3_X1   g658(.A1(new_n852), .A2(new_n208), .A3(new_n674), .ZN(new_n860));
  AOI21_X1  g659(.A(G120gat), .B1(new_n855), .B2(new_n704), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n860), .A2(new_n861), .ZN(G1341gat));
  OAI21_X1  g661(.A(new_n205), .B1(new_n852), .B2(new_n642), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n855), .A2(new_n283), .A3(new_n700), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT119), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n863), .A2(KEYINPUT119), .A3(new_n864), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(G1342gat));
  NOR2_X1   g668(.A1(new_n844), .A2(new_n680), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n854), .A2(new_n282), .A3(new_n471), .A4(new_n870), .ZN(new_n871));
  XOR2_X1   g670(.A(new_n871), .B(KEYINPUT56), .Z(new_n872));
  OAI21_X1  g671(.A(G134gat), .B1(new_n852), .B2(new_n844), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(G1343gat));
  NOR2_X1   g673(.A1(new_n688), .A2(new_n458), .ZN(new_n875));
  AND3_X1   g674(.A1(new_n854), .A2(new_n468), .A3(new_n875), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n876), .A2(new_n320), .A3(new_n582), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n783), .A2(new_n805), .ZN(new_n878));
  XOR2_X1   g677(.A(new_n878), .B(KEYINPUT120), .Z(new_n879));
  AOI21_X1  g678(.A(KEYINPUT57), .B1(new_n849), .B2(new_n457), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT57), .ZN(new_n881));
  OAI21_X1  g680(.A(KEYINPUT121), .B1(new_n674), .B2(new_n841), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n838), .A2(new_n882), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n674), .A2(new_n841), .A3(KEYINPUT121), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n844), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(new_n837), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n700), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(new_n887), .ZN(new_n888));
  AOI211_X1 g687(.A(new_n881), .B(new_n458), .C1(new_n888), .C2(new_n808), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n879), .B1(new_n880), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(G141gat), .B1(new_n890), .B2(new_n583), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n877), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(KEYINPUT58), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT58), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n877), .A2(new_n891), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n893), .A2(new_n895), .ZN(G1344gat));
  NAND2_X1  g695(.A1(new_n876), .A2(new_n704), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(KEYINPUT59), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n898), .A2(new_n317), .A3(new_n318), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n849), .A2(KEYINPUT57), .A3(new_n457), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n457), .B1(new_n887), .B2(new_n806), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(new_n881), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n903), .A2(new_n704), .A3(new_n879), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n904), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n905));
  OR3_X1    g704(.A1(new_n890), .A2(KEYINPUT59), .A3(new_n674), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n899), .A2(new_n905), .A3(new_n906), .ZN(G1345gat));
  INV_X1    g706(.A(G155gat), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n876), .A2(new_n908), .A3(new_n700), .ZN(new_n909));
  OAI21_X1  g708(.A(G155gat), .B1(new_n890), .B2(new_n642), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(G1346gat));
  OAI21_X1  g710(.A(G162gat), .B1(new_n890), .B2(new_n844), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n854), .A2(new_n605), .A3(new_n870), .A4(new_n875), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(G1347gat));
  NOR2_X1   g713(.A1(new_n468), .A2(new_n677), .ZN(new_n915));
  AND3_X1   g714(.A1(new_n849), .A2(new_n471), .A3(new_n915), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n916), .A2(new_n223), .A3(new_n582), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n849), .A2(new_n458), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT117), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n849), .A2(KEYINPUT117), .A3(new_n458), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND4_X1  g721(.A1(new_n922), .A2(new_n467), .A3(new_n582), .A4(new_n915), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n923), .A2(KEYINPUT122), .A3(G169gat), .ZN(new_n924));
  INV_X1    g723(.A(new_n924), .ZN(new_n925));
  AOI21_X1  g724(.A(KEYINPUT122), .B1(new_n923), .B2(G169gat), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n917), .B1(new_n925), .B2(new_n926), .ZN(G1348gat));
  OAI211_X1 g726(.A(new_n467), .B(new_n915), .C1(new_n850), .C2(new_n851), .ZN(new_n928));
  OAI21_X1  g727(.A(G176gat), .B1(new_n928), .B2(new_n674), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n916), .A2(new_n224), .A3(new_n704), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(G1349gat));
  OAI21_X1  g730(.A(G183gat), .B1(new_n928), .B2(new_n642), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT123), .ZN(new_n933));
  AND3_X1   g732(.A1(new_n700), .A2(new_n259), .A3(new_n263), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n933), .B1(new_n916), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n932), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(KEYINPUT60), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT60), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n932), .A2(new_n938), .A3(new_n935), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n937), .A2(new_n939), .ZN(G1350gat));
  NAND3_X1  g739(.A1(new_n916), .A2(new_n242), .A3(new_n618), .ZN(new_n941));
  NAND4_X1  g740(.A1(new_n922), .A2(new_n467), .A3(new_n618), .A4(new_n915), .ZN(new_n942));
  NOR2_X1   g741(.A1(KEYINPUT124), .A2(KEYINPUT61), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n242), .B1(KEYINPUT124), .B2(KEYINPUT61), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  INV_X1    g744(.A(new_n945), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n943), .B1(new_n942), .B2(new_n944), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n941), .B1(new_n946), .B2(new_n947), .ZN(G1351gat));
  AND4_X1   g747(.A1(new_n457), .A2(new_n849), .A3(new_n783), .A4(new_n915), .ZN(new_n949));
  AOI21_X1  g748(.A(G197gat), .B1(new_n949), .B2(new_n582), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n783), .A2(new_n915), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n951), .B1(new_n900), .B2(new_n902), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n582), .A2(G197gat), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n950), .B1(new_n952), .B2(new_n953), .ZN(G1352gat));
  XOR2_X1   g753(.A(KEYINPUT125), .B(G204gat), .Z(new_n955));
  NAND3_X1  g754(.A1(new_n949), .A2(new_n704), .A3(new_n955), .ZN(new_n956));
  OR2_X1    g755(.A1(new_n956), .A2(KEYINPUT62), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(KEYINPUT62), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n952), .A2(new_n704), .ZN(new_n959));
  OAI211_X1 g758(.A(new_n957), .B(new_n958), .C1(new_n955), .C2(new_n959), .ZN(G1353gat));
  NAND3_X1  g759(.A1(new_n949), .A2(new_n334), .A3(new_n700), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n952), .A2(new_n700), .ZN(new_n962));
  AND3_X1   g761(.A1(new_n962), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n963));
  AOI21_X1  g762(.A(KEYINPUT63), .B1(new_n962), .B2(G211gat), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n961), .B1(new_n963), .B2(new_n964), .ZN(G1354gat));
  AOI21_X1  g764(.A(G218gat), .B1(new_n949), .B2(new_n618), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT126), .ZN(new_n967));
  OR2_X1    g766(.A1(new_n952), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n618), .A2(G218gat), .ZN(new_n969));
  XOR2_X1   g768(.A(new_n969), .B(KEYINPUT127), .Z(new_n970));
  AOI21_X1  g769(.A(new_n970), .B1(new_n952), .B2(new_n967), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n966), .B1(new_n968), .B2(new_n971), .ZN(G1355gat));
endmodule


