//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 1 0 1 0 0 0 1 0 0 1 0 0 1 0 0 1 1 1 1 1 0 0 0 1 0 1 0 1 1 1 1 1 1 1 1 0 0 0 0 0 1 0 0 0 0 1 1 0 0 1 0 1 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:39 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1250, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  NOR3_X1   g0006(.A1(new_n206), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0007(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0008(.A1(new_n206), .A2(G50), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(KEYINPUT65), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND3_X1  g0012(.A1(KEYINPUT65), .A2(G1), .A3(G13), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(G20), .ZN(new_n215));
  INV_X1    g0015(.A(G1), .ZN(new_n216));
  INV_X1    g0016(.A(G20), .ZN(new_n217));
  NOR3_X1   g0017(.A1(new_n216), .A2(new_n217), .A3(G13), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n218), .B(G250), .C1(G257), .C2(G264), .ZN(new_n219));
  INV_X1    g0019(.A(KEYINPUT0), .ZN(new_n220));
  OAI22_X1  g0020(.A1(new_n209), .A2(new_n215), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G77), .A2(G244), .B1(G87), .B2(G250), .ZN(new_n222));
  INV_X1    g0022(.A(G116), .ZN(new_n223));
  INV_X1    g0023(.A(G270), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n222), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n226));
  INV_X1    g0026(.A(G50), .ZN(new_n227));
  INV_X1    g0027(.A(G226), .ZN(new_n228));
  INV_X1    g0028(.A(G238), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n226), .B1(new_n227), .B2(new_n228), .C1(new_n202), .C2(new_n229), .ZN(new_n230));
  AOI211_X1 g0030(.A(new_n225), .B(new_n230), .C1(G97), .C2(G257), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(G1), .B2(G20), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n232), .B(KEYINPUT1), .Z(new_n233));
  AOI211_X1 g0033(.A(new_n221), .B(new_n233), .C1(new_n220), .C2(new_n219), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n236), .B(new_n237), .Z(new_n238));
  XOR2_X1   g0038(.A(G250), .B(G257), .Z(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G358));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  NAND3_X1  g0049(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n212), .A2(new_n213), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(KEYINPUT69), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT69), .ZN(new_n253));
  NAND4_X1  g0053(.A1(new_n212), .A2(new_n253), .A3(new_n213), .A4(new_n250), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n255), .B1(new_n216), .B2(G20), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G50), .ZN(new_n257));
  INV_X1    g0057(.A(G13), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(G1), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G20), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(new_n227), .ZN(new_n262));
  OAI21_X1  g0062(.A(G20), .B1(new_n206), .B2(G50), .ZN(new_n263));
  NOR2_X1   g0063(.A1(G20), .A2(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G150), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n217), .A2(G33), .ZN(new_n266));
  OR2_X1    g0066(.A1(KEYINPUT8), .A2(G58), .ZN(new_n267));
  NAND2_X1  g0067(.A1(KEYINPUT8), .A2(G58), .ZN(new_n268));
  AND2_X1   g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  OAI211_X1 g0070(.A(new_n263), .B(new_n265), .C1(new_n266), .C2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(new_n255), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n257), .A2(new_n262), .A3(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(KEYINPUT9), .ZN(new_n275));
  XNOR2_X1  g0075(.A(KEYINPUT3), .B(G33), .ZN(new_n276));
  AOI21_X1  g0076(.A(KEYINPUT67), .B1(new_n276), .B2(G1698), .ZN(new_n277));
  AND2_X1   g0077(.A1(KEYINPUT3), .A2(G33), .ZN(new_n278));
  NOR2_X1   g0078(.A1(KEYINPUT3), .A2(G33), .ZN(new_n279));
  OAI211_X1 g0079(.A(KEYINPUT67), .B(G1698), .C1(new_n278), .C2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  OAI21_X1  g0081(.A(G223), .B1(new_n277), .B2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n276), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G77), .ZN(new_n284));
  INV_X1    g0084(.A(G1698), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n276), .A2(G222), .A3(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n282), .A2(new_n284), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(KEYINPUT68), .ZN(new_n288));
  NAND2_X1  g0088(.A1(G33), .A2(G41), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n214), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT68), .ZN(new_n292));
  NAND4_X1  g0092(.A1(new_n282), .A2(new_n292), .A3(new_n284), .A4(new_n286), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n288), .A2(new_n291), .A3(new_n293), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n216), .B1(G41), .B2(G45), .ZN(new_n295));
  INV_X1    g0095(.A(G274), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n289), .A2(G1), .A3(G13), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(new_n295), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  OR2_X1    g0101(.A1(KEYINPUT66), .A2(G226), .ZN(new_n302));
  NAND2_X1  g0102(.A1(KEYINPUT66), .A2(G226), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n301), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n294), .A2(G190), .A3(new_n298), .A4(new_n304), .ZN(new_n305));
  AND2_X1   g0105(.A1(new_n275), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT10), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT9), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n273), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n294), .A2(new_n298), .A3(new_n304), .ZN(new_n310));
  XNOR2_X1  g0110(.A(KEYINPUT71), .B(G200), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n306), .A2(new_n307), .A3(new_n309), .A4(new_n312), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n312), .A2(new_n309), .A3(new_n305), .A4(new_n275), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(KEYINPUT10), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(G169), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n310), .A2(new_n317), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n310), .A2(G179), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n319), .A2(KEYINPUT70), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT70), .ZN(new_n321));
  NOR3_X1   g0121(.A1(new_n310), .A2(new_n321), .A3(G179), .ZN(new_n322));
  OAI211_X1 g0122(.A(new_n273), .B(new_n318), .C1(new_n320), .C2(new_n322), .ZN(new_n323));
  OAI21_X1  g0123(.A(G238), .B1(new_n277), .B2(new_n281), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n276), .A2(G232), .A3(new_n285), .ZN(new_n325));
  INV_X1    g0125(.A(G107), .ZN(new_n326));
  OAI211_X1 g0126(.A(new_n324), .B(new_n325), .C1(new_n326), .C2(new_n276), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n297), .B1(new_n327), .B2(new_n291), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n301), .A2(G244), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(G179), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n330), .A2(new_n317), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n256), .A2(G77), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n269), .A2(new_n264), .ZN(new_n336));
  XNOR2_X1  g0136(.A(KEYINPUT15), .B(G87), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n336), .B1(new_n266), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(G77), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n217), .A2(new_n339), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n255), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n335), .B(new_n341), .C1(G77), .C2(new_n260), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n333), .A2(new_n334), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n342), .B1(new_n331), .B2(G190), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n330), .A2(new_n311), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n316), .A2(new_n323), .A3(new_n343), .A4(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT72), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n276), .A2(G226), .A3(new_n285), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n276), .A2(G232), .A3(G1698), .ZN(new_n351));
  NAND2_X1  g0151(.A1(G33), .A2(G97), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n350), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n297), .B1(new_n353), .B2(new_n291), .ZN(new_n354));
  XOR2_X1   g0154(.A(KEYINPUT73), .B(KEYINPUT13), .Z(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n301), .A2(G238), .ZN(new_n357));
  AND3_X1   g0157(.A1(new_n354), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n356), .B1(new_n354), .B2(new_n357), .ZN(new_n359));
  OAI21_X1  g0159(.A(G169), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT14), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n354), .A2(new_n357), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n355), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n354), .A2(new_n356), .A3(new_n357), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n366), .A2(KEYINPUT14), .A3(G169), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n362), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n363), .A2(KEYINPUT13), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n369), .A2(G179), .A3(new_n365), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT74), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n369), .A2(KEYINPUT74), .A3(G179), .A4(new_n365), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n368), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n256), .A2(G68), .ZN(new_n376));
  INV_X1    g0176(.A(new_n266), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n377), .A2(G77), .B1(new_n264), .B2(G50), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n378), .B1(new_n217), .B2(G68), .ZN(new_n379));
  AND2_X1   g0179(.A1(new_n379), .A2(new_n255), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n376), .B1(KEYINPUT11), .B2(new_n380), .ZN(new_n381));
  AND2_X1   g0181(.A1(new_n380), .A2(KEYINPUT11), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n259), .A2(G20), .A3(new_n202), .ZN(new_n383));
  XOR2_X1   g0183(.A(new_n383), .B(KEYINPUT12), .Z(new_n384));
  NOR3_X1   g0184(.A1(new_n381), .A2(new_n382), .A3(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n375), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n366), .A2(G200), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n369), .A2(G190), .A3(new_n365), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n385), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n387), .A2(new_n390), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n349), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n228), .A2(G1698), .ZN(new_n393));
  OAI211_X1 g0193(.A(new_n276), .B(new_n393), .C1(G223), .C2(G1698), .ZN(new_n394));
  NAND2_X1  g0194(.A1(G33), .A2(G87), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(new_n291), .ZN(new_n397));
  INV_X1    g0197(.A(G190), .ZN(new_n398));
  AND3_X1   g0198(.A1(new_n299), .A2(G232), .A3(new_n295), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n397), .A2(new_n398), .A3(new_n298), .A4(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n290), .B1(new_n394), .B2(new_n395), .ZN(new_n402));
  NOR3_X1   g0202(.A1(new_n402), .A2(new_n297), .A3(new_n399), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n401), .B1(new_n403), .B2(G200), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n255), .A2(new_n261), .ZN(new_n405));
  OAI211_X1 g0205(.A(new_n267), .B(new_n268), .C1(G1), .C2(new_n217), .ZN(new_n406));
  XNOR2_X1  g0206(.A(new_n406), .B(KEYINPUT77), .ZN(new_n407));
  AOI22_X1  g0207(.A1(new_n405), .A2(new_n407), .B1(new_n261), .B2(new_n270), .ZN(new_n408));
  NAND2_X1  g0208(.A1(G58), .A2(G68), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n203), .A2(new_n205), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(G20), .ZN(new_n411));
  INV_X1    g0211(.A(G159), .ZN(new_n412));
  NOR3_X1   g0212(.A1(new_n412), .A2(G20), .A3(G33), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n411), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(KEYINPUT75), .ZN(new_n416));
  OR2_X1    g0216(.A1(KEYINPUT3), .A2(G33), .ZN(new_n417));
  NAND2_X1  g0217(.A1(KEYINPUT3), .A2(G33), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n417), .A2(new_n217), .A3(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT7), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n417), .A2(KEYINPUT7), .A3(new_n217), .A4(new_n418), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(G68), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT75), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n411), .A2(new_n425), .A3(new_n414), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n416), .A2(KEYINPUT16), .A3(new_n424), .A4(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(new_n255), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n425), .B1(new_n411), .B2(new_n414), .ZN(new_n429));
  AOI211_X1 g0229(.A(KEYINPUT75), .B(new_n413), .C1(new_n410), .C2(G20), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(KEYINPUT76), .B1(new_n421), .B2(new_n422), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT76), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n433), .B1(new_n419), .B2(new_n420), .ZN(new_n434));
  OAI21_X1  g0234(.A(G68), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(KEYINPUT16), .B1(new_n431), .B2(new_n435), .ZN(new_n436));
  OAI211_X1 g0236(.A(new_n404), .B(new_n408), .C1(new_n428), .C2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT17), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n408), .ZN(new_n440));
  INV_X1    g0240(.A(new_n255), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n202), .B1(new_n421), .B2(new_n422), .ZN(new_n442));
  NOR3_X1   g0242(.A1(new_n429), .A2(new_n430), .A3(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n441), .B1(new_n443), .B2(KEYINPUT16), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n431), .A2(new_n435), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT16), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n440), .B1(new_n444), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n448), .A2(KEYINPUT17), .A3(new_n404), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n408), .B1(new_n428), .B2(new_n436), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n403), .A2(G179), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n451), .B1(new_n317), .B2(new_n403), .ZN(new_n452));
  AND3_X1   g0252(.A1(new_n450), .A2(KEYINPUT18), .A3(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(KEYINPUT18), .B1(new_n450), .B2(new_n452), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n439), .B(new_n449), .C1(new_n453), .C2(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n455), .B1(new_n347), .B2(new_n348), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n392), .A2(new_n456), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n260), .A2(G97), .ZN(new_n458));
  OAI21_X1  g0258(.A(G107), .B1(new_n432), .B2(new_n434), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT6), .ZN(new_n460));
  INV_X1    g0260(.A(G97), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n461), .A2(new_n326), .ZN(new_n462));
  NOR2_X1   g0262(.A1(G97), .A2(G107), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n460), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n326), .A2(KEYINPUT6), .A3(G97), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(G20), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n264), .A2(G77), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n459), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n458), .B1(new_n469), .B2(new_n255), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n216), .A2(G33), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n252), .A2(new_n260), .A3(new_n254), .A4(new_n471), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n472), .A2(new_n461), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n470), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g0275(.A1(KEYINPUT79), .A2(G41), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(KEYINPUT5), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT5), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n478), .B1(KEYINPUT79), .B2(G41), .ZN(new_n479));
  INV_X1    g0279(.A(G45), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n480), .A2(G1), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n477), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  AND3_X1   g0282(.A1(new_n482), .A2(G257), .A3(new_n299), .ZN(new_n483));
  OAI211_X1 g0283(.A(G244), .B(new_n285), .C1(new_n278), .C2(new_n279), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT4), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(KEYINPUT78), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n276), .A2(G244), .A3(new_n285), .A4(new_n486), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n276), .A2(G250), .A3(G1698), .ZN(new_n490));
  NAND2_X1  g0290(.A1(G33), .A2(G283), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n488), .A2(new_n489), .A3(new_n490), .A4(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n483), .B1(new_n492), .B2(new_n291), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n482), .A2(new_n296), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(KEYINPUT80), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT80), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n493), .A2(new_n498), .A3(new_n495), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n497), .A2(new_n317), .A3(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n496), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(new_n332), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n475), .A2(new_n500), .A3(new_n502), .ZN(new_n503));
  AOI211_X1 g0303(.A(new_n458), .B(new_n473), .C1(new_n469), .C2(new_n255), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n492), .A2(new_n291), .ZN(new_n505));
  INV_X1    g0305(.A(new_n483), .ZN(new_n506));
  AND4_X1   g0306(.A1(new_n498), .A2(new_n505), .A3(new_n495), .A4(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n498), .B1(new_n493), .B2(new_n495), .ZN(new_n508));
  OAI21_X1  g0308(.A(G190), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n496), .A2(G200), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n504), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT24), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT86), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n217), .B(G87), .C1(new_n278), .C2(new_n279), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(KEYINPUT22), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT22), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n276), .A2(new_n516), .A3(new_n217), .A4(G87), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n377), .A2(G116), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n326), .A2(G20), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT23), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(KEYINPUT23), .B1(new_n326), .B2(G20), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  AND4_X1   g0325(.A1(new_n513), .A2(new_n518), .A3(new_n519), .A4(new_n525), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n524), .B1(new_n515), .B2(new_n517), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n513), .B1(new_n527), .B2(new_n519), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n512), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n518), .A2(new_n519), .A3(new_n525), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(KEYINPUT86), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n527), .A2(new_n513), .A3(new_n519), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n531), .A2(KEYINPUT24), .A3(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n529), .A2(new_n533), .A3(new_n255), .ZN(new_n534));
  NOR3_X1   g0334(.A1(new_n520), .A2(G1), .A3(new_n258), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT25), .ZN(new_n536));
  OR2_X1    g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AND4_X1   g0337(.A1(new_n260), .A2(new_n252), .A3(new_n254), .A4(new_n471), .ZN(new_n538));
  AOI22_X1  g0338(.A1(new_n538), .A2(G107), .B1(new_n536), .B2(new_n535), .ZN(new_n539));
  AND3_X1   g0339(.A1(new_n482), .A2(G264), .A3(new_n299), .ZN(new_n540));
  OAI211_X1 g0340(.A(G250), .B(new_n285), .C1(new_n278), .C2(new_n279), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT88), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n276), .A2(KEYINPUT88), .A3(G250), .A4(new_n285), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n276), .A2(G257), .A3(G1698), .ZN(new_n545));
  NAND2_X1  g0345(.A1(G33), .A2(G294), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n543), .A2(new_n544), .A3(new_n545), .A4(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n540), .B1(new_n547), .B2(new_n291), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n548), .A2(new_n398), .A3(new_n495), .ZN(new_n549));
  AOI211_X1 g0349(.A(new_n494), .B(new_n540), .C1(new_n547), .C2(new_n291), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n549), .B1(new_n550), .B2(G200), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n534), .A2(new_n537), .A3(new_n539), .A4(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n503), .A2(new_n511), .A3(new_n552), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n491), .B(new_n217), .C1(G33), .C2(new_n461), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n251), .B(new_n554), .C1(new_n217), .C2(G116), .ZN(new_n555));
  XOR2_X1   g0355(.A(new_n555), .B(KEYINPUT20), .Z(new_n556));
  NOR2_X1   g0356(.A1(new_n260), .A2(G116), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  OAI21_X1  g0358(.A(KEYINPUT85), .B1(new_n472), .B2(new_n223), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  NOR3_X1   g0360(.A1(new_n472), .A2(KEYINPUT85), .A3(new_n223), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n556), .B(new_n558), .C1(new_n560), .C2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT84), .ZN(new_n563));
  OR2_X1    g0363(.A1(KEYINPUT83), .A2(G303), .ZN(new_n564));
  NAND2_X1  g0364(.A1(KEYINPUT83), .A2(G303), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n566), .A2(new_n276), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n285), .A2(G257), .ZN(new_n568));
  NAND2_X1  g0368(.A1(G264), .A2(G1698), .ZN(new_n569));
  AOI22_X1  g0369(.A1(new_n417), .A2(new_n418), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n563), .B1(new_n567), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n568), .A2(new_n569), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n276), .A2(new_n572), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n573), .B(KEYINPUT84), .C1(new_n276), .C2(new_n566), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n571), .A2(new_n574), .A3(new_n291), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n482), .A2(G270), .A3(new_n299), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n575), .A2(new_n495), .A3(new_n576), .ZN(new_n577));
  AND2_X1   g0377(.A1(new_n577), .A2(G169), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n562), .A2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT21), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n562), .A2(new_n578), .A3(KEYINPUT21), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n577), .A2(new_n332), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n562), .A2(new_n583), .ZN(new_n584));
  XNOR2_X1  g0384(.A(new_n555), .B(KEYINPUT20), .ZN(new_n585));
  INV_X1    g0385(.A(new_n561), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n585), .B1(new_n586), .B2(new_n559), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n577), .A2(G200), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n575), .A2(G190), .A3(new_n495), .A4(new_n576), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n587), .A2(new_n588), .A3(new_n558), .A4(new_n589), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n581), .A2(new_n582), .A3(new_n584), .A4(new_n590), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n553), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n534), .A2(new_n537), .A3(new_n539), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(KEYINPUT87), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT87), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n534), .A2(new_n595), .A3(new_n537), .A4(new_n539), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n550), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(G169), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n550), .A2(G179), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n597), .A2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(G87), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n603), .A2(new_n461), .A3(new_n326), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n352), .A2(new_n217), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n604), .A2(new_n605), .A3(KEYINPUT19), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n217), .B(G68), .C1(new_n278), .C2(new_n279), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n266), .A2(new_n461), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n606), .B(new_n607), .C1(KEYINPUT19), .C2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n255), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n261), .A2(new_n337), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n612), .B1(G87), .B2(new_n538), .ZN(new_n613));
  INV_X1    g0413(.A(new_n311), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n216), .A2(G45), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n299), .A2(G250), .A3(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n229), .A2(new_n285), .ZN(new_n618));
  OAI221_X1 g0418(.A(new_n618), .B1(G244), .B2(new_n285), .C1(new_n278), .C2(new_n279), .ZN(new_n619));
  NAND2_X1  g0419(.A1(G33), .A2(G116), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n617), .B1(new_n621), .B2(new_n291), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n615), .A2(new_n296), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n614), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n613), .A2(KEYINPUT82), .A3(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT82), .ZN(new_n628));
  AOI22_X1  g0428(.A1(new_n255), .A2(new_n609), .B1(new_n261), .B2(new_n337), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n629), .B1(new_n603), .B2(new_n472), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n628), .B1(new_n630), .B2(new_n625), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n290), .B1(new_n620), .B2(new_n619), .ZN(new_n632));
  NOR4_X1   g0432(.A1(new_n632), .A2(new_n398), .A3(new_n623), .A4(new_n617), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n627), .A2(new_n631), .A3(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(G169), .B1(new_n622), .B2(new_n624), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n472), .A2(new_n337), .ZN(new_n637));
  OAI21_X1  g0437(.A(KEYINPUT81), .B1(new_n612), .B2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT81), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n629), .B(new_n639), .C1(new_n337), .C2(new_n472), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n636), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n622), .A2(new_n624), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n332), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n635), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n592), .A2(new_n602), .A3(new_n647), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n457), .A2(new_n648), .ZN(G372));
  INV_X1    g0449(.A(new_n323), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT18), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n403), .A2(new_n317), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n652), .B1(G179), .B2(new_n403), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n651), .B1(new_n448), .B2(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n450), .A2(KEYINPUT18), .A3(new_n452), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AOI22_X1  g0456(.A1(new_n367), .A2(new_n362), .B1(new_n372), .B2(new_n373), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n657), .A2(new_n385), .ZN(new_n658));
  INV_X1    g0458(.A(new_n343), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n658), .B1(new_n659), .B2(new_n390), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n449), .A2(new_n439), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n656), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n650), .B1(new_n662), .B2(new_n316), .ZN(new_n663));
  INV_X1    g0463(.A(new_n503), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT26), .ZN(new_n665));
  NOR3_X1   g0465(.A1(new_n630), .A2(new_n625), .A3(new_n633), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n666), .B1(new_n641), .B2(new_n644), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n664), .A2(new_n665), .A3(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(KEYINPUT26), .B1(new_n646), .B2(new_n503), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n668), .A2(new_n669), .A3(new_n645), .ZN(new_n670));
  AND4_X1   g0470(.A1(new_n503), .A2(new_n511), .A3(new_n667), .A4(new_n552), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n593), .A2(new_n601), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n672), .A2(new_n581), .A3(new_n582), .A4(new_n584), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT89), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n671), .A2(new_n673), .A3(KEYINPUT89), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n670), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n663), .B1(new_n457), .B2(new_n678), .ZN(G369));
  OR2_X1    g0479(.A1(new_n591), .A2(KEYINPUT90), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n258), .A2(G20), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n216), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n682), .A2(KEYINPUT27), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(KEYINPUT27), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n683), .A2(G213), .A3(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(G343), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n562), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n591), .A2(KEYINPUT90), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n680), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n581), .A2(new_n582), .A3(new_n584), .ZN(new_n691));
  OR2_X1    g0491(.A1(new_n691), .A2(new_n688), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n690), .A2(G330), .A3(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n687), .ZN(new_n695));
  INV_X1    g0495(.A(new_n601), .ZN(new_n696));
  AOI22_X1  g0496(.A1(new_n594), .A2(new_n596), .B1(new_n696), .B2(new_n695), .ZN(new_n697));
  INV_X1    g0497(.A(new_n552), .ZN(new_n698));
  OAI22_X1  g0498(.A1(new_n602), .A2(new_n695), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n694), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n691), .A2(new_n695), .ZN(new_n701));
  NOR3_X1   g0501(.A1(new_n697), .A2(new_n701), .A3(new_n698), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n672), .A2(new_n687), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n700), .A2(new_n704), .ZN(G399));
  INV_X1    g0505(.A(new_n218), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(G41), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n604), .A2(G116), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n708), .A2(G1), .A3(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n710), .B1(new_n209), .B2(new_n708), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n711), .B(KEYINPUT28), .ZN(new_n712));
  NOR3_X1   g0512(.A1(new_n678), .A2(KEYINPUT29), .A3(new_n687), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT29), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n665), .B1(new_n646), .B2(new_n503), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT92), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n664), .A2(KEYINPUT26), .A3(new_n667), .ZN(new_n718));
  OAI211_X1 g0518(.A(KEYINPUT92), .B(new_n665), .C1(new_n646), .C2(new_n503), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n717), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n696), .B1(new_n594), .B2(new_n596), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n671), .B1(new_n721), .B2(new_n691), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n720), .A2(new_n645), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n714), .B1(new_n723), .B2(new_n695), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n713), .A2(new_n724), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n592), .A2(new_n602), .A3(new_n647), .A4(new_n695), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT30), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT91), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n583), .A2(new_n728), .ZN(new_n729));
  NOR3_X1   g0529(.A1(new_n577), .A2(KEYINPUT91), .A3(new_n332), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n548), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n642), .B1(new_n497), .B2(new_n499), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n727), .B1(new_n731), .B2(new_n733), .ZN(new_n734));
  XNOR2_X1  g0534(.A(new_n583), .B(new_n728), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n735), .A2(KEYINPUT30), .A3(new_n548), .A4(new_n732), .ZN(new_n736));
  NOR3_X1   g0536(.A1(new_n501), .A2(G179), .A3(new_n643), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n737), .A2(new_n598), .A3(new_n577), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n734), .A2(new_n736), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(new_n687), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n726), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(KEYINPUT31), .ZN(new_n742));
  AOI21_X1  g0542(.A(KEYINPUT31), .B1(new_n739), .B2(new_n687), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(G330), .ZN(new_n746));
  AND2_X1   g0546(.A1(new_n725), .A2(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n712), .B1(new_n747), .B2(G1), .ZN(new_n748));
  XOR2_X1   g0548(.A(new_n748), .B(KEYINPUT93), .Z(G364));
  XNOR2_X1  g0549(.A(new_n693), .B(KEYINPUT94), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n681), .A2(G45), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n708), .A2(G1), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n690), .A2(new_n692), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  OAI211_X1 g0554(.A(new_n750), .B(new_n752), .C1(G330), .C2(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n214), .B1(new_n217), .B2(G169), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n217), .A2(new_n332), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT96), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(G190), .A2(G200), .ZN(new_n760));
  OAI21_X1  g0560(.A(KEYINPUT96), .B1(new_n217), .B2(new_n332), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n759), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(KEYINPUT97), .ZN(new_n763));
  OR2_X1    g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n762), .A2(new_n763), .ZN(new_n765));
  AND2_X1   g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n398), .A2(G200), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n759), .A2(new_n768), .A3(new_n761), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  AOI22_X1  g0570(.A1(new_n767), .A2(G77), .B1(G58), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n757), .A2(G200), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(new_n398), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n771), .B1(new_n227), .B2(new_n774), .ZN(new_n775));
  XOR2_X1   g0575(.A(new_n775), .B(KEYINPUT98), .Z(new_n776));
  NAND2_X1  g0576(.A1(new_n768), .A2(new_n332), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G20), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n772), .A2(G190), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  OAI221_X1 g0581(.A(new_n276), .B1(new_n779), .B2(new_n461), .C1(new_n781), .C2(new_n202), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n217), .A2(G179), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n311), .A2(G190), .A3(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n782), .B1(G87), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n783), .A2(new_n760), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(new_n412), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n788), .B(KEYINPUT32), .ZN(new_n789));
  AND3_X1   g0589(.A1(new_n311), .A2(new_n398), .A3(new_n783), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(new_n326), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NAND4_X1  g0593(.A1(new_n776), .A2(new_n786), .A3(new_n789), .A4(new_n793), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n773), .A2(G326), .B1(new_n778), .B2(G294), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT99), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n790), .A2(G283), .ZN(new_n797));
  INV_X1    g0597(.A(new_n787), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n276), .B1(new_n798), .B2(G329), .ZN(new_n799));
  INV_X1    g0599(.A(G303), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n799), .B1(new_n800), .B2(new_n784), .ZN(new_n801));
  XNOR2_X1  g0601(.A(KEYINPUT33), .B(G317), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n801), .B1(new_n780), .B2(new_n802), .ZN(new_n803));
  AND3_X1   g0603(.A1(new_n796), .A2(new_n797), .A3(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(G311), .ZN(new_n805));
  INV_X1    g0605(.A(G322), .ZN(new_n806));
  OAI221_X1 g0606(.A(new_n804), .B1(new_n805), .B2(new_n766), .C1(new_n806), .C2(new_n769), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n756), .B1(new_n794), .B2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n756), .ZN(new_n809));
  NOR2_X1   g0609(.A1(G13), .A2(G33), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n811), .A2(G20), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n809), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n209), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(new_n480), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n706), .A2(new_n276), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n815), .B(new_n816), .C1(new_n480), .C2(new_n245), .ZN(new_n817));
  INV_X1    g0617(.A(G355), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n276), .A2(new_n218), .ZN(new_n819));
  XOR2_X1   g0619(.A(new_n819), .B(KEYINPUT95), .Z(new_n820));
  OAI221_X1 g0620(.A(new_n817), .B1(G116), .B2(new_n218), .C1(new_n818), .C2(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n808), .B1(new_n813), .B2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n812), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n822), .B1(new_n754), .B2(new_n823), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n755), .B1(new_n752), .B2(new_n824), .ZN(G396));
  INV_X1    g0625(.A(new_n752), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n809), .A2(new_n810), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n770), .A2(G143), .B1(G150), .B2(new_n780), .ZN(new_n829));
  INV_X1    g0629(.A(G137), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n829), .B1(new_n830), .B2(new_n774), .C1(new_n766), .C2(new_n412), .ZN(new_n831));
  XOR2_X1   g0631(.A(new_n831), .B(KEYINPUT101), .Z(new_n832));
  OR2_X1    g0632(.A1(new_n832), .A2(KEYINPUT34), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(KEYINPUT34), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n790), .A2(G68), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n835), .B1(new_n227), .B2(new_n784), .ZN(new_n836));
  XNOR2_X1  g0636(.A(new_n836), .B(KEYINPUT102), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n283), .B(new_n837), .C1(G58), .C2(new_n778), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n798), .A2(G132), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n833), .A2(new_n834), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n283), .B1(new_n787), .B2(new_n805), .ZN(new_n841));
  XNOR2_X1  g0641(.A(KEYINPUT100), .B(G283), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  OAI22_X1  g0643(.A1(new_n781), .A2(new_n843), .B1(new_n774), .B2(new_n800), .ZN(new_n844));
  AOI211_X1 g0644(.A(new_n841), .B(new_n844), .C1(G97), .C2(new_n778), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n790), .A2(G87), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n767), .A2(G116), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n770), .A2(G294), .B1(new_n785), .B2(G107), .ZN(new_n848));
  NAND4_X1  g0648(.A1(new_n845), .A2(new_n846), .A3(new_n847), .A4(new_n848), .ZN(new_n849));
  AND2_X1   g0649(.A1(new_n840), .A2(new_n849), .ZN(new_n850));
  OAI221_X1 g0650(.A(new_n826), .B1(G77), .B2(new_n828), .C1(new_n850), .C2(new_n756), .ZN(new_n851));
  OR2_X1    g0651(.A1(new_n851), .A2(KEYINPUT103), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(KEYINPUT103), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n343), .A2(new_n687), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n344), .A2(new_n345), .B1(new_n342), .B2(new_n687), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n855), .B1(new_n856), .B2(new_n659), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n852), .B(new_n853), .C1(new_n811), .C2(new_n858), .ZN(new_n859));
  XOR2_X1   g0659(.A(new_n859), .B(KEYINPUT104), .Z(new_n860));
  OAI21_X1  g0660(.A(new_n857), .B1(new_n678), .B2(new_n687), .ZN(new_n861));
  AND3_X1   g0661(.A1(new_n668), .A2(new_n669), .A3(new_n645), .ZN(new_n862));
  AND3_X1   g0662(.A1(new_n671), .A2(new_n673), .A3(KEYINPUT89), .ZN(new_n863));
  AOI21_X1  g0663(.A(KEYINPUT89), .B1(new_n671), .B2(new_n673), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n862), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n865), .A2(new_n695), .A3(new_n858), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n861), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n746), .A2(new_n867), .ZN(new_n868));
  OR2_X1    g0668(.A1(new_n868), .A2(KEYINPUT105), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(KEYINPUT105), .ZN(new_n870));
  OR2_X1    g0670(.A1(new_n746), .A2(new_n867), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n869), .A2(new_n752), .A3(new_n870), .A4(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n860), .A2(new_n872), .ZN(G384));
  INV_X1    g0673(.A(KEYINPUT40), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n416), .A2(new_n426), .A3(new_n424), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n446), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n440), .B1(new_n444), .B2(new_n876), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n877), .A2(new_n685), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n437), .B1(new_n877), .B2(new_n653), .ZN(new_n879));
  OAI21_X1  g0679(.A(KEYINPUT37), .B1(new_n879), .B2(new_n878), .ZN(new_n880));
  INV_X1    g0680(.A(new_n685), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n450), .B1(new_n452), .B2(new_n881), .ZN(new_n882));
  XOR2_X1   g0682(.A(KEYINPUT107), .B(KEYINPUT37), .Z(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n882), .A2(new_n437), .A3(new_n884), .ZN(new_n885));
  AOI22_X1  g0685(.A1(new_n455), .A2(new_n878), .B1(new_n880), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(KEYINPUT108), .B1(new_n886), .B2(KEYINPUT38), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(KEYINPUT38), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT108), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT38), .ZN(new_n890));
  AOI21_X1  g0690(.A(KEYINPUT16), .B1(new_n431), .B2(new_n424), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n408), .B1(new_n428), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n881), .ZN(new_n893));
  AND2_X1   g0693(.A1(new_n449), .A2(new_n439), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n893), .B1(new_n894), .B2(new_n656), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n882), .A2(new_n437), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n892), .A2(new_n452), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n893), .A2(new_n897), .A3(new_n437), .ZN(new_n898));
  AOI22_X1  g0698(.A1(new_n896), .A2(new_n884), .B1(new_n898), .B2(KEYINPUT37), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n889), .B(new_n890), .C1(new_n895), .C2(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n887), .A2(new_n888), .A3(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT106), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n902), .B1(new_n387), .B2(new_n695), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n658), .A2(KEYINPUT106), .A3(new_n687), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n387), .B(new_n390), .C1(new_n385), .C2(new_n695), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n857), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT31), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n908), .B1(new_n726), .B2(new_n740), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n901), .B(new_n907), .C1(new_n909), .C2(new_n743), .ZN(new_n910));
  AOI21_X1  g0710(.A(KEYINPUT106), .B1(new_n658), .B2(new_n687), .ZN(new_n911));
  NOR4_X1   g0711(.A1(new_n657), .A2(new_n385), .A3(new_n902), .A4(new_n695), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n906), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n858), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n914), .B1(new_n742), .B2(new_n744), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT109), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n884), .B1(new_n882), .B2(new_n916), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n896), .B(new_n917), .ZN(new_n918));
  AND3_X1   g0718(.A1(new_n455), .A2(new_n450), .A3(new_n881), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n890), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n874), .B1(new_n920), .B2(new_n888), .ZN(new_n921));
  AOI22_X1  g0721(.A1(new_n874), .A2(new_n910), .B1(new_n915), .B2(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n457), .B1(new_n742), .B2(new_n744), .ZN(new_n923));
  XOR2_X1   g0723(.A(new_n922), .B(new_n923), .Z(new_n924));
  AND2_X1   g0724(.A1(new_n924), .A2(G330), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n654), .A2(new_n655), .A3(new_n685), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n866), .A2(new_n855), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n927), .A2(new_n901), .A3(new_n913), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n901), .A2(KEYINPUT39), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT39), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n920), .A2(new_n930), .A3(new_n888), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(KEYINPUT110), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT110), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n929), .A2(new_n934), .A3(new_n931), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n387), .A2(new_n687), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n926), .B(new_n928), .C1(new_n936), .C2(new_n938), .ZN(new_n939));
  OAI211_X1 g0739(.A(new_n392), .B(new_n456), .C1(new_n713), .C2(new_n724), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(new_n663), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n939), .B(new_n941), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n925), .B(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n943), .B1(new_n216), .B2(new_n681), .ZN(new_n944));
  OAI211_X1 g0744(.A(G20), .B(new_n214), .C1(new_n466), .C2(KEYINPUT35), .ZN(new_n945));
  AOI211_X1 g0745(.A(new_n223), .B(new_n945), .C1(KEYINPUT35), .C2(new_n466), .ZN(new_n946));
  XOR2_X1   g0746(.A(new_n946), .B(KEYINPUT36), .Z(new_n947));
  NAND3_X1  g0747(.A1(new_n814), .A2(G77), .A3(new_n409), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(G50), .B2(new_n202), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n949), .A2(G1), .A3(new_n258), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n944), .A2(new_n947), .A3(new_n950), .ZN(G367));
  INV_X1    g0751(.A(new_n511), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n664), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n475), .A2(new_n687), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n702), .A2(new_n956), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n957), .A2(KEYINPUT42), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n503), .B1(new_n602), .B2(new_n952), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(new_n695), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n957), .A2(KEYINPUT42), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n958), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n630), .A2(new_n687), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n667), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(new_n645), .B2(new_n963), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(KEYINPUT43), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n962), .A2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(new_n700), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n955), .B1(new_n503), .B2(new_n695), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n967), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n969), .ZN(new_n971));
  OAI211_X1 g0771(.A(new_n962), .B(new_n966), .C1(new_n700), .C2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n965), .A2(KEYINPUT43), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n973), .B(new_n974), .ZN(new_n975));
  XNOR2_X1  g0775(.A(KEYINPUT111), .B(KEYINPUT41), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n707), .B(new_n976), .Z(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT112), .ZN(new_n979));
  INV_X1    g0779(.A(new_n702), .ZN(new_n980));
  INV_X1    g0780(.A(new_n701), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n980), .B1(new_n699), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n750), .A2(new_n982), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n982), .A2(new_n693), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n725), .A2(new_n746), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n979), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n984), .B1(new_n750), .B2(new_n982), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n747), .A2(KEYINPUT112), .A3(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n704), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT45), .ZN(new_n992));
  NOR3_X1   g0792(.A1(new_n991), .A2(new_n971), .A3(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(KEYINPUT45), .B1(new_n704), .B2(new_n969), .ZN(new_n994));
  OR2_X1    g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  OR3_X1    g0795(.A1(new_n704), .A2(KEYINPUT44), .A3(new_n969), .ZN(new_n996));
  OAI21_X1  g0796(.A(KEYINPUT44), .B1(new_n704), .B2(new_n969), .ZN(new_n997));
  AND2_X1   g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n995), .A2(new_n700), .A3(new_n998), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n997), .B(new_n996), .C1(new_n993), .C2(new_n994), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(new_n968), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n988), .A2(new_n990), .A3(new_n999), .A4(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n978), .B1(new_n1002), .B2(new_n747), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n751), .A2(G1), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n1004), .B(KEYINPUT113), .Z(new_n1005));
  OAI21_X1  g0805(.A(new_n975), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n791), .A2(new_n461), .B1(new_n566), .B2(new_n769), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n773), .A2(G311), .B1(new_n778), .B2(G107), .ZN(new_n1008));
  INV_X1    g0808(.A(G294), .ZN(new_n1009));
  OAI211_X1 g0809(.A(new_n1008), .B(new_n283), .C1(new_n1009), .C2(new_n781), .ZN(new_n1010));
  OAI21_X1  g0810(.A(KEYINPUT46), .B1(new_n784), .B2(new_n223), .ZN(new_n1011));
  OR3_X1    g0811(.A1(new_n784), .A2(KEYINPUT46), .A3(new_n223), .ZN(new_n1012));
  AOI211_X1 g0812(.A(new_n1007), .B(new_n1010), .C1(new_n1011), .C2(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(G317), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n1013), .B1(new_n1014), .B2(new_n787), .C1(new_n766), .C2(new_n843), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT114), .ZN(new_n1016));
  INV_X1    g0816(.A(G150), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n769), .A2(new_n1017), .B1(new_n784), .B2(new_n201), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n283), .B1(new_n773), .B2(G143), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n778), .A2(G68), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n1019), .B(new_n1020), .C1(new_n412), .C2(new_n781), .ZN(new_n1021));
  AOI211_X1 g0821(.A(new_n1018), .B(new_n1021), .C1(G137), .C2(new_n798), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n1022), .B1(new_n227), .B2(new_n766), .C1(new_n339), .C2(new_n791), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1016), .A2(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT47), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n752), .B1(new_n1025), .B2(new_n809), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n816), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n813), .B1(new_n218), .B2(new_n337), .C1(new_n241), .C2(new_n1027), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n1026), .B(new_n1028), .C1(new_n823), .C2(new_n965), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1006), .A2(new_n1029), .ZN(G387));
  NAND2_X1  g0830(.A1(new_n747), .A2(new_n989), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n986), .A2(new_n987), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1031), .A2(new_n1032), .A3(new_n707), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n989), .A2(new_n1005), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT115), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n238), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1035), .B1(new_n1036), .B2(new_n480), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n269), .A2(new_n227), .ZN(new_n1038));
  AOI211_X1 g0838(.A(G116), .B(new_n604), .C1(new_n1038), .C2(KEYINPUT50), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(G68), .A2(G77), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n1038), .A2(KEYINPUT50), .ZN(new_n1041));
  NAND4_X1  g0841(.A1(new_n1039), .A2(new_n480), .A3(new_n1040), .A4(new_n1041), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n238), .A2(KEYINPUT115), .A3(G45), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1037), .A2(new_n816), .A3(new_n1042), .A4(new_n1043), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1044), .B1(G107), .B2(new_n218), .C1(new_n709), .C2(new_n820), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n752), .B1(new_n1045), .B2(new_n813), .ZN(new_n1046));
  XOR2_X1   g0846(.A(new_n1046), .B(KEYINPUT116), .Z(new_n1047));
  AOI22_X1  g0847(.A1(new_n770), .A2(G317), .B1(G311), .B2(new_n780), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n1048), .B1(new_n806), .B2(new_n774), .C1(new_n766), .C2(new_n566), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT48), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1050), .B1(new_n1009), .B2(new_n784), .C1(new_n779), .C2(new_n843), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT49), .ZN(new_n1052));
  OR2_X1    g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n798), .A2(G326), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n283), .B(new_n1054), .C1(new_n791), .C2(new_n223), .ZN(new_n1055));
  OR2_X1    g0855(.A1(new_n1055), .A2(KEYINPUT118), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1055), .A2(KEYINPUT118), .ZN(new_n1058));
  NAND4_X1  g0858(.A1(new_n1053), .A2(new_n1056), .A3(new_n1057), .A4(new_n1058), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n766), .A2(new_n202), .B1(new_n270), .B2(new_n781), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT117), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n276), .B1(new_n787), .B2(new_n1017), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n774), .A2(new_n412), .B1(new_n779), .B2(new_n337), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n1062), .B(new_n1063), .C1(G77), .C2(new_n785), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n770), .A2(G50), .B1(G97), .B2(new_n790), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1061), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  AND2_X1   g0866(.A1(new_n1059), .A2(new_n1066), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n1047), .B1(new_n699), .B2(new_n823), .C1(new_n1067), .C2(new_n756), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1033), .A2(new_n1034), .A3(new_n1068), .ZN(G393));
  INV_X1    g0869(.A(new_n1001), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n1000), .A2(new_n968), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1031), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1002), .A2(new_n707), .A3(new_n1072), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n813), .B1(new_n461), .B2(new_n218), .C1(new_n248), .C2(new_n1027), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n767), .A2(new_n269), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n774), .A2(new_n1017), .B1(new_n412), .B2(new_n769), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT51), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n785), .A2(G68), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n780), .A2(G50), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n283), .B1(new_n798), .B2(G143), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n778), .A2(G77), .ZN(new_n1081));
  AND4_X1   g0881(.A1(new_n846), .A2(new_n1079), .A3(new_n1080), .A4(new_n1081), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n1075), .A2(new_n1077), .A3(new_n1078), .A4(new_n1082), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n781), .A2(new_n566), .B1(new_n779), .B2(new_n223), .ZN(new_n1084));
  XOR2_X1   g0884(.A(new_n1084), .B(KEYINPUT120), .Z(new_n1085));
  OAI21_X1  g0885(.A(new_n283), .B1(new_n787), .B2(new_n806), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n1086), .B(new_n792), .C1(new_n785), .C2(new_n842), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1085), .B(new_n1087), .C1(new_n1009), .C2(new_n766), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n770), .A2(G311), .B1(G317), .B2(new_n773), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT52), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1083), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n752), .B1(new_n1091), .B2(new_n809), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n1074), .B(new_n1092), .C1(new_n969), .C2(new_n823), .ZN(new_n1093));
  INV_X1    g0893(.A(KEYINPUT119), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n999), .A2(new_n1001), .A3(KEYINPUT119), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1095), .A2(new_n1005), .A3(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1073), .A2(new_n1093), .A3(new_n1097), .ZN(G390));
  OAI211_X1 g0898(.A(G330), .B(new_n858), .C1(new_n909), .C2(new_n743), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n913), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n937), .B1(new_n927), .B2(new_n913), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(new_n933), .B2(new_n935), .ZN(new_n1103));
  AND2_X1   g0903(.A1(new_n920), .A2(new_n888), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n723), .A2(new_n695), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n856), .A2(new_n659), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n855), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  AOI211_X1 g0907(.A(new_n937), .B(new_n1104), .C1(new_n1107), .C2(new_n913), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1101), .B1(new_n1103), .B2(new_n1108), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n1104), .A2(new_n937), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1107), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1110), .B1(new_n1111), .B2(new_n1100), .ZN(new_n1112));
  OR2_X1    g0912(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1113));
  AND3_X1   g0913(.A1(new_n929), .A2(new_n934), .A3(new_n931), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n934), .B1(new_n929), .B2(new_n931), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n1112), .B(new_n1113), .C1(new_n1116), .C2(new_n1102), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1109), .A2(new_n1117), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n745), .A2(new_n392), .A3(new_n456), .A4(G330), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n940), .A2(new_n1119), .A3(new_n663), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n927), .B1(new_n1122), .B2(new_n1101), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1113), .A2(new_n1111), .A3(new_n1121), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1120), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1118), .A2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1109), .A2(new_n1117), .A3(new_n1125), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1127), .A2(new_n707), .A3(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1109), .A2(new_n1117), .A3(new_n1005), .ZN(new_n1130));
  INV_X1    g0930(.A(G132), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n791), .A2(new_n227), .B1(new_n1131), .B2(new_n769), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n283), .B1(new_n778), .B2(G159), .ZN(new_n1133));
  INV_X1    g0933(.A(G128), .ZN(new_n1134));
  OAI221_X1 g0934(.A(new_n1133), .B1(new_n781), .B2(new_n830), .C1(new_n1134), .C2(new_n774), .ZN(new_n1135));
  XOR2_X1   g0935(.A(KEYINPUT54), .B(G143), .Z(new_n1136));
  AOI211_X1 g0936(.A(new_n1132), .B(new_n1135), .C1(new_n767), .C2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n798), .A2(G125), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n784), .A2(new_n1017), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n1139), .B(KEYINPUT53), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1137), .A2(new_n1138), .A3(new_n1140), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(new_n1141), .B(KEYINPUT121), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n835), .B1(new_n603), .B2(new_n784), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n780), .A2(G107), .B1(new_n773), .B2(G283), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n770), .A2(G116), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n276), .B1(new_n798), .B2(G294), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n1144), .A2(new_n1145), .A3(new_n1081), .A4(new_n1146), .ZN(new_n1147));
  AOI211_X1 g0947(.A(new_n1143), .B(new_n1147), .C1(new_n767), .C2(G97), .ZN(new_n1148));
  XOR2_X1   g0948(.A(new_n1148), .B(KEYINPUT122), .Z(new_n1149));
  NAND2_X1  g0949(.A1(new_n1142), .A2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n752), .B1(new_n1150), .B2(new_n809), .ZN(new_n1151));
  OAI221_X1 g0951(.A(new_n1151), .B1(new_n269), .B2(new_n828), .C1(new_n1116), .C2(new_n811), .ZN(new_n1152));
  AND2_X1   g0952(.A1(new_n1130), .A2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(KEYINPUT123), .B1(new_n1129), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1129), .A2(KEYINPUT123), .A3(new_n1153), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1155), .A2(new_n1156), .ZN(G378));
  INV_X1    g0957(.A(new_n1120), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1128), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n928), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1160), .B1(new_n1116), .B2(new_n937), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT125), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n274), .A2(new_n685), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT55), .ZN(new_n1164));
  AND3_X1   g0964(.A1(new_n316), .A2(new_n1164), .A3(new_n323), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1164), .B1(new_n316), .B2(new_n323), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1163), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n316), .A2(new_n323), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1168), .A2(KEYINPUT55), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n316), .A2(new_n1164), .A3(new_n323), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1163), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1169), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(KEYINPUT124), .B(KEYINPUT56), .ZN(new_n1173));
  AND3_X1   g0973(.A1(new_n1167), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1173), .B1(new_n1167), .B2(new_n1172), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1162), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n922), .A2(G330), .A3(new_n1176), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n907), .B1(new_n909), .B2(new_n743), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n901), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n874), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n745), .A2(new_n921), .A3(new_n907), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1180), .A2(G330), .A3(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1167), .A2(new_n1172), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1173), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1167), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1186));
  AOI21_X1  g0986(.A(KEYINPUT125), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1182), .A2(new_n1187), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1161), .A2(new_n926), .A3(new_n1177), .A4(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1177), .A2(new_n1188), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1190), .A2(new_n939), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1189), .A2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1159), .A2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT57), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1159), .A2(new_n1192), .A3(KEYINPUT57), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1195), .A2(new_n707), .A3(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1192), .A2(new_n1005), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n810), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n780), .A2(G132), .B1(new_n773), .B2(G125), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1136), .ZN(new_n1201));
  OAI221_X1 g1001(.A(new_n1200), .B1(new_n1134), .B2(new_n769), .C1(new_n784), .C2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(G137), .B2(new_n767), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1203), .B1(new_n1017), .B2(new_n779), .ZN(new_n1204));
  XOR2_X1   g1004(.A(new_n1204), .B(KEYINPUT59), .Z(new_n1205));
  AOI21_X1  g1005(.A(G41), .B1(new_n790), .B2(G159), .ZN(new_n1206));
  AOI21_X1  g1006(.A(G33), .B1(new_n798), .B2(G124), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n227), .B1(new_n278), .B2(G41), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n769), .A2(new_n326), .B1(new_n784), .B2(new_n339), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n780), .A2(G97), .B1(new_n773), .B2(G116), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n790), .A2(G58), .ZN(new_n1212));
  AOI211_X1 g1012(.A(G41), .B(new_n276), .C1(new_n798), .C2(G283), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1211), .A2(new_n1020), .A3(new_n1212), .A4(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n337), .ZN(new_n1215));
  AOI211_X1 g1015(.A(new_n1210), .B(new_n1214), .C1(new_n767), .C2(new_n1215), .ZN(new_n1216));
  XOR2_X1   g1016(.A(new_n1216), .B(KEYINPUT58), .Z(new_n1217));
  NAND3_X1  g1017(.A1(new_n1208), .A2(new_n1209), .A3(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n752), .B1(new_n1218), .B2(new_n809), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1199), .B(new_n1219), .C1(G50), .C2(new_n828), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1198), .A2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1197), .A2(new_n1222), .ZN(G375));
  NAND2_X1  g1023(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(new_n1120), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1226), .A2(new_n977), .A3(new_n1126), .ZN(new_n1227));
  OAI22_X1  g1027(.A1(new_n781), .A2(new_n223), .B1(new_n774), .B2(new_n1009), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1228), .B1(new_n1215), .B2(new_n778), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n276), .B1(new_n798), .B2(G303), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n770), .A2(G283), .B1(G77), .B2(new_n790), .ZN(new_n1231));
  AND3_X1   g1031(.A1(new_n1229), .A2(new_n1230), .A3(new_n1231), .ZN(new_n1232));
  OAI221_X1 g1032(.A(new_n1232), .B1(new_n461), .B2(new_n784), .C1(new_n326), .C2(new_n766), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n774), .A2(new_n1131), .B1(new_n779), .B2(new_n227), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1212), .B1(new_n830), .B2(new_n769), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n276), .B1(new_n781), .B2(new_n1201), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n787), .A2(new_n1134), .ZN(new_n1237));
  NOR4_X1   g1037(.A1(new_n1234), .A2(new_n1235), .A3(new_n1236), .A4(new_n1237), .ZN(new_n1238));
  OAI221_X1 g1038(.A(new_n1238), .B1(new_n1017), .B2(new_n766), .C1(new_n412), .C2(new_n784), .ZN(new_n1239));
  AND2_X1   g1039(.A1(new_n1233), .A2(new_n1239), .ZN(new_n1240));
  OAI22_X1  g1040(.A1(new_n1240), .A2(new_n756), .B1(G68), .B2(new_n828), .ZN(new_n1241));
  AOI211_X1 g1041(.A(new_n752), .B(new_n1241), .C1(new_n1100), .C2(new_n810), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(new_n1224), .B2(new_n1005), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1227), .A2(new_n1243), .ZN(G381));
  NAND2_X1  g1044(.A1(new_n1129), .A2(new_n1153), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(G375), .A2(new_n1245), .ZN(new_n1246));
  OR3_X1    g1046(.A1(G390), .A2(G396), .A3(G393), .ZN(new_n1247));
  NOR4_X1   g1047(.A1(new_n1247), .A2(G387), .A3(G384), .A4(G381), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1246), .A2(new_n1248), .ZN(G407));
  OAI21_X1  g1049(.A(new_n1246), .B1(new_n1248), .B2(new_n686), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(G213), .ZN(G409));
  INV_X1    g1051(.A(G390), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(G387), .A2(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1006), .A2(new_n1029), .A3(G390), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  XNOR2_X1  g1055(.A(G393), .B(G396), .ZN(new_n1256));
  AOI21_X1  g1056(.A(G390), .B1(new_n1006), .B2(new_n1029), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT127), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1256), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1255), .A2(new_n1259), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1253), .A2(new_n1258), .A3(new_n1254), .A4(new_n1256), .ZN(new_n1261));
  AND2_X1   g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1225), .A2(KEYINPUT60), .A3(new_n1120), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1263), .A2(new_n707), .A3(new_n1126), .ZN(new_n1264));
  AOI21_X1  g1064(.A(KEYINPUT60), .B1(new_n1225), .B2(new_n1120), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1243), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1266), .A2(new_n860), .A3(new_n872), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1265), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1268), .A2(new_n707), .A3(new_n1126), .A4(new_n1263), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1269), .A2(G384), .A3(new_n1243), .ZN(new_n1270));
  INV_X1    g1070(.A(G213), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1271), .A2(G343), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(G2897), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1267), .A2(new_n1270), .A3(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1273), .B1(new_n1267), .B2(new_n1270), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  AND3_X1   g1077(.A1(new_n1159), .A2(KEYINPUT57), .A3(new_n1192), .ZN(new_n1278));
  AOI21_X1  g1078(.A(KEYINPUT57), .B1(new_n1159), .B2(new_n1192), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1221), .B1(new_n1280), .B2(new_n707), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1245), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1192), .A2(KEYINPUT126), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT126), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1189), .A2(new_n1191), .A3(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1283), .A2(new_n1005), .A3(new_n1285), .ZN(new_n1286));
  OAI211_X1 g1086(.A(new_n1286), .B(new_n1220), .C1(new_n978), .C2(new_n1193), .ZN(new_n1287));
  AOI22_X1  g1087(.A1(new_n1281), .A2(G378), .B1(new_n1282), .B2(new_n1287), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1277), .B1(new_n1288), .B2(new_n1272), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1156), .ZN(new_n1290));
  OAI211_X1 g1090(.A(new_n1197), .B(new_n1222), .C1(new_n1290), .C2(new_n1154), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1287), .A2(new_n1282), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1267), .A2(new_n1270), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1272), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1293), .A2(new_n1295), .A3(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(KEYINPUT62), .B1(new_n1289), .B2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT61), .ZN(new_n1299));
  AOI211_X1 g1099(.A(new_n1272), .B(new_n1294), .C1(new_n1291), .C2(new_n1292), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT62), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1299), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1262), .B1(new_n1298), .B2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1273), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1294), .A2(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(new_n1274), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1306), .B1(new_n1293), .B2(new_n1296), .ZN(new_n1307));
  OAI21_X1  g1107(.A(KEYINPUT63), .B1(new_n1307), .B2(new_n1300), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT63), .ZN(new_n1310));
  AOI21_X1  g1110(.A(KEYINPUT61), .B1(new_n1297), .B2(new_n1310), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1308), .A2(new_n1309), .A3(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1303), .A2(new_n1312), .ZN(G405));
  NAND2_X1  g1113(.A1(G375), .A2(new_n1282), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1314), .A2(new_n1291), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1262), .A2(new_n1315), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1309), .A2(new_n1291), .A3(new_n1314), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  XNOR2_X1  g1118(.A(new_n1318), .B(new_n1295), .ZN(G402));
endmodule


