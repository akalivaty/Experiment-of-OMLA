//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 1 0 1 1 0 0 0 0 1 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 0 1 1 0 1 0 0 1 1 0 1 0 0 0 1 1 0 1 0 1 0 0 0 0 0 0 1 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:03 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1241, new_n1242, new_n1243, new_n1244, new_n1245,
    new_n1246, new_n1247;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(new_n204));
  XOR2_X1   g0004(.A(new_n204), .B(KEYINPUT64), .Z(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  OAI21_X1  g0009(.A(G250), .B1(G257), .B2(G264), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  XOR2_X1   g0011(.A(KEYINPUT65), .B(KEYINPUT0), .Z(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(G58), .ZN(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(G50), .ZN(new_n220));
  OAI22_X1  g0020(.A1(new_n211), .A2(new_n212), .B1(new_n216), .B2(new_n220), .ZN(new_n221));
  AOI21_X1  g0021(.A(new_n221), .B1(new_n212), .B2(new_n211), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT66), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n207), .B1(new_n226), .B2(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT1), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n223), .A2(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G250), .B(G257), .Z(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT67), .ZN(new_n242));
  XOR2_X1   g0042(.A(G58), .B(G77), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G116), .Z(new_n245));
  XNOR2_X1  g0045(.A(G97), .B(G107), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  INV_X1    g0048(.A(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(KEYINPUT3), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT3), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G33), .ZN(new_n252));
  AND2_X1   g0052(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n253), .A2(G232), .A3(G1698), .ZN(new_n254));
  INV_X1    g0054(.A(G1698), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n253), .A2(G226), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G33), .A2(G97), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n254), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G274), .ZN(new_n261));
  INV_X1    g0061(.A(G41), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(KEYINPUT68), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT68), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G41), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G45), .ZN(new_n267));
  AOI211_X1 g0067(.A(G1), .B(new_n261), .C1(new_n266), .C2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n259), .ZN(new_n269));
  INV_X1    g0069(.A(G1), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n270), .B1(G41), .B2(G45), .ZN(new_n271));
  AND2_X1   g0071(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n268), .B1(G238), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n260), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(KEYINPUT13), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT73), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT13), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n260), .A2(new_n273), .A3(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n275), .A2(new_n276), .A3(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n274), .A2(KEYINPUT73), .A3(KEYINPUT13), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n279), .A2(G169), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(KEYINPUT14), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT14), .ZN(new_n283));
  NAND4_X1  g0083(.A1(new_n279), .A2(new_n283), .A3(G169), .A4(new_n280), .ZN(new_n284));
  AND2_X1   g0084(.A1(new_n275), .A2(new_n278), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G179), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n282), .A2(new_n284), .A3(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G13), .ZN(new_n288));
  NOR3_X1   g0088(.A1(new_n288), .A2(new_n214), .A3(G1), .ZN(new_n289));
  NAND3_X1  g0089(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(new_n213), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT70), .ZN(new_n293));
  XNOR2_X1  g0093(.A(new_n292), .B(new_n293), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n214), .A2(G1), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n294), .A2(G68), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n214), .A2(G33), .ZN(new_n298));
  INV_X1    g0098(.A(G77), .ZN(new_n299));
  OAI22_X1  g0099(.A1(new_n298), .A2(new_n299), .B1(new_n214), .B2(G68), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n214), .A2(new_n249), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n301), .A2(new_n202), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n291), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  XNOR2_X1  g0103(.A(KEYINPUT75), .B(KEYINPUT11), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  OR2_X1    g0105(.A1(new_n303), .A2(new_n304), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n289), .A2(new_n218), .ZN(new_n307));
  XNOR2_X1  g0107(.A(new_n307), .B(KEYINPUT12), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n297), .A2(new_n305), .A3(new_n306), .A4(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n279), .A2(G200), .A3(new_n280), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT74), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n279), .A2(KEYINPUT74), .A3(G200), .A4(new_n280), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n309), .B1(new_n285), .B2(G190), .ZN(new_n315));
  AOI22_X1  g0115(.A1(new_n287), .A2(new_n309), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(G200), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n250), .A2(new_n252), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n318), .A2(G1698), .ZN(new_n319));
  AOI22_X1  g0119(.A1(new_n319), .A2(G223), .B1(G33), .B2(G87), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n318), .A2(new_n255), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(G226), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(new_n259), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n268), .B1(G232), .B2(new_n272), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n317), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n324), .A2(new_n325), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n326), .B1(new_n328), .B2(G190), .ZN(new_n329));
  XOR2_X1   g0129(.A(KEYINPUT8), .B(G58), .Z(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n289), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n291), .A2(new_n295), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n333), .B1(new_n334), .B2(new_n331), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(KEYINPUT7), .B1(new_n318), .B2(new_n214), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT7), .ZN(new_n338));
  AOI211_X1 g0138(.A(new_n338), .B(G20), .C1(new_n250), .C2(new_n252), .ZN(new_n339));
  OAI21_X1  g0139(.A(G68), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(G58), .A2(G68), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n214), .B1(new_n219), .B2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(G159), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n301), .A2(new_n343), .ZN(new_n344));
  OAI21_X1  g0144(.A(KEYINPUT76), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n341), .ZN(new_n346));
  OAI21_X1  g0146(.A(G20), .B1(new_n346), .B2(new_n201), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT76), .ZN(new_n348));
  NOR2_X1   g0148(.A1(G20), .A2(G33), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(G159), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n347), .A2(new_n348), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n345), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n340), .A2(new_n352), .A3(KEYINPUT16), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(new_n291), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n340), .A2(new_n347), .A3(new_n350), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT16), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n336), .B1(new_n355), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n329), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(KEYINPUT17), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT17), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n329), .A2(new_n362), .A3(new_n359), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n355), .A2(new_n358), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(new_n335), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n327), .A2(G169), .ZN(new_n368));
  INV_X1    g0168(.A(G179), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n368), .B1(new_n369), .B2(new_n327), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n367), .A2(new_n370), .A3(KEYINPUT18), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT18), .ZN(new_n372));
  INV_X1    g0172(.A(G169), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n373), .B1(new_n324), .B2(new_n325), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n374), .B1(new_n328), .B2(G179), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n372), .B1(new_n375), .B2(new_n359), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n371), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n365), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n332), .A2(new_n202), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n380), .B1(new_n334), .B2(new_n202), .ZN(new_n381));
  XNOR2_X1  g0181(.A(new_n381), .B(KEYINPUT69), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n203), .A2(G20), .ZN(new_n383));
  INV_X1    g0183(.A(G150), .ZN(new_n384));
  OAI221_X1 g0184(.A(new_n383), .B1(new_n384), .B2(new_n301), .C1(new_n331), .C2(new_n298), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(new_n291), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n382), .A2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  OR2_X1    g0188(.A1(new_n388), .A2(KEYINPUT9), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n268), .B1(G226), .B2(new_n272), .ZN(new_n390));
  AOI22_X1  g0190(.A1(new_n321), .A2(G223), .B1(G77), .B2(new_n318), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n319), .A2(G222), .ZN(new_n392));
  AND2_X1   g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n390), .B1(new_n393), .B2(new_n269), .ZN(new_n394));
  INV_X1    g0194(.A(G190), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  XNOR2_X1  g0196(.A(KEYINPUT71), .B(G200), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n396), .B1(new_n397), .B2(new_n394), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n388), .A2(KEYINPUT9), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n389), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(KEYINPUT10), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT10), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n389), .A2(new_n398), .A3(new_n402), .A4(new_n399), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n394), .A2(G179), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n388), .B1(new_n373), .B2(new_n394), .ZN(new_n406));
  AOI22_X1  g0206(.A1(new_n401), .A2(new_n403), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  XNOR2_X1  g0207(.A(KEYINPUT68), .B(G41), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n270), .B(G274), .C1(new_n408), .C2(G45), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n269), .A2(new_n271), .ZN(new_n410));
  INV_X1    g0210(.A(G244), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n409), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  AOI22_X1  g0212(.A1(new_n321), .A2(G238), .B1(G107), .B2(new_n318), .ZN(new_n413));
  INV_X1    g0213(.A(G232), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n253), .A2(new_n255), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n413), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n412), .B1(new_n416), .B2(new_n259), .ZN(new_n417));
  AND2_X1   g0217(.A1(new_n417), .A2(G190), .ZN(new_n418));
  INV_X1    g0218(.A(new_n397), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  AOI22_X1  g0220(.A1(new_n330), .A2(new_n349), .B1(G20), .B2(G77), .ZN(new_n421));
  XNOR2_X1  g0221(.A(KEYINPUT15), .B(G87), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n421), .B1(new_n298), .B2(new_n422), .ZN(new_n423));
  AOI22_X1  g0223(.A1(new_n423), .A2(new_n291), .B1(new_n299), .B2(new_n289), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n294), .A2(G77), .A3(new_n296), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NOR3_X1   g0226(.A1(new_n418), .A2(new_n420), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n416), .A2(new_n259), .ZN(new_n428));
  INV_X1    g0228(.A(new_n412), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n430), .A2(G179), .ZN(new_n431));
  AOI22_X1  g0231(.A1(new_n430), .A2(new_n373), .B1(new_n425), .B2(new_n424), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT72), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n431), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n426), .B1(G169), .B2(new_n417), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(KEYINPUT72), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n427), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  AND4_X1   g0237(.A1(new_n316), .A2(new_n379), .A3(new_n407), .A4(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n321), .A2(G250), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n253), .A2(KEYINPUT4), .A3(G244), .A4(new_n255), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n250), .A2(new_n252), .A3(G244), .A4(new_n255), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT4), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(G33), .A2(G283), .ZN(new_n445));
  XNOR2_X1  g0245(.A(new_n445), .B(KEYINPUT77), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n440), .A2(new_n441), .A3(new_n444), .A4(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(new_n259), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT5), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n270), .B(G45), .C1(new_n449), .C2(G41), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n450), .B1(new_n408), .B2(new_n449), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n451), .A2(new_n259), .ZN(new_n452));
  AOI22_X1  g0252(.A1(new_n452), .A2(G257), .B1(G274), .B2(new_n451), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n448), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(G200), .ZN(new_n455));
  OAI21_X1  g0255(.A(G107), .B1(new_n337), .B2(new_n339), .ZN(new_n456));
  INV_X1    g0256(.A(G107), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n457), .A2(KEYINPUT6), .A3(G97), .ZN(new_n458));
  INV_X1    g0258(.A(new_n246), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n458), .B1(new_n459), .B2(KEYINPUT6), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(G20), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n349), .A2(G77), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n456), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(new_n291), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n332), .A2(G97), .ZN(new_n465));
  AOI211_X1 g0265(.A(new_n291), .B(new_n289), .C1(new_n270), .C2(G33), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n465), .B1(new_n466), .B2(G97), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n448), .A2(G190), .A3(new_n453), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n455), .A2(new_n464), .A3(new_n467), .A4(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n454), .A2(new_n373), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n464), .A2(new_n467), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n448), .A2(new_n369), .A3(new_n453), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n470), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  AND2_X1   g0273(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(G250), .ZN(new_n475));
  OAI21_X1  g0275(.A(KEYINPUT80), .B1(new_n415), .B2(new_n475), .ZN(new_n476));
  AOI22_X1  g0276(.A1(new_n321), .A2(G257), .B1(G33), .B2(G294), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT80), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n319), .A2(new_n478), .A3(G250), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n476), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(new_n259), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n451), .A2(G274), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n452), .A2(G264), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(G200), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n253), .A2(new_n214), .A3(G87), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(KEYINPUT22), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT22), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n253), .A2(new_n488), .A3(new_n214), .A4(G87), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT23), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n491), .B1(new_n214), .B2(G107), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n457), .A2(KEYINPUT23), .A3(G20), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(G33), .A2(G116), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n494), .B1(G20), .B2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n490), .A2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT24), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n496), .B1(new_n487), .B2(new_n489), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(KEYINPUT24), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n500), .A2(new_n291), .A3(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n289), .A2(KEYINPUT25), .A3(new_n457), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT25), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n505), .B1(new_n332), .B2(G107), .ZN(new_n506));
  AOI22_X1  g0306(.A1(new_n466), .A2(G107), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n480), .A2(new_n259), .B1(G264), .B2(new_n452), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n508), .A2(G190), .A3(new_n482), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n485), .A2(new_n503), .A3(new_n507), .A4(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n270), .A2(G45), .A3(G274), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n270), .A2(G45), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(G250), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n511), .B1(new_n259), .B2(new_n513), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n250), .A2(new_n252), .A3(G244), .A4(G1698), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n250), .A2(new_n252), .A3(G238), .A4(new_n255), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n515), .A2(new_n516), .A3(new_n495), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n514), .B1(new_n517), .B2(new_n259), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(G190), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT79), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n466), .A2(G87), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT19), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n214), .B1(new_n257), .B2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(G87), .ZN(new_n525));
  INV_X1    g0325(.A(G97), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n525), .A2(new_n526), .A3(new_n457), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n250), .A2(new_n252), .A3(new_n214), .A4(G68), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n523), .B1(new_n298), .B2(new_n526), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n531), .A2(new_n291), .B1(new_n289), .B2(new_n422), .ZN(new_n532));
  AND2_X1   g0332(.A1(new_n522), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n518), .A2(KEYINPUT79), .A3(G190), .ZN(new_n534));
  INV_X1    g0334(.A(new_n518), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n397), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n521), .A2(new_n533), .A3(new_n534), .A4(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n466), .ZN(new_n538));
  XOR2_X1   g0338(.A(new_n422), .B(KEYINPUT78), .Z(new_n539));
  OAI21_X1  g0339(.A(new_n532), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n518), .A2(new_n369), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n540), .B(new_n541), .C1(G169), .C2(new_n518), .ZN(new_n542));
  AND2_X1   g0342(.A1(new_n537), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n474), .A2(new_n510), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n484), .A2(new_n373), .ZN(new_n545));
  INV_X1    g0345(.A(new_n502), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n291), .B1(new_n501), .B2(KEYINPUT24), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n507), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n508), .A2(new_n369), .A3(new_n482), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n545), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n452), .A2(G270), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n250), .A2(new_n252), .A3(G257), .A4(new_n255), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n250), .A2(new_n252), .A3(G264), .A4(G1698), .ZN(new_n553));
  INV_X1    g0353(.A(G303), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n552), .B(new_n553), .C1(new_n253), .C2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n259), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n551), .A2(new_n482), .A3(new_n556), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n557), .A2(new_n369), .ZN(new_n558));
  INV_X1    g0358(.A(G116), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n559), .B1(new_n270), .B2(G33), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n292), .A2(new_n293), .ZN(new_n561));
  NOR3_X1   g0361(.A1(new_n289), .A2(new_n291), .A3(KEYINPUT70), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n289), .A2(new_n559), .ZN(new_n564));
  AOI21_X1  g0364(.A(G20), .B1(new_n249), .B2(G97), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n446), .A2(new_n565), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n291), .B1(new_n214), .B2(G116), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  AND3_X1   g0368(.A1(new_n566), .A2(new_n568), .A3(KEYINPUT20), .ZN(new_n569));
  AOI21_X1  g0369(.A(KEYINPUT20), .B1(new_n566), .B2(new_n568), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n563), .B(new_n564), .C1(new_n569), .C2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n558), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n571), .A2(KEYINPUT21), .A3(G169), .A4(new_n557), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n571), .B1(G200), .B2(new_n557), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n576), .B1(new_n395), .B2(new_n557), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n571), .A2(G169), .A3(new_n557), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT21), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n550), .A2(new_n575), .A3(new_n577), .A4(new_n580), .ZN(new_n581));
  NOR3_X1   g0381(.A1(new_n439), .A2(new_n544), .A3(new_n581), .ZN(G372));
  NAND2_X1  g0382(.A1(new_n314), .A2(new_n315), .ZN(new_n583));
  AND2_X1   g0383(.A1(new_n434), .A2(new_n436), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n287), .A2(new_n309), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n365), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  OR2_X1    g0387(.A1(new_n587), .A2(new_n378), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n401), .A2(new_n403), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n588), .A2(new_n589), .B1(new_n405), .B2(new_n406), .ZN(new_n590));
  AND3_X1   g0390(.A1(new_n470), .A2(new_n471), .A3(new_n472), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n543), .A2(new_n591), .A3(KEYINPUT26), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT26), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n537), .A2(new_n542), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n593), .B1(new_n594), .B2(new_n473), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n542), .ZN(new_n597));
  AND4_X1   g0397(.A1(new_n510), .A2(new_n473), .A3(new_n469), .A4(new_n543), .ZN(new_n598));
  AND2_X1   g0398(.A1(new_n557), .A2(G169), .ZN(new_n599));
  AOI21_X1  g0399(.A(KEYINPUT21), .B1(new_n599), .B2(new_n571), .ZN(new_n600));
  OAI21_X1  g0400(.A(KEYINPUT81), .B1(new_n574), .B2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT81), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n580), .A2(new_n602), .A3(new_n573), .A4(new_n572), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n601), .A2(new_n550), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n598), .A2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT82), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n597), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n598), .A2(new_n604), .A3(KEYINPUT82), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n438), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n590), .A2(new_n610), .ZN(G369));
  NOR2_X1   g0411(.A1(new_n288), .A2(G20), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n270), .ZN(new_n613));
  AND2_X1   g0413(.A1(new_n613), .A2(KEYINPUT27), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n613), .A2(KEYINPUT27), .ZN(new_n615));
  INV_X1    g0415(.A(G213), .ZN(new_n616));
  NOR3_X1   g0416(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  AND2_X1   g0417(.A1(new_n617), .A2(G343), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n571), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n619), .B1(new_n574), .B2(new_n600), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n601), .A2(new_n603), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n577), .B(new_n620), .C1(new_n621), .C2(new_n619), .ZN(new_n622));
  INV_X1    g0422(.A(G330), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n550), .A2(new_n618), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n548), .A2(new_n618), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n510), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n625), .B1(new_n550), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n624), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n618), .B1(new_n575), .B2(new_n580), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n625), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n629), .A2(new_n631), .ZN(G399));
  NOR2_X1   g0432(.A1(new_n527), .A2(G116), .ZN(new_n633));
  XOR2_X1   g0433(.A(new_n633), .B(KEYINPUT83), .Z(new_n634));
  NOR2_X1   g0434(.A1(new_n209), .A2(new_n408), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(G1), .ZN(new_n637));
  OAI22_X1  g0437(.A1(new_n634), .A2(new_n637), .B1(new_n220), .B2(new_n636), .ZN(new_n638));
  XNOR2_X1  g0438(.A(new_n638), .B(KEYINPUT28), .ZN(new_n639));
  NOR3_X1   g0439(.A1(new_n557), .A2(new_n535), .A3(new_n369), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n448), .A2(new_n453), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n640), .A2(new_n508), .A3(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT30), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n557), .A2(new_n369), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n484), .A2(new_n645), .A3(new_n454), .A4(new_n535), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n640), .A2(new_n641), .A3(KEYINPUT30), .A4(new_n508), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n644), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT31), .ZN(new_n649));
  AND3_X1   g0449(.A1(new_n648), .A2(new_n649), .A3(new_n618), .ZN(new_n650));
  AND3_X1   g0450(.A1(new_n550), .A2(new_n575), .A3(new_n580), .ZN(new_n651));
  INV_X1    g0451(.A(new_n618), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n598), .A2(new_n651), .A3(new_n577), .A4(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n649), .B1(new_n648), .B2(new_n618), .ZN(new_n654));
  AOI211_X1 g0454(.A(new_n623), .B(new_n650), .C1(new_n653), .C2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n609), .A2(new_n652), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT29), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  OR2_X1    g0458(.A1(new_n544), .A2(new_n651), .ZN(new_n659));
  INV_X1    g0459(.A(new_n597), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n618), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(KEYINPUT29), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n655), .B1(new_n658), .B2(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n639), .B1(new_n663), .B2(G1), .ZN(G364));
  NOR2_X1   g0464(.A1(G13), .A2(G33), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n666), .A2(G20), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n213), .B1(G20), .B2(new_n373), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n253), .A2(new_n208), .ZN(new_n670));
  XNOR2_X1  g0470(.A(new_n670), .B(KEYINPUT84), .ZN(new_n671));
  XOR2_X1   g0471(.A(G355), .B(KEYINPUT85), .Z(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n673), .B1(G116), .B2(new_n208), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(KEYINPUT86), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n244), .A2(new_n267), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n253), .A2(new_n209), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n677), .B1(G45), .B2(new_n220), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n675), .B1(new_n676), .B2(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n674), .A2(KEYINPUT86), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n669), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n270), .B1(new_n612), .B2(G45), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n635), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n214), .A2(new_n395), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT87), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n369), .A2(G200), .ZN(new_n688));
  AND3_X1   g0488(.A1(new_n686), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n687), .B1(new_n686), .B2(new_n688), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(G322), .ZN(new_n693));
  INV_X1    g0493(.A(G283), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n214), .A2(G190), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n397), .A2(new_n369), .A3(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n397), .A2(new_n369), .A3(new_n686), .ZN(new_n697));
  OAI221_X1 g0497(.A(new_n693), .B1(new_n694), .B2(new_n696), .C1(new_n554), .C2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n695), .A2(new_n688), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(G179), .A2(G200), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n695), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  AOI22_X1  g0503(.A1(G311), .A2(new_n700), .B1(new_n703), .B2(G329), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n369), .A2(new_n317), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(new_n686), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  XOR2_X1   g0507(.A(KEYINPUT89), .B(G326), .Z(new_n708));
  AOI21_X1  g0508(.A(new_n253), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n705), .A2(new_n695), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(G317), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(KEYINPUT33), .ZN(new_n713));
  OR2_X1    g0513(.A1(new_n712), .A2(KEYINPUT33), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n711), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n214), .B1(new_n701), .B2(G190), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(G294), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n704), .A2(new_n709), .A3(new_n715), .A4(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n697), .ZN(new_n720));
  AOI22_X1  g0520(.A1(new_n692), .A2(G58), .B1(G87), .B2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n696), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(G107), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n318), .B1(new_n711), .B2(G68), .ZN(new_n724));
  AOI22_X1  g0524(.A1(G50), .A2(new_n707), .B1(new_n700), .B2(G77), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n721), .A2(new_n723), .A3(new_n724), .A4(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n702), .A2(new_n343), .ZN(new_n727));
  XOR2_X1   g0527(.A(KEYINPUT88), .B(KEYINPUT32), .Z(new_n728));
  XNOR2_X1  g0528(.A(new_n727), .B(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n729), .B1(new_n526), .B2(new_n716), .ZN(new_n730));
  OAI22_X1  g0530(.A1(new_n698), .A2(new_n719), .B1(new_n726), .B2(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n685), .B1(new_n731), .B2(new_n668), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n681), .A2(new_n732), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n733), .B1(new_n622), .B2(new_n667), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n624), .A2(new_n684), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n622), .A2(new_n623), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n734), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(G396));
  AOI21_X1  g0538(.A(new_n618), .B1(new_n607), .B2(new_n608), .ZN(new_n739));
  INV_X1    g0539(.A(new_n431), .ZN(new_n740));
  OAI211_X1 g0540(.A(new_n426), .B(new_n433), .C1(G169), .C2(new_n417), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n426), .A2(new_n618), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  AND4_X1   g0543(.A1(new_n436), .A2(new_n740), .A3(new_n741), .A4(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n744), .B1(new_n437), .B2(new_n742), .ZN(new_n745));
  XNOR2_X1  g0545(.A(new_n739), .B(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n684), .B1(new_n746), .B2(new_n655), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n747), .B1(new_n655), .B2(new_n746), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n668), .A2(new_n665), .ZN(new_n749));
  XOR2_X1   g0549(.A(new_n749), .B(KEYINPUT90), .Z(new_n750));
  OAI21_X1  g0550(.A(new_n684), .B1(new_n750), .B2(G77), .ZN(new_n751));
  INV_X1    g0551(.A(G311), .ZN(new_n752));
  OAI22_X1  g0552(.A1(new_n710), .A2(new_n694), .B1(new_n702), .B2(new_n752), .ZN(new_n753));
  OAI221_X1 g0553(.A(new_n318), .B1(new_n716), .B2(new_n526), .C1(new_n706), .C2(new_n554), .ZN(new_n754));
  AOI211_X1 g0554(.A(new_n753), .B(new_n754), .C1(G116), .C2(new_n700), .ZN(new_n755));
  AOI22_X1  g0555(.A1(G87), .A2(new_n722), .B1(new_n720), .B2(G107), .ZN(new_n756));
  INV_X1    g0556(.A(G294), .ZN(new_n757));
  OAI211_X1 g0557(.A(new_n755), .B(new_n756), .C1(new_n757), .C2(new_n691), .ZN(new_n758));
  AOI22_X1  g0558(.A1(G137), .A2(new_n707), .B1(new_n700), .B2(G159), .ZN(new_n759));
  INV_X1    g0559(.A(G143), .ZN(new_n760));
  OAI221_X1 g0560(.A(new_n759), .B1(new_n384), .B2(new_n710), .C1(new_n760), .C2(new_n691), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  XNOR2_X1  g0562(.A(KEYINPUT91), .B(KEYINPUT34), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n696), .A2(new_n218), .ZN(new_n765));
  INV_X1    g0565(.A(G132), .ZN(new_n766));
  OAI221_X1 g0566(.A(new_n253), .B1(new_n716), .B2(new_n217), .C1(new_n766), .C2(new_n702), .ZN(new_n767));
  AOI211_X1 g0567(.A(new_n765), .B(new_n767), .C1(G50), .C2(new_n720), .ZN(new_n768));
  INV_X1    g0568(.A(new_n763), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n768), .B1(new_n761), .B2(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n758), .B1(new_n764), .B2(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n751), .B1(new_n771), .B2(new_n668), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n437), .A2(new_n742), .ZN(new_n773));
  INV_X1    g0573(.A(new_n744), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n772), .B1(new_n775), .B2(new_n666), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n748), .A2(new_n776), .ZN(G384));
  XNOR2_X1  g0577(.A(new_n460), .B(KEYINPUT92), .ZN(new_n778));
  INV_X1    g0578(.A(KEYINPUT35), .ZN(new_n779));
  AOI211_X1 g0579(.A(new_n559), .B(new_n216), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n780), .B1(new_n779), .B2(new_n778), .ZN(new_n781));
  INV_X1    g0581(.A(KEYINPUT36), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n341), .A2(G77), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n220), .A2(new_n783), .B1(G50), .B2(new_n218), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n270), .A2(G13), .ZN(new_n785));
  AOI22_X1  g0585(.A1(new_n781), .A2(new_n782), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(KEYINPUT16), .B1(new_n340), .B2(new_n352), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n335), .B1(new_n354), .B2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(KEYINPUT94), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  OAI211_X1 g0590(.A(KEYINPUT94), .B(new_n335), .C1(new_n354), .C2(new_n787), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n790), .A2(new_n617), .A3(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(KEYINPUT95), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND4_X1  g0594(.A1(new_n790), .A2(KEYINPUT95), .A3(new_n617), .A4(new_n791), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n370), .A2(new_n790), .A3(new_n791), .ZN(new_n796));
  NAND4_X1  g0596(.A1(new_n794), .A2(new_n360), .A3(new_n795), .A4(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(KEYINPUT37), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n367), .A2(new_n370), .ZN(new_n799));
  XOR2_X1   g0599(.A(new_n617), .B(KEYINPUT96), .Z(new_n800));
  NAND2_X1  g0600(.A1(new_n367), .A2(new_n800), .ZN(new_n801));
  XOR2_X1   g0601(.A(KEYINPUT97), .B(KEYINPUT37), .Z(new_n802));
  AND4_X1   g0602(.A1(new_n799), .A2(new_n801), .A3(new_n360), .A4(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n798), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n794), .A2(new_n795), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n806), .B1(new_n365), .B2(new_n378), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n805), .A2(KEYINPUT38), .A3(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(KEYINPUT98), .ZN(new_n809));
  INV_X1    g0609(.A(KEYINPUT38), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n803), .B1(new_n797), .B2(KEYINPUT37), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n364), .A2(new_n377), .B1(new_n794), .B2(new_n795), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n810), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n808), .A2(new_n809), .A3(new_n813), .ZN(new_n814));
  NAND4_X1  g0614(.A1(new_n805), .A2(KEYINPUT98), .A3(new_n807), .A4(KEYINPUT38), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(KEYINPUT99), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n584), .A2(new_n652), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n820), .B1(new_n739), .B2(new_n775), .ZN(new_n821));
  AND2_X1   g0621(.A1(new_n281), .A2(KEYINPUT14), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n284), .A2(new_n286), .ZN(new_n823));
  OAI211_X1 g0623(.A(new_n309), .B(new_n618), .C1(new_n822), .C2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(KEYINPUT93), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND4_X1  g0626(.A1(new_n287), .A2(KEYINPUT93), .A3(new_n309), .A4(new_n618), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n309), .A2(new_n618), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n826), .A2(new_n827), .B1(new_n316), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n821), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n814), .A2(KEYINPUT99), .A3(new_n815), .ZN(new_n831));
  AND3_X1   g0631(.A1(new_n818), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n377), .A2(new_n800), .ZN(new_n833));
  OAI21_X1  g0633(.A(KEYINPUT100), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n814), .A2(KEYINPUT39), .A3(new_n815), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n379), .A2(new_n801), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n799), .A2(new_n801), .A3(new_n360), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(new_n802), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n810), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT39), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n839), .A2(new_n840), .A3(new_n808), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n835), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n586), .A2(new_n618), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n818), .A2(new_n830), .A3(new_n831), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT100), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n848), .B(new_n849), .C1(new_n377), .C2(new_n800), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n834), .A2(new_n847), .A3(new_n850), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n658), .A2(new_n438), .A3(new_n662), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(new_n590), .ZN(new_n853));
  XOR2_X1   g0653(.A(new_n851), .B(new_n853), .Z(new_n854));
  NAND2_X1  g0654(.A1(new_n839), .A2(new_n808), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n826), .A2(new_n827), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n316), .A2(new_n828), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n650), .ZN(new_n859));
  NOR3_X1   g0659(.A1(new_n544), .A2(new_n581), .A3(new_n618), .ZN(new_n860));
  INV_X1    g0660(.A(new_n654), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n775), .B(new_n859), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  NAND4_X1  g0663(.A1(new_n855), .A2(KEYINPUT40), .A3(new_n858), .A4(new_n863), .ZN(new_n864));
  AND3_X1   g0664(.A1(new_n814), .A2(KEYINPUT99), .A3(new_n815), .ZN(new_n865));
  AOI21_X1  g0665(.A(KEYINPUT99), .B1(new_n814), .B2(new_n815), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT101), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n863), .A2(new_n858), .A3(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(KEYINPUT101), .B1(new_n829), .B2(new_n862), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NOR3_X1   g0670(.A1(new_n865), .A2(new_n866), .A3(new_n870), .ZN(new_n871));
  OAI211_X1 g0671(.A(G330), .B(new_n864), .C1(new_n871), .C2(KEYINPUT40), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n438), .A2(new_n655), .ZN(new_n873));
  INV_X1    g0673(.A(new_n864), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n867), .B1(new_n863), .B2(new_n858), .ZN(new_n875));
  NOR3_X1   g0675(.A1(new_n829), .A2(new_n862), .A3(KEYINPUT101), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n818), .A2(new_n831), .A3(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT40), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n874), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n653), .A2(new_n654), .ZN(new_n881));
  AND3_X1   g0681(.A1(new_n438), .A2(new_n881), .A3(new_n859), .ZN(new_n882));
  AOI22_X1  g0682(.A1(new_n872), .A2(new_n873), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(KEYINPUT102), .B1(new_n854), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n854), .A2(new_n883), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n884), .B(new_n885), .C1(new_n270), .C2(new_n612), .ZN(new_n886));
  NOR3_X1   g0686(.A1(new_n854), .A2(KEYINPUT102), .A3(new_n883), .ZN(new_n887));
  OAI221_X1 g0687(.A(new_n786), .B1(new_n782), .B2(new_n781), .C1(new_n886), .C2(new_n887), .ZN(G367));
  INV_X1    g0688(.A(new_n677), .ZN(new_n889));
  OAI221_X1 g0689(.A(new_n669), .B1(new_n208), .B2(new_n422), .C1(new_n239), .C2(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n685), .B1(new_n890), .B2(KEYINPUT109), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n891), .B1(KEYINPUT109), .B2(new_n890), .ZN(new_n892));
  AOI22_X1  g0692(.A1(G50), .A2(new_n700), .B1(new_n703), .B2(G137), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n893), .B1(new_n760), .B2(new_n706), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n716), .A2(new_n218), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n253), .B1(new_n710), .B2(new_n343), .ZN(new_n896));
  NOR3_X1   g0696(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  AOI22_X1  g0697(.A1(G58), .A2(new_n720), .B1(new_n722), .B2(G77), .ZN(new_n898));
  OAI211_X1 g0698(.A(new_n897), .B(new_n898), .C1(new_n384), .C2(new_n691), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n899), .B(KEYINPUT110), .ZN(new_n900));
  OAI22_X1  g0700(.A1(new_n706), .A2(new_n752), .B1(new_n710), .B2(new_n757), .ZN(new_n901));
  OAI221_X1 g0701(.A(new_n318), .B1(new_n716), .B2(new_n457), .C1(new_n694), .C2(new_n699), .ZN(new_n902));
  AOI211_X1 g0702(.A(new_n901), .B(new_n902), .C1(G317), .C2(new_n703), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n696), .A2(new_n526), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n904), .B1(new_n692), .B2(G303), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT46), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n906), .B1(new_n697), .B2(new_n559), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n720), .A2(KEYINPUT46), .A3(G116), .ZN(new_n908));
  NAND4_X1  g0708(.A1(new_n903), .A2(new_n905), .A3(new_n907), .A4(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(KEYINPUT47), .B1(new_n900), .B2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n668), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n900), .A2(KEYINPUT47), .A3(new_n909), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n892), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n652), .A2(new_n533), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(new_n542), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n917), .B1(new_n543), .B2(new_n916), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n918), .B(KEYINPUT103), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n915), .B1(new_n667), .B2(new_n919), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n682), .B(KEYINPUT108), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n471), .A2(new_n618), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n474), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n591), .A2(new_n618), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n631), .A2(new_n926), .ZN(new_n927));
  XOR2_X1   g0727(.A(new_n927), .B(KEYINPUT45), .Z(new_n928));
  XOR2_X1   g0728(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  OR3_X1    g0730(.A1(new_n631), .A2(new_n926), .A3(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n930), .B1(new_n631), .B2(new_n926), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n928), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n629), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND4_X1  g0735(.A1(new_n928), .A2(new_n629), .A3(new_n931), .A4(new_n932), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n628), .B(new_n630), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n938), .B(new_n624), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n663), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n663), .B1(new_n937), .B2(new_n940), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n635), .B(KEYINPUT41), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n922), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT106), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n628), .A2(new_n630), .ZN(new_n946));
  OAI21_X1  g0746(.A(KEYINPUT42), .B1(new_n946), .B2(new_n924), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n473), .B1(new_n924), .B2(new_n550), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(new_n652), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT105), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OR3_X1    g0752(.A1(new_n946), .A2(KEYINPUT42), .A3(new_n924), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n950), .A2(new_n951), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(KEYINPUT104), .A2(KEYINPUT43), .ZN(new_n957));
  AND2_X1   g0757(.A1(KEYINPUT104), .A2(KEYINPUT43), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n919), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n956), .A2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT43), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n959), .B1(new_n961), .B2(new_n919), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n954), .B2(new_n955), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n960), .A2(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(new_n926), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n629), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n945), .B1(new_n964), .B2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(new_n966), .ZN(new_n968));
  NAND4_X1  g0768(.A1(new_n960), .A2(KEYINPUT106), .A3(new_n968), .A4(new_n963), .ZN(new_n969));
  AOI22_X1  g0769(.A1(new_n967), .A2(new_n969), .B1(new_n966), .B2(new_n964), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n920), .B1(new_n944), .B2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(G387));
  NAND2_X1  g0772(.A1(new_n939), .A2(new_n922), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n671), .A2(new_n634), .B1(new_n457), .B2(new_n209), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n974), .B(KEYINPUT111), .Z(new_n975));
  OAI21_X1  g0775(.A(new_n267), .B1(new_n218), .B2(new_n299), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n330), .A2(new_n202), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n976), .B1(new_n977), .B2(KEYINPUT50), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(KEYINPUT50), .B2(new_n977), .ZN(new_n979));
  OAI221_X1 g0779(.A(new_n677), .B1(new_n634), .B2(new_n979), .C1(new_n236), .C2(new_n267), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n975), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n685), .B1(new_n981), .B2(new_n669), .ZN(new_n982));
  INV_X1    g0782(.A(new_n667), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n706), .A2(new_n343), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT113), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n318), .B1(new_n711), .B2(new_n330), .ZN(new_n986));
  XNOR2_X1  g0786(.A(KEYINPUT112), .B(G150), .ZN(new_n987));
  AOI22_X1  g0787(.A1(G68), .A2(new_n700), .B1(new_n703), .B2(new_n987), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n985), .A2(new_n986), .A3(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n539), .A2(new_n716), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n691), .A2(new_n202), .B1(new_n299), .B2(new_n697), .ZN(new_n991));
  NOR4_X1   g0791(.A1(new_n989), .A2(new_n904), .A3(new_n990), .A4(new_n991), .ZN(new_n992));
  AOI22_X1  g0792(.A1(G322), .A2(new_n707), .B1(new_n700), .B2(G303), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n993), .B1(new_n752), .B2(new_n710), .C1(new_n712), .C2(new_n691), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT48), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n995), .B1(new_n694), .B2(new_n716), .C1(new_n757), .C2(new_n697), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT49), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n253), .B1(new_n703), .B2(new_n708), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n559), .B2(new_n696), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n1000), .B1(new_n996), .B2(new_n997), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n992), .B1(new_n998), .B2(new_n1001), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n982), .B1(new_n628), .B2(new_n983), .C1(new_n1002), .C2(new_n911), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n663), .A2(new_n939), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT114), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1006), .A2(new_n635), .A3(new_n940), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1008));
  OAI211_X1 g0808(.A(new_n973), .B(new_n1003), .C1(new_n1007), .C2(new_n1008), .ZN(G393));
  INV_X1    g0809(.A(KEYINPUT115), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n935), .A2(new_n1010), .A3(new_n936), .ZN(new_n1011));
  OR3_X1    g0811(.A1(new_n933), .A2(new_n1010), .A3(new_n934), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(new_n922), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT118), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n965), .A2(new_n667), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n247), .A2(new_n889), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n669), .B1(new_n526), .B2(new_n208), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n684), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n691), .A2(new_n343), .B1(new_n384), .B2(new_n706), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT51), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n253), .B1(new_n710), .B2(new_n202), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n331), .A2(new_n699), .B1(new_n760), .B2(new_n702), .ZN(new_n1023));
  AOI211_X1 g0823(.A(new_n1022), .B(new_n1023), .C1(G77), .C2(new_n717), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(G68), .A2(new_n720), .B1(new_n722), .B2(G87), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1021), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n691), .A2(new_n752), .B1(new_n712), .B2(new_n706), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n1027), .B(KEYINPUT52), .Z(new_n1028));
  XNOR2_X1  g0828(.A(KEYINPUT116), .B(KEYINPUT117), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n723), .B1(new_n694), .B2(new_n697), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(G303), .A2(new_n711), .B1(new_n703), .B2(G322), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1032), .B(new_n318), .C1(new_n757), .C2(new_n699), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n1031), .B(new_n1033), .C1(G116), .C2(new_n717), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1030), .A2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1026), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1019), .B1(new_n1037), .B2(new_n668), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1016), .A2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1014), .A2(new_n1015), .A3(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n921), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n1039), .ZN(new_n1042));
  OAI21_X1  g0842(.A(KEYINPUT118), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1011), .A2(new_n1012), .A3(new_n940), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n937), .A2(new_n940), .ZN(new_n1045));
  NOR3_X1   g0845(.A1(new_n1045), .A2(new_n209), .A3(new_n408), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n1040), .A2(new_n1043), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n1047), .ZN(G390));
  OAI21_X1  g0848(.A(new_n845), .B1(new_n821), .B2(new_n829), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1049), .A2(new_n835), .A3(new_n841), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n829), .B(KEYINPUT119), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n820), .B1(new_n661), .B2(new_n775), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n845), .B(new_n855), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1053));
  AND4_X1   g0853(.A1(G330), .A2(new_n881), .A3(new_n859), .A4(new_n775), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1054), .A2(new_n858), .ZN(new_n1055));
  AND3_X1   g0855(.A1(new_n1050), .A2(new_n1053), .A3(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1055), .B1(new_n1050), .B2(new_n1053), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n843), .A2(new_n665), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n684), .B1(new_n750), .B2(new_n330), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n699), .A2(new_n526), .B1(new_n702), .B2(new_n757), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n318), .B1(new_n716), .B2(new_n299), .C1(new_n706), .C2(new_n694), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n1061), .B(new_n1062), .C1(G107), .C2(new_n711), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n765), .B1(G87), .B2(new_n720), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n1063), .B(new_n1064), .C1(new_n559), .C2(new_n691), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n720), .A2(new_n987), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT53), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n711), .A2(G137), .ZN(new_n1068));
  INV_X1    g0868(.A(G128), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(KEYINPUT54), .B(G143), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n1068), .B1(new_n1069), .B2(new_n706), .C1(new_n699), .C2(new_n1070), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n691), .A2(new_n766), .B1(new_n202), .B2(new_n696), .ZN(new_n1072));
  INV_X1    g0872(.A(G125), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n253), .B1(new_n716), .B2(new_n343), .C1(new_n1073), .C2(new_n702), .ZN(new_n1074));
  OR3_X1    g0874(.A1(new_n1071), .A2(new_n1072), .A3(new_n1074), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1065), .B1(new_n1067), .B2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1060), .B1(new_n1076), .B2(new_n668), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n1058), .A2(new_n922), .B1(new_n1059), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(KEYINPUT120), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n655), .A2(new_n775), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1051), .A2(new_n1080), .ZN(new_n1081));
  AND2_X1   g0881(.A1(new_n1055), .A2(new_n1052), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1080), .A2(new_n829), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(new_n1055), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n821), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n1081), .A2(new_n1082), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n852), .A2(new_n590), .A3(new_n873), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n636), .B1(new_n1058), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1087), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1079), .B1(new_n1089), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1050), .A2(new_n1053), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1055), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1050), .A2(new_n1055), .A3(new_n1053), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1099), .A2(new_n1088), .A3(new_n1100), .ZN(new_n1101));
  AND4_X1   g0901(.A1(new_n1079), .A2(new_n1095), .A3(new_n1101), .A4(new_n635), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1078), .B1(new_n1096), .B2(new_n1102), .ZN(G378));
  NAND2_X1  g0903(.A1(new_n878), .A2(new_n879), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n407), .A2(KEYINPUT122), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n407), .A2(KEYINPUT122), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n387), .B(new_n617), .C1(new_n1106), .C2(new_n1107), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1107), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n387), .A2(new_n617), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1110), .A2(new_n1111), .A3(new_n1105), .ZN(new_n1112));
  AND3_X1   g0912(.A1(new_n1108), .A2(new_n1109), .A3(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1109), .B1(new_n1108), .B2(new_n1112), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(new_n1116));
  AND4_X1   g0916(.A1(G330), .A2(new_n1104), .A3(new_n864), .A4(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1116), .B1(new_n880), .B2(G330), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n851), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n872), .A2(new_n1115), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n865), .A2(new_n866), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n833), .B1(new_n1121), .B2(new_n830), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n846), .B1(new_n1122), .B2(new_n849), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n1104), .A2(new_n1116), .A3(G330), .A4(new_n864), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1120), .A2(new_n1123), .A3(new_n834), .A4(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1119), .A2(new_n922), .A3(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n685), .B1(new_n202), .B2(new_n749), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(new_n1127), .B(KEYINPUT121), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n716), .A2(new_n384), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n706), .A2(new_n1073), .B1(new_n710), .B2(new_n766), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n1129), .B(new_n1130), .C1(G137), .C2(new_n700), .ZN(new_n1131));
  OAI221_X1 g0931(.A(new_n1131), .B1(new_n1069), .B2(new_n691), .C1(new_n697), .C2(new_n1070), .ZN(new_n1132));
  OR2_X1    g0932(.A1(new_n1132), .A2(KEYINPUT59), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(KEYINPUT59), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n722), .A2(G159), .ZN(new_n1135));
  AOI211_X1 g0935(.A(G33), .B(G41), .C1(new_n703), .C2(G124), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n1133), .A2(new_n1134), .A3(new_n1135), .A4(new_n1136), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n692), .A2(G107), .B1(G77), .B2(new_n720), .ZN(new_n1138));
  OAI221_X1 g0938(.A(new_n1138), .B1(new_n217), .B2(new_n696), .C1(new_n539), .C2(new_n699), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n706), .A2(new_n559), .B1(new_n710), .B2(new_n526), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n318), .B(new_n266), .C1(new_n702), .C2(new_n694), .ZN(new_n1141));
  NOR4_X1   g0941(.A1(new_n1139), .A2(new_n895), .A3(new_n1140), .A4(new_n1141), .ZN(new_n1142));
  OR2_X1    g0942(.A1(new_n1142), .A2(KEYINPUT58), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1142), .A2(KEYINPUT58), .ZN(new_n1144));
  OAI221_X1 g0944(.A(new_n202), .B1(G33), .B2(G41), .C1(new_n253), .C2(new_n408), .ZN(new_n1145));
  AND4_X1   g0945(.A1(new_n1137), .A2(new_n1143), .A3(new_n1144), .A4(new_n1145), .ZN(new_n1146));
  OAI221_X1 g0946(.A(new_n1128), .B1(new_n911), .B2(new_n1146), .C1(new_n1115), .C2(new_n666), .ZN(new_n1147));
  AND2_X1   g0947(.A1(new_n1126), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1101), .A2(new_n1093), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1119), .A2(new_n1125), .A3(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(KEYINPUT57), .ZN(new_n1151));
  AND2_X1   g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n1119), .A2(new_n1125), .A3(KEYINPUT57), .A4(new_n1149), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n635), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1148), .B1(new_n1152), .B2(new_n1154), .ZN(G375));
  NAND2_X1  g0955(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1094), .A2(new_n942), .A3(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n990), .B1(G77), .B2(new_n722), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n318), .B1(new_n706), .B2(new_n757), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n710), .A2(new_n559), .B1(new_n702), .B2(new_n554), .ZN(new_n1160));
  AOI211_X1 g0960(.A(new_n1159), .B(new_n1160), .C1(G107), .C2(new_n700), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n692), .A2(G283), .B1(G97), .B2(new_n720), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1158), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n692), .A2(G137), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(G58), .A2(new_n722), .B1(new_n720), .B2(G159), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n710), .A2(new_n1070), .B1(new_n702), .B2(new_n1069), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1166), .B1(G132), .B2(new_n707), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n253), .B1(new_n699), .B2(new_n384), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1168), .B1(G50), .B2(new_n717), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n1164), .A2(new_n1165), .A3(new_n1167), .A4(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n911), .B1(new_n1163), .B2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n684), .B1(new_n750), .B2(G68), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n1171), .B(new_n1172), .C1(new_n1051), .C2(new_n665), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(new_n1092), .B2(new_n922), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1157), .A2(new_n1174), .ZN(G381));
  NAND2_X1  g0975(.A1(new_n1089), .A2(new_n1095), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(new_n1078), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(G375), .A2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n971), .A2(new_n1047), .ZN(new_n1179));
  OR2_X1    g0979(.A1(G393), .A2(G396), .ZN(new_n1180));
  NOR4_X1   g0980(.A1(new_n1179), .A2(G384), .A3(G381), .A4(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1178), .A2(new_n1181), .ZN(G407));
  NOR2_X1   g0982(.A1(new_n616), .A2(G343), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1178), .A2(new_n1183), .ZN(new_n1184));
  OR2_X1    g0984(.A1(new_n1184), .A2(KEYINPUT123), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(KEYINPUT123), .ZN(new_n1186));
  NAND4_X1  g0986(.A1(new_n1185), .A2(G213), .A3(G407), .A4(new_n1186), .ZN(G409));
  XNOR2_X1  g0987(.A(G393), .B(new_n737), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT127), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1179), .A2(new_n1189), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n971), .A2(new_n1047), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1188), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT61), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(G387), .A2(G390), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1188), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1194), .A2(new_n1179), .A3(new_n1195), .A4(new_n1189), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1192), .A2(new_n1193), .A3(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT124), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT60), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n635), .B(new_n1094), .C1(new_n1199), .C2(new_n1200), .ZN(new_n1201));
  AND2_X1   g1001(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1174), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(G384), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  OAI211_X1 g1005(.A(G384), .B(new_n1174), .C1(new_n1201), .C2(new_n1202), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1183), .A2(KEYINPUT125), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1183), .A2(G2897), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1208), .A2(new_n1210), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .A4(new_n1209), .ZN(new_n1212));
  AND3_X1   g1012(.A1(new_n1211), .A2(KEYINPUT126), .A3(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(KEYINPUT126), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  OAI211_X1 g1015(.A(G378), .B(new_n1148), .C1(new_n1152), .C2(new_n1154), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n942), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1126), .B(new_n1147), .C1(new_n1150), .C2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1177), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1216), .A2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1183), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1197), .B1(new_n1215), .B2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1225));
  NOR3_X1   g1025(.A1(new_n1223), .A2(KEYINPUT63), .A3(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT63), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1183), .B1(new_n1216), .B2(new_n1220), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1225), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1227), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1224), .B1(new_n1226), .B2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT62), .ZN(new_n1232));
  AND3_X1   g1032(.A1(new_n1228), .A2(new_n1232), .A3(new_n1229), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1193), .B1(new_n1228), .B2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1232), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1236));
  NOR3_X1   g1036(.A1(new_n1233), .A2(new_n1235), .A3(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1192), .A2(new_n1196), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1231), .B1(new_n1237), .B2(new_n1239), .ZN(G405));
  NAND2_X1  g1040(.A1(G375), .A2(new_n1219), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(new_n1216), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1239), .A2(new_n1242), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1238), .A2(new_n1216), .A3(new_n1241), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(new_n1225), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1243), .A2(new_n1229), .A3(new_n1244), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(G402));
endmodule


