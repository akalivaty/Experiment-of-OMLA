//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 0 1 0 1 1 0 1 1 1 0 1 0 0 0 1 0 1 0 0 1 1 0 1 1 0 0 0 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:01 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n224,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1258, new_n1259, new_n1260, new_n1261,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XOR2_X1   g0007(.A(new_n207), .B(KEYINPUT0), .Z(new_n208));
  AOI22_X1  g0008(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n210));
  NAND3_X1  g0010(.A1(new_n209), .A2(new_n210), .A3(KEYINPUT65), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n213));
  NAND3_X1  g0013(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  AOI21_X1  g0014(.A(KEYINPUT65), .B1(new_n209), .B2(new_n210), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n205), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT1), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  INV_X1    g0018(.A(G20), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n202), .A2(G50), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT64), .Z(new_n222));
  AOI211_X1 g0022(.A(new_n208), .B(new_n217), .C1(new_n220), .C2(new_n222), .ZN(G361));
  XOR2_X1   g0023(.A(G250), .B(G257), .Z(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(G270), .ZN(new_n225));
  XOR2_X1   g0025(.A(KEYINPUT67), .B(G264), .Z(new_n226));
  XNOR2_X1  g0026(.A(new_n225), .B(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n228));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G226), .B(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n227), .B(new_n232), .Z(G358));
  XOR2_X1   g0033(.A(G87), .B(G116), .Z(new_n234));
  XNOR2_X1  g0034(.A(G97), .B(G107), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G50), .B(G68), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G58), .B(G77), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n236), .B(new_n239), .Z(G351));
  INV_X1    g0040(.A(G1), .ZN(new_n241));
  NAND3_X1  g0041(.A1(new_n241), .A2(G13), .A3(G20), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n242), .A2(KEYINPUT70), .ZN(new_n243));
  INV_X1    g0043(.A(KEYINPUT70), .ZN(new_n244));
  NAND4_X1  g0044(.A1(new_n244), .A2(new_n241), .A3(G13), .A4(G20), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  NOR2_X1   g0046(.A1(new_n246), .A2(G97), .ZN(new_n247));
  NAND3_X1  g0047(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(new_n218), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n241), .A2(G33), .ZN(new_n251));
  AND3_X1   g0051(.A1(new_n246), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n247), .B1(new_n252), .B2(G97), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G107), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G97), .ZN(new_n256));
  INV_X1    g0056(.A(G97), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G107), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT6), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n256), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n255), .A2(KEYINPUT6), .A3(G97), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G20), .ZN(new_n263));
  NOR2_X1   g0063(.A1(G20), .A2(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G77), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT7), .ZN(new_n267));
  XNOR2_X1  g0067(.A(KEYINPUT3), .B(G33), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n267), .B1(new_n268), .B2(G20), .ZN(new_n269));
  INV_X1    g0069(.A(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(KEYINPUT3), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT3), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n274), .A2(KEYINPUT7), .A3(new_n219), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n255), .B1(new_n269), .B2(new_n275), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n249), .B1(new_n266), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(KEYINPUT76), .ZN(new_n278));
  AOI21_X1  g0078(.A(KEYINPUT7), .B1(new_n274), .B2(new_n219), .ZN(new_n279));
  AOI211_X1 g0079(.A(new_n267), .B(G20), .C1(new_n271), .C2(new_n273), .ZN(new_n280));
  OAI21_X1  g0080(.A(G107), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  AOI22_X1  g0081(.A1(new_n262), .A2(G20), .B1(G77), .B2(new_n264), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT76), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n283), .A2(new_n284), .A3(new_n249), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n254), .B1(new_n278), .B2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT77), .ZN(new_n287));
  NAND2_X1  g0087(.A1(G33), .A2(G41), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n288), .A2(G1), .A3(G13), .ZN(new_n289));
  INV_X1    g0089(.A(G41), .ZN(new_n290));
  OAI211_X1 g0090(.A(new_n241), .B(G45), .C1(new_n290), .C2(KEYINPUT5), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT5), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n292), .A2(G41), .ZN(new_n293));
  OAI211_X1 g0093(.A(G257), .B(new_n289), .C1(new_n291), .C2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G45), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n296), .A2(G1), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n290), .A2(KEYINPUT5), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n292), .A2(G41), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n297), .A2(new_n298), .A3(new_n299), .A4(G274), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G1698), .ZN(new_n302));
  NAND4_X1  g0102(.A1(new_n271), .A2(new_n273), .A3(G244), .A4(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT4), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n268), .A2(KEYINPUT4), .A3(G244), .A4(new_n302), .ZN(new_n306));
  NAND2_X1  g0106(.A1(G33), .A2(G283), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n268), .A2(G250), .A3(G1698), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n305), .A2(new_n306), .A3(new_n307), .A4(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n289), .ZN(new_n310));
  AOI211_X1 g0110(.A(new_n295), .B(new_n301), .C1(new_n309), .C2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G200), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n287), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n309), .A2(new_n310), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n314), .A2(new_n300), .A3(new_n294), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n315), .A2(KEYINPUT77), .A3(G200), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n311), .A2(G190), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n286), .A2(new_n313), .A3(new_n316), .A4(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n268), .A2(new_n219), .A3(G68), .ZN(new_n319));
  NAND2_X1  g0119(.A1(G33), .A2(G97), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT19), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n219), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G87), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n323), .A2(new_n257), .A3(new_n255), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n219), .A2(G33), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n321), .B1(new_n326), .B2(new_n257), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n319), .A2(new_n325), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(new_n249), .ZN(new_n329));
  INV_X1    g0129(.A(new_n246), .ZN(new_n330));
  XNOR2_X1  g0130(.A(KEYINPUT15), .B(G87), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n246), .A2(new_n250), .A3(G87), .A4(new_n251), .ZN(new_n333));
  AND3_X1   g0133(.A1(new_n329), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n289), .B(G250), .C1(G1), .C2(new_n296), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n297), .A2(G274), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n268), .A2(G244), .A3(G1698), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n268), .A2(G238), .A3(new_n302), .ZN(new_n339));
  NAND2_X1  g0139(.A1(G33), .A2(G116), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n337), .B1(new_n341), .B2(new_n310), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(G190), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n334), .B(new_n343), .C1(new_n312), .C2(new_n342), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n341), .A2(new_n310), .ZN(new_n345));
  INV_X1    g0145(.A(new_n337), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(G169), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n246), .A2(new_n250), .A3(new_n251), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n329), .B(new_n332), .C1(new_n350), .C2(new_n331), .ZN(new_n351));
  INV_X1    g0151(.A(G179), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n342), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n349), .A2(new_n351), .A3(new_n353), .ZN(new_n354));
  AND2_X1   g0154(.A1(new_n344), .A2(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n284), .B1(new_n283), .B2(new_n249), .ZN(new_n356));
  AOI211_X1 g0156(.A(KEYINPUT76), .B(new_n250), .C1(new_n281), .C2(new_n282), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n253), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n311), .A2(new_n352), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n315), .A2(new_n348), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n358), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  AND3_X1   g0161(.A1(new_n318), .A2(new_n355), .A3(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(G1), .B1(new_n290), .B2(new_n296), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(G274), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n241), .B1(G41), .B2(G45), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n289), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(G226), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n364), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n274), .A2(new_n302), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n369), .A2(G223), .B1(G77), .B2(new_n274), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n268), .A2(KEYINPUT68), .A3(G222), .A4(new_n302), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT68), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n268), .A2(new_n302), .ZN(new_n373));
  INV_X1    g0173(.A(G222), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n372), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n370), .A2(new_n371), .A3(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n368), .B1(new_n376), .B2(new_n310), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n378), .A2(G179), .ZN(new_n379));
  INV_X1    g0179(.A(G50), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n330), .A2(new_n380), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n246), .B(new_n250), .C1(G1), .C2(new_n219), .ZN(new_n382));
  INV_X1    g0182(.A(G58), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n383), .A2(KEYINPUT8), .ZN(new_n384));
  XNOR2_X1  g0184(.A(KEYINPUT69), .B(G58), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n384), .B1(new_n385), .B2(KEYINPUT8), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n386), .A2(new_n326), .ZN(new_n387));
  OAI21_X1  g0187(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n388));
  INV_X1    g0188(.A(G150), .ZN(new_n389));
  INV_X1    g0189(.A(new_n264), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n388), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n387), .A2(new_n391), .ZN(new_n392));
  OAI221_X1 g0192(.A(new_n381), .B1(new_n380), .B2(new_n382), .C1(new_n392), .C2(new_n250), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n393), .B1(G169), .B2(new_n377), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n379), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(G190), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT9), .ZN(new_n397));
  OAI22_X1  g0197(.A1(new_n378), .A2(new_n396), .B1(new_n393), .B2(new_n397), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n392), .A2(new_n250), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n381), .B1(new_n382), .B2(new_n380), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  OAI22_X1  g0201(.A1(new_n401), .A2(KEYINPUT9), .B1(new_n312), .B2(new_n377), .ZN(new_n402));
  OAI21_X1  g0202(.A(KEYINPUT10), .B1(new_n398), .B2(new_n402), .ZN(new_n403));
  AOI22_X1  g0203(.A1(G200), .A2(new_n378), .B1(new_n393), .B2(new_n397), .ZN(new_n404));
  AOI22_X1  g0204(.A1(new_n401), .A2(KEYINPUT9), .B1(G190), .B2(new_n377), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT10), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n395), .B1(new_n403), .B2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT18), .ZN(new_n409));
  OAI21_X1  g0209(.A(G68), .B1(new_n279), .B2(new_n280), .ZN(new_n410));
  INV_X1    g0210(.A(G68), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n202), .B1(new_n385), .B2(new_n411), .ZN(new_n412));
  AOI22_X1  g0212(.A1(new_n412), .A2(G20), .B1(G159), .B2(new_n264), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT16), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n250), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n410), .A2(new_n413), .A3(KEYINPUT16), .ZN(new_n417));
  INV_X1    g0217(.A(new_n386), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n382), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n386), .A2(new_n246), .ZN(new_n420));
  AOI22_X1  g0220(.A1(new_n416), .A2(new_n417), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n271), .A2(new_n273), .A3(G226), .A4(G1698), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n271), .A2(new_n273), .A3(G223), .A4(new_n302), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n422), .B(new_n423), .C1(new_n270), .C2(new_n323), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n310), .ZN(new_n425));
  INV_X1    g0225(.A(G232), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n364), .B1(new_n366), .B2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n425), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(G169), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n425), .A2(G179), .A3(new_n428), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n409), .B1(new_n421), .B2(new_n433), .ZN(new_n434));
  AND2_X1   g0234(.A1(KEYINPUT69), .A2(G58), .ZN(new_n435));
  NOR2_X1   g0235(.A1(KEYINPUT69), .A2(G58), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n201), .B1(new_n437), .B2(G68), .ZN(new_n438));
  INV_X1    g0238(.A(G159), .ZN(new_n439));
  OAI22_X1  g0239(.A1(new_n438), .A2(new_n219), .B1(new_n439), .B2(new_n390), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n411), .B1(new_n269), .B2(new_n275), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n415), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n442), .A2(new_n417), .A3(new_n249), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n419), .B1(new_n330), .B2(new_n418), .ZN(new_n444));
  AOI22_X1  g0244(.A1(new_n443), .A2(new_n444), .B1(new_n430), .B2(new_n431), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(KEYINPUT18), .ZN(new_n446));
  OR2_X1    g0246(.A1(new_n396), .A2(KEYINPUT75), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n396), .A2(KEYINPUT75), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  AOI211_X1 g0249(.A(new_n449), .B(new_n427), .C1(new_n310), .C2(new_n424), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n312), .B1(new_n425), .B2(new_n428), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n452), .A2(new_n444), .A3(new_n443), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(KEYINPUT17), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT17), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n452), .A2(new_n443), .A3(new_n455), .A4(new_n444), .ZN(new_n456));
  AOI22_X1  g0256(.A1(new_n434), .A2(new_n446), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n274), .A2(G107), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n268), .A2(G1698), .ZN(new_n459));
  INV_X1    g0259(.A(G238), .ZN(new_n460));
  OAI221_X1 g0260(.A(new_n458), .B1(new_n459), .B2(new_n460), .C1(new_n426), .C2(new_n373), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(new_n310), .ZN(new_n462));
  INV_X1    g0262(.A(G244), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n364), .B1(new_n366), .B2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n348), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n464), .B1(new_n461), .B2(new_n310), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(new_n352), .ZN(new_n469));
  INV_X1    g0269(.A(G77), .ZN(new_n470));
  OR2_X1    g0270(.A1(new_n382), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n330), .A2(new_n470), .ZN(new_n472));
  NAND2_X1  g0272(.A1(G20), .A2(G77), .ZN(new_n473));
  XNOR2_X1  g0273(.A(KEYINPUT8), .B(G58), .ZN(new_n474));
  OAI221_X1 g0274(.A(new_n473), .B1(new_n331), .B2(new_n326), .C1(new_n390), .C2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(new_n249), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n471), .A2(new_n472), .A3(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n467), .A2(new_n469), .A3(new_n477), .ZN(new_n478));
  AND3_X1   g0278(.A1(new_n471), .A2(new_n472), .A3(new_n476), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n468), .A2(G190), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n479), .B(new_n480), .C1(new_n312), .C2(new_n468), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n408), .A2(new_n457), .A3(new_n478), .A4(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n330), .A2(new_n411), .ZN(new_n483));
  XNOR2_X1  g0283(.A(new_n483), .B(KEYINPUT12), .ZN(new_n484));
  OR2_X1    g0284(.A1(new_n382), .A2(new_n411), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n390), .A2(new_n380), .ZN(new_n486));
  OAI22_X1  g0286(.A1(new_n326), .A2(new_n470), .B1(new_n219), .B2(G68), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n249), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  XNOR2_X1  g0288(.A(new_n488), .B(KEYINPUT11), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n484), .A2(new_n485), .A3(new_n489), .ZN(new_n490));
  XNOR2_X1  g0290(.A(new_n490), .B(KEYINPUT74), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT13), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n268), .A2(G226), .A3(new_n302), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n493), .B(new_n320), .C1(new_n459), .C2(new_n426), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(new_n310), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n364), .B1(new_n366), .B2(new_n460), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n492), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  AOI211_X1 g0298(.A(KEYINPUT13), .B(new_n496), .C1(new_n494), .C2(new_n310), .ZN(new_n499));
  OAI21_X1  g0299(.A(G169), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g0300(.A1(KEYINPUT72), .A2(KEYINPUT14), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  OAI211_X1 g0303(.A(G169), .B(new_n501), .C1(new_n498), .C2(new_n499), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n495), .A2(new_n497), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n492), .A2(KEYINPUT71), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT73), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n495), .B(new_n497), .C1(KEYINPUT71), .C2(new_n492), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n507), .A2(new_n508), .A3(new_n509), .A4(G179), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n503), .A2(new_n504), .A3(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n507), .A2(G179), .A3(new_n509), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(KEYINPUT73), .ZN(new_n513));
  NAND2_X1  g0313(.A1(KEYINPUT72), .A2(KEYINPUT14), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n491), .B1(new_n511), .B2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(new_n490), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n507), .A2(G190), .A3(new_n509), .ZN(new_n518));
  OAI21_X1  g0318(.A(G200), .B1(new_n498), .B2(new_n499), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n516), .A2(new_n520), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n482), .A2(new_n521), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n243), .A2(KEYINPUT25), .A3(new_n255), .A4(new_n245), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT81), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT25), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n527), .B1(new_n246), .B2(G107), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n523), .A2(new_n524), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n526), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n252), .A2(G107), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT23), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n532), .B1(new_n219), .B2(G107), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n255), .A2(KEYINPUT23), .A3(G20), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n219), .A2(G33), .A3(G116), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n271), .A2(new_n273), .A3(new_n219), .A4(G87), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(KEYINPUT22), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT22), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n268), .A2(new_n540), .A3(new_n219), .A4(G87), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n537), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(KEYINPUT24), .ZN(new_n543));
  INV_X1    g0343(.A(new_n543), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n249), .B1(new_n542), .B2(KEYINPUT24), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n530), .B(new_n531), .C1(new_n544), .C2(new_n545), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n271), .A2(new_n273), .A3(G250), .A4(new_n302), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n271), .A2(new_n273), .A3(G257), .A4(G1698), .ZN(new_n548));
  INV_X1    g0348(.A(G294), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n547), .B(new_n548), .C1(new_n270), .C2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n310), .ZN(new_n551));
  OAI211_X1 g0351(.A(G264), .B(new_n289), .C1(new_n291), .C2(new_n293), .ZN(new_n552));
  AND2_X1   g0352(.A1(new_n552), .A2(new_n300), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT82), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n552), .A2(new_n300), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n557), .B1(new_n310), .B2(new_n550), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(KEYINPUT82), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n556), .A2(new_n559), .A3(new_n396), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n554), .A2(new_n312), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n546), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n348), .B1(new_n556), .B2(new_n559), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n551), .A2(G179), .A3(new_n553), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT83), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n558), .A2(KEYINPUT83), .A3(G179), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n546), .B1(new_n563), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(KEYINPUT84), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT84), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n546), .B(new_n571), .C1(new_n563), .C2(new_n568), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n562), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT21), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n271), .A2(new_n273), .A3(G264), .A4(G1698), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT79), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n268), .A2(KEYINPUT79), .A3(G264), .A4(G1698), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n274), .A2(G303), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n268), .A2(G257), .A3(new_n302), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n577), .A2(new_n578), .A3(new_n579), .A4(new_n580), .ZN(new_n581));
  AND2_X1   g0381(.A1(new_n581), .A2(new_n310), .ZN(new_n582));
  OAI211_X1 g0382(.A(G270), .B(new_n289), .C1(new_n291), .C2(new_n293), .ZN(new_n583));
  AND3_X1   g0383(.A1(new_n583), .A2(KEYINPUT78), .A3(new_n300), .ZN(new_n584));
  AOI21_X1  g0384(.A(KEYINPUT78), .B1(new_n583), .B2(new_n300), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  OAI21_X1  g0386(.A(G169), .B1(new_n582), .B2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(G116), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n330), .A2(new_n588), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n589), .B1(new_n350), .B2(new_n588), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n248), .A2(new_n218), .B1(G20), .B2(new_n588), .ZN(new_n591));
  AOI21_X1  g0391(.A(G20), .B1(G33), .B2(G283), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n270), .A2(G97), .ZN(new_n593));
  AND3_X1   g0393(.A1(new_n592), .A2(new_n593), .A3(KEYINPUT80), .ZN(new_n594));
  AOI21_X1  g0394(.A(KEYINPUT80), .B1(new_n592), .B2(new_n593), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n591), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT20), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  OAI211_X1 g0398(.A(KEYINPUT20), .B(new_n591), .C1(new_n594), .C2(new_n595), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n590), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n574), .B1(new_n587), .B2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(new_n585), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n583), .A2(KEYINPUT78), .A3(new_n300), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n581), .A2(new_n310), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(G200), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n607), .B(new_n600), .C1(new_n606), .C2(new_n449), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n598), .A2(new_n599), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n609), .B(new_n589), .C1(new_n588), .C2(new_n350), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n610), .A2(new_n606), .A3(KEYINPUT21), .A4(G169), .ZN(new_n611));
  NOR3_X1   g0411(.A1(new_n582), .A2(new_n586), .A3(new_n352), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n610), .ZN(new_n613));
  AND4_X1   g0413(.A1(new_n601), .A2(new_n608), .A3(new_n611), .A4(new_n613), .ZN(new_n614));
  AND4_X1   g0414(.A1(new_n362), .A2(new_n522), .A3(new_n573), .A4(new_n614), .ZN(G372));
  INV_X1    g0415(.A(new_n395), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n434), .A2(new_n446), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n520), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n516), .B1(new_n619), .B2(new_n478), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n454), .A2(new_n456), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n618), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n403), .A2(new_n407), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n616), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n601), .A2(new_n611), .A3(new_n613), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n569), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n560), .A2(new_n561), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n528), .A2(new_n529), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n531), .B1(new_n629), .B2(new_n525), .ZN(new_n630));
  INV_X1    g0430(.A(new_n545), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n630), .B1(new_n631), .B2(new_n543), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n628), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n362), .A2(new_n627), .A3(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n354), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n315), .A2(G179), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n311), .A2(G169), .ZN(new_n637));
  NOR3_X1   g0437(.A1(new_n286), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n638), .A2(KEYINPUT26), .A3(new_n355), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT26), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n344), .A2(new_n354), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n640), .B1(new_n361), .B2(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n635), .B1(new_n639), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n634), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n625), .B1(new_n522), .B2(new_n644), .ZN(new_n645));
  XNOR2_X1  g0445(.A(new_n645), .B(KEYINPUT85), .ZN(G369));
  INV_X1    g0446(.A(G330), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n241), .A2(new_n219), .A3(G13), .ZN(new_n648));
  OR2_X1    g0448(.A1(new_n648), .A2(KEYINPUT27), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT86), .ZN(new_n650));
  OR2_X1    g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n649), .A2(new_n650), .ZN(new_n652));
  INV_X1    g0452(.A(G213), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n653), .B1(new_n648), .B2(KEYINPUT27), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n651), .A2(new_n652), .A3(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(G343), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n614), .B1(new_n600), .B2(new_n658), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n601), .A2(new_n613), .A3(new_n611), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n660), .A2(new_n610), .A3(new_n657), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(KEYINPUT87), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT87), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n659), .A2(new_n664), .A3(new_n661), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n647), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n570), .A2(new_n572), .ZN(new_n667));
  OAI211_X1 g0467(.A(new_n667), .B(new_n633), .C1(new_n632), .C2(new_n658), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n556), .A2(new_n559), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(G169), .ZN(new_n670));
  AND2_X1   g0470(.A1(new_n566), .A2(new_n567), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n632), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n657), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n668), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n666), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n626), .A2(new_n657), .ZN(new_n676));
  AOI22_X1  g0476(.A1(new_n573), .A2(new_n676), .B1(new_n672), .B2(new_n658), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n675), .A2(new_n677), .ZN(G399));
  NOR2_X1   g0478(.A1(new_n324), .A2(G116), .ZN(new_n679));
  XOR2_X1   g0479(.A(new_n679), .B(KEYINPUT88), .Z(new_n680));
  INV_X1    g0480(.A(new_n206), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n681), .A2(G41), .ZN(new_n682));
  NOR3_X1   g0482(.A1(new_n680), .A2(new_n241), .A3(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n221), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n683), .B1(new_n684), .B2(new_n682), .ZN(new_n685));
  XNOR2_X1  g0485(.A(KEYINPUT89), .B(KEYINPUT28), .ZN(new_n686));
  XNOR2_X1  g0486(.A(new_n685), .B(new_n686), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n573), .A2(new_n362), .A3(new_n614), .A4(new_n658), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n604), .A2(G179), .A3(new_n605), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n558), .A2(new_n342), .A3(new_n314), .A4(new_n294), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT30), .ZN(new_n691));
  NOR3_X1   g0491(.A1(new_n689), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n691), .B1(new_n689), .B2(new_n690), .ZN(new_n693));
  NOR3_X1   g0493(.A1(new_n558), .A2(new_n342), .A3(G179), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n694), .A2(new_n315), .A3(new_n606), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n692), .B1(new_n696), .B2(KEYINPUT90), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT90), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n693), .A2(new_n695), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT31), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n658), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(KEYINPUT91), .B1(new_n688), .B2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n702), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n705), .B1(new_n697), .B2(new_n699), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT91), .ZN(new_n707));
  AND4_X1   g0507(.A1(new_n342), .A2(new_n558), .A3(new_n314), .A4(new_n294), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n612), .A2(new_n708), .A3(KEYINPUT30), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n709), .A2(new_n693), .A3(new_n695), .ZN(new_n710));
  AND2_X1   g0510(.A1(new_n710), .A2(new_n657), .ZN(new_n711));
  OAI22_X1  g0511(.A1(new_n706), .A2(new_n707), .B1(KEYINPUT31), .B2(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(G330), .B1(new_n704), .B2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n318), .A2(new_n633), .A3(new_n361), .A4(new_n355), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n715), .B1(new_n667), .B2(new_n626), .ZN(new_n716));
  AOI21_X1  g0516(.A(KEYINPUT26), .B1(new_n638), .B2(new_n355), .ZN(new_n717));
  NOR3_X1   g0517(.A1(new_n361), .A2(new_n640), .A3(new_n641), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n354), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n658), .B1(new_n716), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(KEYINPUT29), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n657), .B1(new_n634), .B2(new_n643), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT29), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n721), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n714), .A2(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n687), .B1(new_n726), .B2(G1), .ZN(G364));
  INV_X1    g0527(.A(G13), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(G20), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n241), .B1(new_n729), .B2(G45), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n682), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n666), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n663), .A2(new_n665), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n733), .B1(G330), .B2(new_n734), .ZN(new_n735));
  AND2_X1   g0535(.A1(new_n735), .A2(KEYINPUT92), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n735), .A2(KEYINPUT92), .ZN(new_n737));
  XNOR2_X1  g0537(.A(new_n732), .B(KEYINPUT93), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n681), .A2(new_n274), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(G355), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n741), .B1(G116), .B2(new_n206), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n222), .A2(new_n296), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n681), .A2(new_n268), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n745), .B1(new_n239), .B2(G45), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n742), .B1(new_n743), .B2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(G13), .A2(G33), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(G20), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n218), .B1(G20), .B2(new_n348), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n739), .B1(new_n747), .B2(new_n753), .ZN(new_n754));
  NOR3_X1   g0554(.A1(new_n219), .A2(new_n312), .A3(G179), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(G190), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(new_n323), .ZN(new_n757));
  NAND2_X1  g0557(.A1(G20), .A2(G179), .ZN(new_n758));
  NOR3_X1   g0558(.A1(new_n758), .A2(new_n312), .A3(G190), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR3_X1   g0560(.A1(new_n449), .A2(new_n312), .A3(new_n758), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  OAI221_X1 g0562(.A(new_n268), .B1(new_n411), .B2(new_n760), .C1(new_n762), .C2(new_n380), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G179), .A2(G200), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n764), .A2(G20), .A3(new_n396), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(G159), .ZN(new_n767));
  AOI211_X1 g0567(.A(new_n757), .B(new_n763), .C1(KEYINPUT32), .C2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n449), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n758), .A2(G200), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n219), .B1(new_n764), .B2(G190), .ZN(new_n772));
  OAI22_X1  g0572(.A1(new_n771), .A2(new_n385), .B1(new_n257), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n755), .A2(new_n396), .ZN(new_n774));
  OAI22_X1  g0574(.A1(new_n767), .A2(KEYINPUT32), .B1(new_n774), .B2(new_n255), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  AND3_X1   g0576(.A1(new_n770), .A2(KEYINPUT94), .A3(new_n396), .ZN(new_n777));
  AOI21_X1  g0577(.A(KEYINPUT94), .B1(new_n770), .B2(new_n396), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  OAI211_X1 g0579(.A(new_n768), .B(new_n776), .C1(new_n470), .C2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(G311), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(G322), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n771), .A2(new_n783), .B1(new_n549), .B2(new_n772), .ZN(new_n784));
  INV_X1    g0584(.A(new_n774), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n784), .B1(G283), .B2(new_n785), .ZN(new_n786));
  XOR2_X1   g0586(.A(KEYINPUT33), .B(G317), .Z(new_n787));
  NOR2_X1   g0587(.A1(new_n760), .A2(new_n787), .ZN(new_n788));
  AOI211_X1 g0588(.A(new_n268), .B(new_n788), .C1(G329), .C2(new_n766), .ZN(new_n789));
  INV_X1    g0589(.A(new_n756), .ZN(new_n790));
  AOI22_X1  g0590(.A1(new_n761), .A2(G326), .B1(G303), .B2(new_n790), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n786), .A2(new_n789), .A3(new_n791), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n780), .B1(new_n782), .B2(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n754), .B1(new_n793), .B2(new_n751), .ZN(new_n794));
  INV_X1    g0594(.A(new_n750), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n794), .B1(new_n734), .B2(new_n795), .ZN(new_n796));
  XNOR2_X1  g0596(.A(new_n796), .B(KEYINPUT95), .ZN(new_n797));
  NOR3_X1   g0597(.A1(new_n736), .A2(new_n737), .A3(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(G396));
  NAND2_X1  g0599(.A1(new_n477), .A2(new_n657), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n481), .A2(new_n478), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(KEYINPUT100), .ZN(new_n802));
  INV_X1    g0602(.A(KEYINPUT100), .ZN(new_n803));
  NAND4_X1  g0603(.A1(new_n481), .A2(new_n478), .A3(new_n803), .A4(new_n800), .ZN(new_n804));
  AND2_X1   g0604(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n660), .A2(new_n672), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n715), .A2(new_n806), .ZN(new_n807));
  OAI211_X1 g0607(.A(new_n658), .B(new_n805), .C1(new_n719), .C2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(KEYINPUT101), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND4_X1  g0610(.A1(new_n644), .A2(KEYINPUT101), .A3(new_n658), .A4(new_n805), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n478), .A2(new_n658), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n813), .B1(new_n802), .B2(new_n804), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  OR2_X1    g0615(.A1(new_n722), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n812), .A2(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n732), .B1(new_n817), .B2(new_n713), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n818), .B1(new_n713), .B2(new_n817), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT102), .ZN(new_n820));
  INV_X1    g0620(.A(new_n751), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n821), .A2(new_n749), .ZN(new_n822));
  AOI22_X1  g0622(.A1(new_n761), .A2(G137), .B1(G150), .B2(new_n759), .ZN(new_n823));
  INV_X1    g0623(.A(G143), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n823), .B1(new_n824), .B2(new_n771), .ZN(new_n825));
  INV_X1    g0625(.A(new_n779), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n825), .B1(G159), .B2(new_n826), .ZN(new_n827));
  XNOR2_X1  g0627(.A(KEYINPUT98), .B(KEYINPUT34), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  AND2_X1   g0629(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n827), .A2(new_n829), .ZN(new_n831));
  INV_X1    g0631(.A(G132), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n268), .B1(new_n832), .B2(new_n765), .C1(new_n774), .C2(new_n411), .ZN(new_n833));
  OAI22_X1  g0633(.A1(new_n756), .A2(new_n380), .B1(new_n385), .B2(new_n772), .ZN(new_n834));
  NOR4_X1   g0634(.A1(new_n830), .A2(new_n831), .A3(new_n833), .A4(new_n834), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n826), .A2(G116), .B1(G283), .B2(new_n759), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT96), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n836), .A2(new_n837), .B1(G303), .B2(new_n761), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n838), .B1(new_n837), .B2(new_n836), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n839), .B(KEYINPUT97), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n274), .B1(new_n765), .B2(new_n781), .C1(new_n257), .C2(new_n772), .ZN(new_n841));
  OAI22_X1  g0641(.A1(new_n774), .A2(new_n323), .B1(new_n756), .B2(new_n255), .ZN(new_n842));
  INV_X1    g0642(.A(new_n771), .ZN(new_n843));
  AOI211_X1 g0643(.A(new_n841), .B(new_n842), .C1(G294), .C2(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n835), .B1(new_n840), .B2(new_n844), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n739), .B1(G77), .B2(new_n822), .C1(new_n845), .C2(new_n821), .ZN(new_n846));
  OR2_X1    g0646(.A1(new_n846), .A2(KEYINPUT99), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(KEYINPUT99), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n847), .B(new_n848), .C1(new_n749), .C2(new_n815), .ZN(new_n849));
  AND3_X1   g0649(.A1(new_n819), .A2(new_n820), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n820), .B1(new_n819), .B2(new_n849), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(G384));
  OR2_X1    g0653(.A1(new_n262), .A2(KEYINPUT35), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n854), .A2(G116), .A3(new_n220), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n855), .B1(KEYINPUT35), .B2(new_n262), .ZN(new_n856));
  OR2_X1    g0656(.A1(new_n856), .A2(KEYINPUT36), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(KEYINPUT36), .ZN(new_n858));
  AOI211_X1 g0658(.A(new_n470), .B(new_n221), .C1(new_n437), .C2(G68), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n411), .A2(G50), .ZN(new_n860));
  OAI211_X1 g0660(.A(G1), .B(new_n728), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n857), .A2(new_n858), .A3(new_n861), .ZN(new_n862));
  XOR2_X1   g0662(.A(new_n862), .B(KEYINPUT103), .Z(new_n863));
  INV_X1    g0663(.A(KEYINPUT37), .ZN(new_n864));
  NOR2_X1   g0664(.A1(KEYINPUT104), .A2(KEYINPUT16), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n865), .B1(new_n440), .B2(new_n441), .ZN(new_n866));
  INV_X1    g0666(.A(new_n865), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n410), .A2(new_n413), .A3(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n866), .A2(new_n868), .A3(new_n249), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(new_n444), .ZN(new_n870));
  INV_X1    g0670(.A(new_n655), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n421), .A2(new_n452), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n870), .A2(new_n432), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n864), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n443), .A2(new_n444), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n432), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n871), .ZN(new_n877));
  AND4_X1   g0677(.A1(new_n864), .A2(new_n876), .A3(new_n877), .A4(new_n453), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n874), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n870), .A2(new_n871), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n880), .B1(new_n617), .B2(new_n621), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT38), .ZN(new_n882));
  NOR3_X1   g0682(.A1(new_n879), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n617), .A2(new_n621), .ZN(new_n884));
  INV_X1    g0684(.A(new_n877), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n876), .A2(new_n877), .A3(new_n453), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(KEYINPUT37), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n876), .A2(new_n877), .A3(new_n864), .A4(new_n453), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(KEYINPUT38), .B1(new_n886), .B2(new_n890), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n883), .A2(new_n891), .ZN(new_n892));
  OR2_X1    g0692(.A1(KEYINPUT107), .A2(KEYINPUT31), .ZN(new_n893));
  AND3_X1   g0693(.A1(new_n710), .A2(new_n657), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n893), .B1(new_n710), .B2(new_n657), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n688), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n491), .A2(new_n657), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n516), .A2(new_n520), .A3(new_n898), .ZN(new_n899));
  AOI22_X1  g0699(.A1(new_n512), .A2(KEYINPUT73), .B1(KEYINPUT72), .B2(KEYINPUT14), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n900), .A2(new_n504), .A3(new_n510), .A4(new_n503), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n491), .B(new_n657), .C1(new_n901), .C2(new_n619), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n897), .A2(new_n903), .A3(new_n815), .ZN(new_n904));
  OAI21_X1  g0704(.A(KEYINPUT40), .B1(new_n892), .B2(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n882), .B1(new_n879), .B2(new_n881), .ZN(new_n906));
  AND3_X1   g0706(.A1(new_n880), .A2(new_n873), .A3(new_n453), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n889), .B1(new_n907), .B2(new_n864), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n908), .B(KEYINPUT38), .C1(new_n457), .C2(new_n880), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n906), .A2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT40), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n814), .B1(new_n688), .B2(new_n896), .ZN(new_n912));
  NAND4_X1  g0712(.A1(new_n910), .A2(new_n911), .A3(new_n912), .A4(new_n903), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n905), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(G330), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n522), .A2(G330), .A3(new_n897), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n914), .A2(new_n522), .A3(new_n897), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n725), .A2(new_n522), .ZN(new_n920));
  INV_X1    g0720(.A(new_n625), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  XOR2_X1   g0722(.A(new_n919), .B(new_n922), .Z(new_n923));
  INV_X1    g0723(.A(KEYINPUT105), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n445), .B1(new_n421), .B2(new_n452), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n864), .B1(new_n925), .B2(new_n877), .ZN(new_n926));
  OAI22_X1  g0726(.A1(new_n926), .A2(new_n878), .B1(new_n457), .B2(new_n877), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n924), .B1(new_n927), .B2(new_n882), .ZN(new_n928));
  OAI21_X1  g0728(.A(KEYINPUT39), .B1(new_n910), .B2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n891), .ZN(new_n930));
  NOR2_X1   g0730(.A1(KEYINPUT105), .A2(KEYINPUT39), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n930), .A2(new_n909), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n929), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(KEYINPUT106), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n901), .A2(new_n491), .A3(new_n658), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT106), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n929), .A2(new_n937), .A3(new_n932), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n934), .A2(new_n936), .A3(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n478), .A2(new_n657), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n940), .B1(new_n810), .B2(new_n811), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n942), .A2(new_n910), .A3(new_n903), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n618), .A2(new_n655), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n939), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n923), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n241), .B2(new_n729), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n923), .A2(new_n946), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n863), .B1(new_n948), .B2(new_n949), .ZN(G367));
  OAI211_X1 g0750(.A(new_n318), .B(new_n361), .C1(new_n286), .C2(new_n658), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n638), .A2(new_n657), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n573), .A2(new_n676), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n957), .A2(KEYINPUT42), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n361), .B1(new_n951), .B2(new_n667), .ZN(new_n959));
  AOI22_X1  g0759(.A1(new_n957), .A2(KEYINPUT42), .B1(new_n658), .B2(new_n959), .ZN(new_n960));
  OR2_X1    g0760(.A1(new_n658), .A2(new_n334), .ZN(new_n961));
  OR2_X1    g0761(.A1(new_n961), .A2(new_n354), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n355), .A2(new_n961), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  AOI22_X1  g0764(.A1(new_n958), .A2(new_n960), .B1(KEYINPUT43), .B2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n964), .A2(KEYINPUT43), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT108), .ZN(new_n968));
  OAI21_X1  g0768(.A(KEYINPUT109), .B1(new_n675), .B2(new_n954), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT109), .ZN(new_n970));
  NAND4_X1  g0770(.A1(new_n666), .A2(new_n970), .A3(new_n674), .A4(new_n953), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n968), .B1(new_n969), .B2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(new_n972), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n969), .A2(new_n971), .A3(new_n968), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n967), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n974), .ZN(new_n976));
  INV_X1    g0776(.A(new_n967), .ZN(new_n977));
  NOR3_X1   g0777(.A1(new_n976), .A2(new_n977), .A3(new_n972), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n966), .B1(new_n975), .B2(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n977), .B1(new_n976), .B2(new_n972), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n973), .A2(new_n967), .A3(new_n974), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n980), .A2(new_n981), .A3(new_n965), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n979), .A2(new_n982), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n682), .B(KEYINPUT41), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n955), .B1(new_n674), .B2(new_n676), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n666), .B(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(new_n726), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n677), .A2(new_n953), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n988), .B(KEYINPUT45), .Z(new_n989));
  NOR2_X1   g0789(.A1(new_n677), .A2(new_n953), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT44), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n989), .A2(new_n675), .A3(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n675), .B1(new_n989), .B2(new_n991), .ZN(new_n994));
  NOR3_X1   g0794(.A1(new_n987), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(new_n726), .ZN(new_n996));
  OAI211_X1 g0796(.A(KEYINPUT110), .B(new_n984), .C1(new_n995), .C2(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n984), .B1(new_n995), .B2(new_n996), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT110), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n731), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n983), .B1(new_n997), .B2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n227), .A2(new_n745), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n752), .B1(new_n206), .B2(new_n331), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n739), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(G317), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n274), .B1(new_n765), .B2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(KEYINPUT46), .B1(new_n790), .B2(G116), .ZN(new_n1007));
  AOI211_X1 g0807(.A(new_n1006), .B(new_n1007), .C1(G294), .C2(new_n759), .ZN(new_n1008));
  INV_X1    g0808(.A(G303), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n762), .A2(new_n781), .B1(new_n1009), .B2(new_n771), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n774), .A2(new_n257), .B1(new_n255), .B2(new_n772), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n790), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n826), .A2(G283), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n1008), .A2(new_n1012), .A3(new_n1013), .A4(new_n1014), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n779), .A2(new_n380), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n772), .A2(new_n411), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n774), .A2(new_n470), .ZN(new_n1018));
  AOI211_X1 g0818(.A(new_n1017), .B(new_n1018), .C1(G143), .C2(new_n761), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n268), .B1(new_n760), .B2(new_n439), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1020), .B1(G137), .B2(new_n766), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n843), .A2(G150), .B1(new_n437), .B2(new_n790), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1019), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1015), .B1(new_n1016), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT47), .ZN(new_n1025));
  OR2_X1    g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n821), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1004), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n962), .A2(new_n963), .A3(new_n750), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n1030), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n1001), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n1032), .ZN(G387));
  NAND2_X1  g0833(.A1(new_n986), .A2(new_n731), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n745), .B1(new_n232), .B2(G45), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1035), .B1(new_n680), .B2(new_n740), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n474), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(new_n380), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n296), .B1(new_n411), .B2(new_n470), .C1(new_n1038), .C2(KEYINPUT50), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n680), .B(new_n1039), .C1(KEYINPUT50), .C2(new_n1038), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n1036), .A2(new_n1040), .B1(G107), .B2(new_n206), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n738), .B1(new_n1041), .B2(new_n752), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n772), .A2(new_n331), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(new_n843), .B2(G50), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1044), .B1(new_n470), .B2(new_n756), .C1(new_n439), .C2(new_n762), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n779), .A2(new_n411), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n386), .A2(new_n760), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n268), .B1(new_n389), .B2(new_n765), .C1(new_n774), .C2(new_n257), .ZN(new_n1048));
  NOR4_X1   g0848(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n761), .A2(G322), .B1(G311), .B2(new_n759), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1050), .B1(new_n1005), .B2(new_n771), .C1(new_n779), .C2(new_n1009), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT48), .ZN(new_n1052));
  INV_X1    g0852(.A(G283), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n1052), .B1(new_n1053), .B2(new_n772), .C1(new_n549), .C2(new_n756), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT49), .ZN(new_n1055));
  OR2_X1    g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n268), .B1(new_n766), .B2(G326), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n588), .B2(new_n774), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1049), .B1(new_n1056), .B2(new_n1059), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n1042), .B1(new_n674), .B2(new_n795), .C1(new_n1060), .C2(new_n821), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n987), .A2(new_n682), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n986), .A2(new_n726), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n1034), .B(new_n1061), .C1(new_n1062), .C2(new_n1063), .ZN(G393));
  OAI21_X1  g0864(.A(new_n994), .B1(new_n993), .B2(KEYINPUT111), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n994), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT111), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1066), .A2(new_n1067), .A3(new_n992), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1065), .A2(new_n1068), .A3(new_n987), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT113), .ZN(new_n1070));
  NOR3_X1   g0870(.A1(new_n995), .A2(G41), .A3(new_n681), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1065), .A2(new_n1068), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1073), .A2(new_n731), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n236), .A2(new_n745), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n752), .B1(new_n257), .B2(new_n206), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n739), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n762), .A2(new_n389), .B1(new_n439), .B2(new_n771), .ZN(new_n1078));
  INV_X1    g0878(.A(KEYINPUT51), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n1078), .A2(new_n1079), .B1(new_n1037), .B2(new_n826), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n774), .A2(new_n323), .B1(new_n756), .B2(new_n411), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n268), .B1(new_n765), .B2(new_n824), .C1(new_n760), .C2(new_n380), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n772), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n1081), .B(new_n1082), .C1(G77), .C2(new_n1083), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n1080), .B(new_n1084), .C1(new_n1079), .C2(new_n1078), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n843), .A2(G311), .B1(G317), .B2(new_n761), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1086), .B(KEYINPUT52), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n774), .A2(new_n255), .B1(new_n756), .B2(new_n1053), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n274), .B1(new_n765), .B2(new_n783), .C1(new_n760), .C2(new_n1009), .ZN(new_n1089));
  AOI211_X1 g0889(.A(new_n1088), .B(new_n1089), .C1(G116), .C2(new_n1083), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(new_n549), .B2(new_n779), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1085), .B1(new_n1087), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT112), .ZN(new_n1093));
  OR2_X1    g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n821), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1077), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1096), .B1(new_n953), .B2(new_n795), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1074), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1072), .A2(new_n1099), .ZN(G390));
  INV_X1    g0900(.A(new_n903), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n935), .B1(new_n941), .B2(new_n1101), .ZN(new_n1102));
  AND3_X1   g0902(.A1(new_n929), .A2(new_n937), .A3(new_n932), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n937), .B1(new_n929), .B2(new_n932), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1102), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  OAI211_X1 g0905(.A(G330), .B(new_n815), .C1(new_n704), .C2(new_n712), .ZN(new_n1106));
  OR2_X1    g0906(.A1(new_n1106), .A2(new_n1101), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n802), .A2(new_n804), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n720), .A2(new_n1108), .B1(new_n478), .B2(new_n657), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n936), .B(new_n892), .C1(new_n1109), .C2(new_n903), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1105), .A2(new_n1107), .A3(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n934), .A2(new_n938), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1110), .B1(new_n1113), .B2(new_n1102), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n912), .A2(G330), .A3(new_n903), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1112), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n920), .A2(new_n921), .A3(new_n916), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n720), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n940), .B1(new_n1119), .B2(new_n805), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n903), .B1(new_n912), .B2(G330), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1120), .B1(new_n1121), .B2(KEYINPUT114), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n897), .A2(G330), .A3(new_n815), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n1101), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n1106), .B2(new_n1101), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1122), .B1(new_n1125), .B2(KEYINPUT114), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1106), .A2(new_n1101), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n941), .B1(new_n1127), .B2(new_n1115), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1118), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1116), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1125), .A2(KEYINPUT114), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT114), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1109), .B1(new_n1124), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1128), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1117), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n1136), .B(new_n1112), .C1(new_n1114), .C2(new_n1115), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1130), .A2(new_n1137), .A3(new_n682), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n1112), .B(new_n731), .C1(new_n1114), .C2(new_n1115), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT116), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n749), .B1(new_n934), .B2(new_n938), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n774), .A2(new_n411), .B1(new_n756), .B2(new_n323), .ZN(new_n1142));
  OAI221_X1 g0942(.A(new_n274), .B1(new_n765), .B2(new_n549), .C1(new_n760), .C2(new_n255), .ZN(new_n1143));
  AOI211_X1 g0943(.A(new_n1142), .B(new_n1143), .C1(G283), .C2(new_n761), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n771), .A2(new_n588), .B1(new_n470), .B2(new_n772), .ZN(new_n1145));
  OR2_X1    g0945(.A1(new_n1145), .A2(KEYINPUT115), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1145), .A2(KEYINPUT115), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n826), .A2(G97), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n1144), .A2(new_n1146), .A3(new_n1147), .A4(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(G128), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n762), .A2(new_n1150), .B1(new_n380), .B2(new_n774), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n771), .A2(new_n832), .B1(new_n439), .B2(new_n772), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n790), .A2(G150), .ZN(new_n1154));
  OR2_X1    g0954(.A1(new_n1154), .A2(KEYINPUT53), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n274), .B1(G137), .B2(new_n759), .ZN(new_n1156));
  INV_X1    g0956(.A(G125), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1156), .B1(new_n1157), .B2(new_n765), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1158), .B1(KEYINPUT53), .B2(new_n1154), .ZN(new_n1159));
  XOR2_X1   g0959(.A(KEYINPUT54), .B(G143), .Z(new_n1160));
  NAND2_X1  g0960(.A1(new_n826), .A2(new_n1160), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n1153), .A2(new_n1155), .A3(new_n1159), .A4(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n821), .B1(new_n1149), .B2(new_n1162), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n739), .B1(new_n418), .B2(new_n822), .ZN(new_n1164));
  OR3_X1    g0964(.A1(new_n1141), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  AND3_X1   g0965(.A1(new_n1139), .A2(new_n1140), .A3(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1140), .B1(new_n1139), .B2(new_n1165), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1138), .B1(new_n1166), .B2(new_n1167), .ZN(G378));
  NAND2_X1  g0968(.A1(new_n1137), .A2(new_n1118), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT57), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n623), .A2(new_n616), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n401), .A2(new_n655), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1172), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n408), .A2(new_n1174), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1173), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1176), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n408), .A2(new_n1174), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n395), .B(new_n1172), .C1(new_n403), .C2(new_n407), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1178), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  AND2_X1   g0981(.A1(new_n1177), .A2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(new_n914), .B2(G330), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n647), .B(new_n1182), .C1(new_n905), .C2(new_n913), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  NAND4_X1  g0986(.A1(new_n1186), .A2(new_n943), .A3(new_n944), .A4(new_n939), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n915), .A2(new_n1182), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n914), .A2(G330), .A3(new_n1183), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1190), .A2(new_n945), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1170), .B1(new_n1187), .B2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1169), .A2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1193), .A2(new_n682), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n946), .B1(KEYINPUT118), .B2(new_n1186), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT118), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1190), .A2(new_n945), .A3(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1195), .A2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(KEYINPUT57), .B1(new_n1198), .B2(new_n1169), .ZN(new_n1199));
  OR2_X1    g0999(.A1(new_n1194), .A2(new_n1199), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n732), .B1(new_n822), .B2(G50), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1183), .A2(new_n749), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n380), .B1(G33), .B2(G41), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(new_n274), .B2(new_n290), .ZN(new_n1204));
  AOI211_X1 g1004(.A(G41), .B(new_n268), .C1(new_n766), .C2(G283), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1205), .B1(new_n257), .B2(new_n760), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n1017), .B(new_n1206), .C1(G77), .C2(new_n790), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n762), .A2(new_n588), .B1(new_n255), .B2(new_n771), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n774), .A2(new_n385), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  OAI211_X1 g1010(.A(new_n1207), .B(new_n1210), .C1(new_n331), .C2(new_n779), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT58), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1204), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n762), .A2(new_n1157), .B1(new_n832), .B2(new_n760), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n843), .A2(G128), .B1(G150), .B2(new_n1083), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1160), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1215), .B1(new_n756), .B2(new_n1216), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n1214), .B(new_n1217), .C1(G137), .C2(new_n826), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(KEYINPUT117), .B(KEYINPUT59), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  AOI211_X1 g1020(.A(G33), .B(G41), .C1(new_n766), .C2(G124), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1220), .B(new_n1221), .C1(new_n439), .C2(new_n774), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1223));
  OAI221_X1 g1023(.A(new_n1213), .B1(new_n1212), .B2(new_n1211), .C1(new_n1222), .C2(new_n1223), .ZN(new_n1224));
  AOI211_X1 g1024(.A(new_n1201), .B(new_n1202), .C1(new_n751), .C2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(new_n1198), .B2(new_n731), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1200), .A2(new_n1226), .ZN(G375));
  AOI21_X1  g1027(.A(new_n730), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1101), .A2(new_n748), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n739), .B1(G68), .B2(new_n822), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n771), .A2(new_n1053), .B1(new_n257), .B2(new_n756), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(G294), .B2(new_n761), .ZN(new_n1232));
  OAI221_X1 g1032(.A(new_n274), .B1(new_n765), .B2(new_n1009), .C1(new_n760), .C2(new_n588), .ZN(new_n1233));
  NOR3_X1   g1033(.A1(new_n1233), .A2(new_n1018), .A3(new_n1043), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n1232), .B(new_n1234), .C1(new_n255), .C2(new_n779), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n779), .A2(new_n389), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n756), .A2(new_n439), .B1(new_n380), .B2(new_n772), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(new_n843), .B2(G137), .ZN(new_n1238));
  OAI221_X1 g1038(.A(new_n268), .B1(new_n1150), .B2(new_n765), .C1(new_n1216), .C2(new_n760), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1209), .B1(new_n761), .B2(G132), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1238), .A2(new_n1240), .A3(new_n1241), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1235), .B1(new_n1236), .B2(new_n1242), .ZN(new_n1243));
  OR2_X1    g1043(.A1(new_n1243), .A2(KEYINPUT119), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n821), .B1(new_n1243), .B2(KEYINPUT119), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1230), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1228), .B1(new_n1229), .B2(new_n1246), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1134), .A2(new_n1117), .A3(new_n1135), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1129), .A2(new_n984), .A3(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1247), .A2(new_n1249), .ZN(G381));
  AND2_X1   g1050(.A1(new_n1139), .A2(new_n1165), .ZN(new_n1251));
  AND2_X1   g1051(.A1(new_n1138), .A2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(G375), .A2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(G381), .ZN(new_n1255));
  NOR4_X1   g1055(.A1(G390), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1254), .A2(new_n1032), .A3(new_n1255), .A4(new_n1256), .ZN(G407));
  NOR2_X1   g1057(.A1(new_n653), .A2(G343), .ZN(new_n1258));
  XNOR2_X1  g1058(.A(new_n1258), .B(KEYINPUT120), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1254), .A2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(G407), .A2(G213), .A3(new_n1261), .ZN(G409));
  INV_X1    g1062(.A(KEYINPUT61), .ZN(new_n1263));
  OAI211_X1 g1063(.A(G378), .B(new_n1226), .C1(new_n1194), .C2(new_n1199), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1198), .A2(new_n1169), .A3(new_n984), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1187), .A2(new_n1191), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1225), .B1(new_n1266), .B2(new_n731), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1265), .A2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(new_n1252), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1264), .A2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(KEYINPUT121), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1258), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT121), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1264), .A2(new_n1273), .A3(new_n1269), .ZN(new_n1274));
  NOR3_X1   g1074(.A1(new_n1126), .A2(new_n1118), .A3(new_n1128), .ZN(new_n1275));
  OAI211_X1 g1075(.A(new_n682), .B(new_n1129), .C1(new_n1275), .C2(KEYINPUT60), .ZN(new_n1276));
  AND2_X1   g1076(.A1(new_n1275), .A2(KEYINPUT60), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1247), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1278), .A2(G384), .ZN(new_n1279));
  OAI211_X1 g1079(.A(new_n852), .B(new_n1247), .C1(new_n1276), .C2(new_n1277), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1271), .A2(new_n1272), .A3(new_n1274), .A4(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT125), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1283), .B1(new_n1270), .B2(new_n1259), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  AOI211_X1 g1085(.A(KEYINPUT125), .B(new_n1260), .C1(new_n1264), .C2(new_n1269), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1285), .A2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(G2897), .ZN(new_n1289));
  NOR3_X1   g1089(.A1(new_n1281), .A2(new_n1289), .A3(new_n1259), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT123), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT122), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1272), .B1(new_n1293), .B2(new_n1289), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1294), .B1(new_n1293), .B2(new_n1289), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1292), .B1(new_n1281), .B2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1295), .ZN(new_n1297));
  AOI211_X1 g1097(.A(KEYINPUT123), .B(new_n1297), .C1(new_n1279), .C2(new_n1280), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1291), .B1(new_n1296), .B2(new_n1298), .ZN(new_n1299));
  OAI221_X1 g1099(.A(new_n1263), .B1(new_n1282), .B2(KEYINPUT62), .C1(new_n1288), .C2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT62), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1301), .B1(new_n1288), .B2(new_n1281), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1098), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1303), .B1(new_n1001), .B2(new_n1031), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1000), .A2(new_n997), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1305), .A2(new_n982), .A3(new_n979), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(G390), .A2(new_n1306), .A3(new_n1030), .ZN(new_n1307));
  XNOR2_X1  g1107(.A(G393), .B(new_n798), .ZN(new_n1308));
  AND3_X1   g1108(.A1(new_n1304), .A2(new_n1307), .A3(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1308), .B1(new_n1304), .B2(new_n1307), .ZN(new_n1310));
  OAI22_X1  g1110(.A1(new_n1300), .A2(new_n1302), .B1(new_n1309), .B2(new_n1310), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1271), .A2(new_n1272), .A3(new_n1274), .ZN(new_n1312));
  NOR2_X1   g1112(.A1(new_n1296), .A2(new_n1298), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(new_n1313), .A2(new_n1290), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT124), .ZN(new_n1315));
  AND3_X1   g1115(.A1(new_n1312), .A2(new_n1314), .A3(new_n1315), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1315), .B1(new_n1312), .B2(new_n1314), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT63), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1282), .A2(new_n1319), .ZN(new_n1320));
  OAI211_X1 g1120(.A(KEYINPUT63), .B(new_n1281), .C1(new_n1284), .C2(new_n1286), .ZN(new_n1321));
  NOR3_X1   g1121(.A1(new_n1309), .A2(new_n1310), .A3(KEYINPUT61), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1320), .A2(new_n1321), .A3(new_n1322), .ZN(new_n1323));
  NOR3_X1   g1123(.A1(new_n1318), .A2(KEYINPUT126), .A3(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT126), .ZN(new_n1325));
  AND3_X1   g1125(.A1(new_n1320), .A2(new_n1321), .A3(new_n1322), .ZN(new_n1326));
  AND3_X1   g1126(.A1(new_n1264), .A2(new_n1273), .A3(new_n1269), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1273), .B1(new_n1264), .B2(new_n1269), .ZN(new_n1328));
  NOR3_X1   g1128(.A1(new_n1327), .A2(new_n1328), .A3(new_n1258), .ZN(new_n1329));
  OAI21_X1  g1129(.A(KEYINPUT124), .B1(new_n1329), .B2(new_n1299), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1312), .A2(new_n1314), .A3(new_n1315), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1330), .A2(new_n1331), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1325), .B1(new_n1326), .B2(new_n1332), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1311), .B1(new_n1324), .B2(new_n1333), .ZN(G405));
  NOR2_X1   g1134(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1335));
  XOR2_X1   g1135(.A(new_n1335), .B(new_n1281), .Z(new_n1336));
  AOI21_X1  g1136(.A(new_n1253), .B1(new_n1200), .B2(new_n1226), .ZN(new_n1337));
  INV_X1    g1137(.A(new_n1264), .ZN(new_n1338));
  OAI21_X1  g1138(.A(KEYINPUT127), .B1(new_n1337), .B2(new_n1338), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1339), .B1(KEYINPUT127), .B2(new_n1337), .ZN(new_n1340));
  XNOR2_X1  g1140(.A(new_n1336), .B(new_n1340), .ZN(G402));
endmodule


