//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 0 0 1 0 0 1 0 1 0 1 1 1 1 1 1 0 0 0 0 0 0 1 1 1 0 0 1 0 0 0 0 0 1 0 0 1 1 1 0 1 1 0 1 0 0 1 0 1 1 1 1 0 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n808, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n840, new_n841, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n896, new_n897, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n973, new_n974, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1012, new_n1013;
  INV_X1    g000(.A(G230gat), .ZN(new_n202));
  INV_X1    g001(.A(G233gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G85gat), .A2(G92gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(KEYINPUT7), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT100), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n207), .B(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT101), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n210), .B1(new_n206), .B2(KEYINPUT7), .ZN(new_n211));
  OR3_X1    g010(.A1(new_n206), .A2(new_n210), .A3(KEYINPUT7), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n209), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(G99gat), .A2(G106gat), .ZN(new_n214));
  INV_X1    g013(.A(G85gat), .ZN(new_n215));
  INV_X1    g014(.A(G92gat), .ZN(new_n216));
  AOI22_X1  g015(.A1(KEYINPUT8), .A2(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n213), .A2(new_n217), .ZN(new_n218));
  XOR2_X1   g017(.A(G99gat), .B(G106gat), .Z(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(G57gat), .B(G64gat), .ZN(new_n221));
  AOI21_X1  g020(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n222));
  OR2_X1    g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  XOR2_X1   g022(.A(G71gat), .B(G78gat), .Z(new_n224));
  XNOR2_X1  g023(.A(new_n223), .B(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(new_n219), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n213), .A2(new_n227), .A3(new_n217), .ZN(new_n228));
  AND3_X1   g027(.A1(new_n220), .A2(new_n226), .A3(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT102), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n227), .B1(new_n213), .B2(new_n217), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n220), .A2(new_n230), .A3(new_n228), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n233), .A2(new_n234), .A3(new_n225), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(KEYINPUT104), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT104), .ZN(new_n237));
  NAND4_X1  g036(.A1(new_n233), .A2(new_n234), .A3(new_n237), .A4(new_n225), .ZN(new_n238));
  AOI211_X1 g037(.A(KEYINPUT10), .B(new_n229), .C1(new_n236), .C2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT10), .ZN(new_n240));
  AOI211_X1 g039(.A(new_n240), .B(new_n225), .C1(new_n234), .C2(new_n233), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n205), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(G120gat), .B(G148gat), .ZN(new_n243));
  XNOR2_X1  g042(.A(G176gat), .B(G204gat), .ZN(new_n244));
  XOR2_X1   g043(.A(new_n243), .B(new_n244), .Z(new_n245));
  AOI21_X1  g044(.A(new_n229), .B1(new_n236), .B2(new_n238), .ZN(new_n246));
  OAI211_X1 g045(.A(new_n242), .B(new_n245), .C1(new_n205), .C2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n245), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n246), .A2(new_n240), .ZN(new_n249));
  INV_X1    g048(.A(new_n241), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n204), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n246), .A2(new_n205), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n248), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n247), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT21), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n225), .A2(new_n256), .ZN(new_n257));
  XOR2_X1   g056(.A(G127gat), .B(G155gat), .Z(new_n258));
  XNOR2_X1  g057(.A(new_n257), .B(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(G15gat), .B(G22gat), .ZN(new_n260));
  OR2_X1    g059(.A1(new_n260), .A2(G1gat), .ZN(new_n261));
  AOI21_X1  g060(.A(G8gat), .B1(new_n261), .B2(KEYINPUT94), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT16), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n260), .B1(new_n263), .B2(G1gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n261), .A2(new_n264), .ZN(new_n265));
  OR2_X1    g064(.A1(new_n262), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n262), .A2(new_n265), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n268), .B1(new_n256), .B2(new_n225), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n259), .B(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(G231gat), .A2(G233gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n271), .B(KEYINPUT99), .ZN(new_n272));
  XOR2_X1   g071(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n273));
  XNOR2_X1  g072(.A(new_n272), .B(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(G183gat), .B(G211gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n274), .B(new_n275), .ZN(new_n276));
  XOR2_X1   g075(.A(new_n270), .B(new_n276), .Z(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  AOI21_X1  g077(.A(KEYINPUT15), .B1(G43gat), .B2(G50gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(KEYINPUT92), .B(G50gat), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n279), .B1(new_n280), .B2(G43gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(KEYINPUT93), .ZN(new_n282));
  XNOR2_X1  g081(.A(G43gat), .B(G50gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(KEYINPUT15), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(G29gat), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n286), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n287));
  XOR2_X1   g086(.A(KEYINPUT14), .B(G29gat), .Z(new_n288));
  OAI21_X1  g087(.A(new_n287), .B1(new_n288), .B2(G36gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n285), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n289), .B1(new_n281), .B2(KEYINPUT93), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(new_n284), .ZN(new_n292));
  AND3_X1   g091(.A1(new_n290), .A2(new_n292), .A3(KEYINPUT17), .ZN(new_n293));
  AOI21_X1  g092(.A(KEYINPUT17), .B1(new_n290), .B2(new_n292), .ZN(new_n294));
  OAI211_X1 g093(.A(new_n233), .B(new_n234), .C1(new_n293), .C2(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(G190gat), .B(G218gat), .ZN(new_n296));
  AND2_X1   g095(.A1(G232gat), .A2(G233gat), .ZN(new_n297));
  AOI22_X1  g096(.A1(new_n296), .A2(KEYINPUT103), .B1(KEYINPUT41), .B2(new_n297), .ZN(new_n298));
  AND2_X1   g097(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n290), .A2(new_n292), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n233), .ZN(new_n302));
  INV_X1    g101(.A(new_n234), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n299), .A2(new_n304), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n296), .A2(KEYINPUT103), .ZN(new_n306));
  AND2_X1   g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n305), .A2(new_n306), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n297), .A2(KEYINPUT41), .ZN(new_n309));
  XNOR2_X1  g108(.A(G134gat), .B(G162gat), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n309), .B(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  OR3_X1    g111(.A1(new_n307), .A2(new_n308), .A3(new_n312), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n312), .B1(new_n307), .B2(new_n308), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n255), .A2(new_n278), .A3(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT84), .ZN(new_n317));
  XNOR2_X1  g116(.A(G78gat), .B(G106gat), .ZN(new_n318));
  XNOR2_X1  g117(.A(new_n318), .B(G22gat), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  AND2_X1   g119(.A1(G228gat), .A2(G233gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(G155gat), .A2(G162gat), .ZN(new_n322));
  OR2_X1    g121(.A1(G155gat), .A2(G162gat), .ZN(new_n323));
  XNOR2_X1  g122(.A(G141gat), .B(G148gat), .ZN(new_n324));
  OAI211_X1 g123(.A(new_n322), .B(new_n323), .C1(new_n324), .C2(KEYINPUT2), .ZN(new_n325));
  INV_X1    g124(.A(G141gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(G148gat), .ZN(new_n327));
  INV_X1    g126(.A(G148gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(G141gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(G155gat), .B(G162gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n322), .A2(KEYINPUT2), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n330), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n325), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(G197gat), .B(G204gat), .ZN(new_n336));
  INV_X1    g135(.A(G218gat), .ZN(new_n337));
  INV_X1    g136(.A(G211gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(KEYINPUT77), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT77), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(G211gat), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n337), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(KEYINPUT76), .B(KEYINPUT22), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n336), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(KEYINPUT78), .ZN(new_n345));
  XNOR2_X1  g144(.A(G211gat), .B(G218gat), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT29), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n344), .A2(KEYINPUT78), .A3(new_n346), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n348), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT3), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n335), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n325), .A2(new_n352), .A3(new_n333), .ZN(new_n354));
  AOI22_X1  g153(.A1(new_n348), .A2(new_n350), .B1(new_n349), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n321), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n355), .A2(new_n321), .ZN(new_n357));
  OR2_X1    g156(.A1(new_n344), .A2(new_n346), .ZN(new_n358));
  AOI21_X1  g157(.A(KEYINPUT29), .B1(new_n344), .B2(new_n346), .ZN(new_n359));
  AOI21_X1  g158(.A(KEYINPUT3), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n357), .B1(new_n335), .B2(new_n360), .ZN(new_n361));
  XNOR2_X1  g160(.A(KEYINPUT31), .B(G50gat), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  AND3_X1   g162(.A1(new_n356), .A2(new_n361), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n363), .B1(new_n356), .B2(new_n361), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n320), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n356), .A2(new_n361), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(new_n362), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n356), .A2(new_n361), .A3(new_n363), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n368), .A2(new_n319), .A3(new_n369), .ZN(new_n370));
  AND2_X1   g169(.A1(new_n366), .A2(new_n370), .ZN(new_n371));
  XOR2_X1   g170(.A(G8gat), .B(G36gat), .Z(new_n372));
  XNOR2_X1  g171(.A(new_n372), .B(KEYINPUT80), .ZN(new_n373));
  XNOR2_X1  g172(.A(G64gat), .B(G92gat), .ZN(new_n374));
  XOR2_X1   g173(.A(new_n373), .B(new_n374), .Z(new_n375));
  INV_X1    g174(.A(new_n348), .ZN(new_n376));
  INV_X1    g175(.A(new_n350), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT79), .ZN(new_n379));
  NAND2_X1  g178(.A1(G226gat), .A2(G233gat), .ZN(new_n380));
  XNOR2_X1  g179(.A(KEYINPUT68), .B(G190gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(KEYINPUT27), .B(G183gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT70), .ZN(new_n384));
  AND2_X1   g183(.A1(new_n384), .A2(KEYINPUT28), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n384), .A2(KEYINPUT28), .ZN(new_n386));
  NOR3_X1   g185(.A1(new_n383), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  AND2_X1   g186(.A1(new_n383), .A2(new_n385), .ZN(new_n388));
  NAND2_X1  g187(.A1(G169gat), .A2(G176gat), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  NOR2_X1   g189(.A1(G169gat), .A2(G176gat), .ZN(new_n391));
  OR3_X1    g190(.A1(new_n390), .A2(new_n391), .A3(KEYINPUT26), .ZN(new_n392));
  NAND2_X1  g191(.A1(G183gat), .A2(G190gat), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n391), .A2(KEYINPUT26), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  NOR3_X1   g194(.A1(new_n387), .A2(new_n388), .A3(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(G183gat), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT24), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n398), .A2(new_n397), .ZN(new_n399));
  AOI22_X1  g198(.A1(new_n381), .A2(new_n397), .B1(G190gat), .B2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT67), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT66), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n393), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(KEYINPUT66), .A2(G183gat), .A3(G190gat), .ZN(new_n404));
  AND4_X1   g203(.A1(new_n401), .A2(new_n403), .A3(new_n398), .A4(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(KEYINPUT24), .B1(new_n393), .B2(new_n402), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n401), .B1(new_n406), .B2(new_n404), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n400), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(KEYINPUT69), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT69), .ZN(new_n410));
  OAI211_X1 g209(.A(new_n400), .B(new_n410), .C1(new_n405), .C2(new_n407), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n391), .A2(KEYINPUT23), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT23), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n413), .B1(G169gat), .B2(G176gat), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n412), .A2(new_n389), .A3(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT25), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n409), .A2(new_n411), .A3(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT65), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n393), .A2(new_n398), .ZN(new_n420));
  NAND3_X1  g219(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n421));
  INV_X1    g220(.A(G190gat), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n397), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n420), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n415), .B1(new_n419), .B2(new_n424), .ZN(new_n425));
  OR2_X1    g224(.A1(new_n424), .A2(new_n419), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(new_n416), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n396), .B1(new_n418), .B2(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n380), .B1(new_n429), .B2(KEYINPUT29), .ZN(new_n430));
  AOI21_X1  g229(.A(KEYINPUT25), .B1(new_n425), .B2(new_n426), .ZN(new_n431));
  OR2_X1    g230(.A1(new_n415), .A2(new_n416), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n432), .B1(new_n408), .B2(KEYINPUT69), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n431), .B1(new_n433), .B2(new_n411), .ZN(new_n434));
  OAI211_X1 g233(.A(G226gat), .B(G233gat), .C1(new_n434), .C2(new_n396), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n379), .B1(new_n430), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n349), .B1(new_n434), .B2(new_n396), .ZN(new_n437));
  AOI21_X1  g236(.A(KEYINPUT79), .B1(new_n437), .B2(new_n380), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n378), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n422), .A2(KEYINPUT68), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT68), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(G190gat), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n440), .A2(new_n442), .A3(new_n397), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(new_n421), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n403), .A2(new_n398), .A3(new_n404), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(KEYINPUT67), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n406), .A2(new_n401), .A3(new_n404), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n444), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n417), .B1(new_n448), .B2(new_n410), .ZN(new_n449));
  INV_X1    g248(.A(new_n411), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n428), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n396), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n380), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n453), .B1(new_n380), .B2(new_n437), .ZN(new_n454));
  INV_X1    g253(.A(new_n378), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n375), .B1(new_n439), .B2(new_n456), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n457), .A2(KEYINPUT30), .ZN(new_n458));
  XOR2_X1   g257(.A(G1gat), .B(G29gat), .Z(new_n459));
  XNOR2_X1  g258(.A(G57gat), .B(G85gat), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n459), .B(new_n460), .ZN(new_n461));
  XNOR2_X1  g260(.A(KEYINPUT83), .B(KEYINPUT0), .ZN(new_n462));
  XNOR2_X1  g261(.A(new_n461), .B(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(G225gat), .A2(G233gat), .ZN(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  AND3_X1   g265(.A1(new_n330), .A2(new_n331), .A3(new_n332), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n331), .B1(new_n332), .B2(new_n330), .ZN(new_n468));
  OAI21_X1  g267(.A(KEYINPUT3), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT1), .ZN(new_n470));
  INV_X1    g269(.A(G113gat), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n471), .A2(G120gat), .ZN(new_n472));
  INV_X1    g271(.A(G120gat), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n473), .A2(G113gat), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n470), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(KEYINPUT71), .A2(G134gat), .ZN(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  NOR2_X1   g276(.A1(KEYINPUT71), .A2(G134gat), .ZN(new_n478));
  INV_X1    g277(.A(G127gat), .ZN(new_n479));
  NOR3_X1   g278(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(G134gat), .ZN(new_n481));
  OAI21_X1  g280(.A(KEYINPUT72), .B1(new_n481), .B2(G127gat), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT72), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n483), .A2(new_n479), .A3(G134gat), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n475), .B1(new_n480), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n473), .A2(G113gat), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n471), .A2(G120gat), .ZN(new_n488));
  AOI21_X1  g287(.A(KEYINPUT1), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  XNOR2_X1  g288(.A(G127gat), .B(G134gat), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n486), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n469), .A2(new_n354), .A3(new_n492), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n486), .A2(new_n325), .A3(new_n333), .A4(new_n491), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n493), .A2(KEYINPUT4), .A3(new_n494), .ZN(new_n495));
  OR2_X1    g294(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n466), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  AND2_X1   g296(.A1(new_n482), .A2(new_n484), .ZN(new_n498));
  INV_X1    g297(.A(new_n478), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n499), .A2(G127gat), .A3(new_n476), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n489), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(new_n491), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n334), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n465), .B1(new_n503), .B2(new_n494), .ZN(new_n504));
  OAI21_X1  g303(.A(KEYINPUT5), .B1(new_n504), .B2(KEYINPUT82), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT82), .ZN(new_n506));
  AOI211_X1 g305(.A(new_n506), .B(new_n465), .C1(new_n503), .C2(new_n494), .ZN(new_n507));
  NOR3_X1   g306(.A1(new_n497), .A2(new_n505), .A3(new_n507), .ZN(new_n508));
  AOI211_X1 g307(.A(KEYINPUT5), .B(new_n466), .C1(new_n495), .C2(new_n496), .ZN(new_n509));
  OAI211_X1 g308(.A(KEYINPUT6), .B(new_n464), .C1(new_n508), .C2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT5), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n497), .A2(new_n511), .ZN(new_n512));
  OR2_X1    g311(.A1(new_n504), .A2(KEYINPUT82), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n504), .A2(KEYINPUT82), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n513), .A2(KEYINPUT5), .A3(new_n514), .ZN(new_n515));
  OAI211_X1 g314(.A(new_n512), .B(new_n463), .C1(new_n515), .C2(new_n497), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT6), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n505), .A2(new_n507), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n495), .A2(new_n496), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n519), .B1(new_n466), .B2(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n463), .B1(new_n522), .B2(new_n512), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n510), .B1(new_n518), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n439), .A2(new_n456), .A3(new_n375), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n458), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n430), .A2(new_n435), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n528), .A2(new_n378), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n430), .A2(new_n379), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n530), .B1(new_n454), .B2(new_n379), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n529), .B1(new_n531), .B2(new_n378), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT30), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n375), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  OAI21_X1  g334(.A(KEYINPUT81), .B1(new_n532), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n439), .A2(new_n456), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT81), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n537), .A2(new_n538), .A3(new_n534), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n371), .B1(new_n527), .B2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n492), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n542), .B1(new_n434), .B2(new_n396), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n451), .A2(new_n492), .A3(new_n452), .ZN(new_n544));
  NAND2_X1  g343(.A1(G227gat), .A2(G233gat), .ZN(new_n545));
  XOR2_X1   g344(.A(new_n545), .B(KEYINPUT64), .Z(new_n546));
  NAND3_X1  g345(.A1(new_n543), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT32), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(KEYINPUT33), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  XOR2_X1   g349(.A(G71gat), .B(G99gat), .Z(new_n551));
  XNOR2_X1  g350(.A(G15gat), .B(G43gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT74), .ZN(new_n555));
  OR2_X1    g354(.A1(new_n553), .A2(KEYINPUT73), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT33), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n557), .B1(new_n553), .B2(KEYINPUT73), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n548), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  AND3_X1   g358(.A1(new_n547), .A2(new_n555), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n555), .B1(new_n547), .B2(new_n559), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n554), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT75), .ZN(new_n563));
  NOR3_X1   g362(.A1(new_n434), .A2(new_n542), .A3(new_n396), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n492), .B1(new_n451), .B2(new_n452), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n545), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(KEYINPUT34), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n546), .A2(KEYINPUT34), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n569), .B1(new_n543), .B2(new_n544), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n563), .B1(new_n567), .B2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT34), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n543), .A2(new_n544), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n573), .B1(new_n574), .B2(new_n545), .ZN(new_n575));
  NOR3_X1   g374(.A1(new_n575), .A2(KEYINPUT75), .A3(new_n570), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n562), .B1(new_n572), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n547), .A2(new_n559), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(KEYINPUT74), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n547), .A2(new_n555), .A3(new_n559), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  OAI21_X1  g380(.A(KEYINPUT75), .B1(new_n575), .B2(new_n570), .ZN(new_n582));
  AOI22_X1  g381(.A1(new_n543), .A2(new_n544), .B1(G227gat), .B2(G233gat), .ZN(new_n583));
  OAI211_X1 g382(.A(new_n571), .B(new_n563), .C1(new_n573), .C2(new_n583), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n581), .A2(new_n582), .A3(new_n584), .A4(new_n554), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n577), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT36), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n577), .A2(new_n585), .A3(KEYINPUT36), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n317), .B1(new_n541), .B2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT86), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n592), .B1(new_n521), .B2(new_n466), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n521), .A2(new_n592), .A3(new_n466), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n503), .A2(new_n465), .A3(new_n494), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n596), .A2(KEYINPUT88), .A3(KEYINPUT39), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(KEYINPUT39), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT88), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n594), .A2(new_n595), .A3(new_n597), .A4(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(KEYINPUT87), .B(KEYINPUT39), .ZN(new_n602));
  INV_X1    g401(.A(new_n595), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n602), .B1(new_n603), .B2(new_n593), .ZN(new_n604));
  XOR2_X1   g403(.A(new_n463), .B(KEYINPUT85), .Z(new_n605));
  NAND3_X1  g404(.A1(new_n601), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT40), .ZN(new_n607));
  OR2_X1    g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n605), .B1(new_n522), .B2(new_n512), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n609), .B1(new_n606), .B2(new_n607), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n538), .B1(new_n537), .B2(new_n534), .ZN(new_n611));
  AOI211_X1 g410(.A(KEYINPUT81), .B(new_n535), .C1(new_n439), .C2(new_n456), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n533), .B1(new_n532), .B2(new_n375), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(new_n525), .ZN(new_n615));
  OAI211_X1 g414(.A(new_n608), .B(new_n610), .C1(new_n613), .C2(new_n615), .ZN(new_n616));
  OAI211_X1 g415(.A(new_n455), .B(new_n530), .C1(new_n454), .C2(new_n379), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT37), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n618), .B1(new_n528), .B2(new_n378), .ZN(new_n619));
  AOI21_X1  g418(.A(KEYINPUT38), .B1(new_n617), .B2(new_n619), .ZN(new_n620));
  OAI211_X1 g419(.A(new_n620), .B(new_n375), .C1(new_n532), .C2(KEYINPUT37), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n510), .B1(new_n518), .B2(new_n609), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n622), .A2(new_n457), .ZN(new_n623));
  AND3_X1   g422(.A1(new_n439), .A2(KEYINPUT37), .A3(new_n456), .ZN(new_n624));
  AOI21_X1  g423(.A(KEYINPUT37), .B1(new_n439), .B2(new_n456), .ZN(new_n625));
  INV_X1    g424(.A(new_n375), .ZN(new_n626));
  NOR3_X1   g425(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT38), .ZN(new_n628));
  OAI211_X1 g427(.A(new_n621), .B(new_n623), .C1(new_n627), .C2(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n616), .A2(new_n629), .A3(new_n371), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n464), .B1(new_n508), .B2(new_n509), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n631), .A2(new_n517), .A3(new_n516), .ZN(new_n632));
  AOI22_X1  g431(.A1(new_n532), .A2(new_n375), .B1(new_n632), .B2(new_n510), .ZN(new_n633));
  OAI211_X1 g432(.A(new_n633), .B(new_n614), .C1(new_n611), .C2(new_n612), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n366), .A2(new_n370), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AND3_X1   g435(.A1(new_n577), .A2(KEYINPUT36), .A3(new_n585), .ZN(new_n637));
  AOI21_X1  g436(.A(KEYINPUT36), .B1(new_n577), .B2(new_n585), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n636), .A2(new_n639), .A3(KEYINPUT84), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n591), .A2(new_n630), .A3(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT89), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n586), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n577), .A2(new_n585), .A3(KEYINPUT89), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n613), .A2(new_n615), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT35), .ZN(new_n647));
  AND3_X1   g446(.A1(new_n371), .A2(new_n647), .A3(new_n622), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n645), .A2(new_n646), .A3(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT90), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n650), .B1(new_n586), .B2(new_n371), .ZN(new_n651));
  AOI211_X1 g450(.A(KEYINPUT90), .B(new_n635), .C1(new_n577), .C2(new_n585), .ZN(new_n652));
  NOR3_X1   g451(.A1(new_n651), .A2(new_n652), .A3(new_n634), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n649), .B1(new_n653), .B2(new_n647), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n641), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT95), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n268), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n266), .A2(KEYINPUT95), .A3(new_n267), .ZN(new_n658));
  OAI211_X1 g457(.A(new_n657), .B(new_n658), .C1(new_n293), .C2(new_n294), .ZN(new_n659));
  NAND2_X1  g458(.A1(G229gat), .A2(G233gat), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n301), .A2(new_n266), .A3(new_n267), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT18), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND4_X1  g463(.A1(new_n659), .A2(KEYINPUT18), .A3(new_n660), .A4(new_n661), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n268), .A2(new_n300), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n661), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(KEYINPUT96), .B(KEYINPUT13), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(new_n660), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(G113gat), .B(G141gat), .ZN(new_n671));
  XNOR2_X1  g470(.A(KEYINPUT91), .B(G197gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XOR2_X1   g472(.A(KEYINPUT11), .B(G169gat), .Z(new_n674));
  XNOR2_X1  g473(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(KEYINPUT12), .ZN(new_n676));
  NAND4_X1  g475(.A1(new_n664), .A2(new_n665), .A3(new_n670), .A4(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT97), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  AOI22_X1  g478(.A1(new_n662), .A2(new_n663), .B1(new_n667), .B2(new_n669), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n676), .B1(new_n680), .B2(new_n665), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  AOI211_X1 g481(.A(new_n678), .B(new_n676), .C1(new_n680), .C2(new_n665), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n655), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(KEYINPUT98), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT98), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n655), .A2(new_n687), .A3(new_n684), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n316), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n524), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(G1gat), .ZN(G1324gat));
  INV_X1    g491(.A(new_n646), .ZN(new_n693));
  INV_X1    g492(.A(new_n316), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n687), .B1(new_n655), .B2(new_n684), .ZN(new_n695));
  INV_X1    g494(.A(new_n684), .ZN(new_n696));
  AOI211_X1 g495(.A(KEYINPUT98), .B(new_n696), .C1(new_n641), .C2(new_n654), .ZN(new_n697));
  OAI211_X1 g496(.A(new_n693), .B(new_n694), .C1(new_n695), .C2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT105), .ZN(new_n699));
  AND3_X1   g498(.A1(new_n698), .A2(new_n699), .A3(G8gat), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n699), .B1(new_n698), .B2(G8gat), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g501(.A(KEYINPUT16), .B(G8gat), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  NAND4_X1  g503(.A1(new_n689), .A2(KEYINPUT42), .A3(new_n693), .A4(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT42), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n706), .B1(new_n698), .B2(new_n703), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(KEYINPUT106), .B1(new_n702), .B2(new_n708), .ZN(new_n709));
  AND2_X1   g508(.A1(new_n705), .A2(new_n707), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n698), .A2(G8gat), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(KEYINPUT105), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n698), .A2(new_n699), .A3(G8gat), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT106), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n710), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n709), .A2(new_n716), .ZN(G1325gat));
  INV_X1    g516(.A(new_n689), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n639), .B(KEYINPUT107), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(G15gat), .B1(new_n718), .B2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(new_n645), .ZN(new_n722));
  OR2_X1    g521(.A1(new_n722), .A2(G15gat), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n721), .B1(new_n718), .B2(new_n723), .ZN(G1326gat));
  NAND2_X1  g523(.A1(new_n689), .A2(new_n635), .ZN(new_n725));
  XNOR2_X1  g524(.A(KEYINPUT43), .B(G22gat), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n725), .B(new_n726), .ZN(G1327gat));
  INV_X1    g526(.A(KEYINPUT44), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n586), .A2(new_n371), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(KEYINPUT90), .ZN(new_n730));
  INV_X1    g529(.A(new_n634), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n586), .A2(new_n650), .A3(new_n371), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n730), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(KEYINPUT35), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n541), .A2(new_n590), .ZN(new_n735));
  AOI22_X1  g534(.A1(new_n734), .A2(new_n649), .B1(new_n735), .B2(new_n630), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n728), .B1(new_n736), .B2(new_n315), .ZN(new_n737));
  INV_X1    g536(.A(new_n315), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n655), .A2(KEYINPUT44), .A3(new_n738), .ZN(new_n739));
  AND2_X1   g538(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n254), .A2(new_n278), .ZN(new_n741));
  INV_X1    g540(.A(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT110), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n743), .B1(new_n682), .B2(new_n683), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n680), .A2(new_n665), .ZN(new_n745));
  INV_X1    g544(.A(new_n676), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n747), .A2(new_n678), .A3(new_n677), .ZN(new_n748));
  INV_X1    g547(.A(new_n683), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n748), .A2(new_n749), .A3(KEYINPUT110), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n744), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n742), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n740), .A2(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(G29gat), .B1(new_n753), .B2(new_n524), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n686), .A2(new_n688), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n742), .A2(new_n315), .ZN(new_n756));
  AND2_X1   g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n757), .A2(new_n286), .A3(new_n690), .ZN(new_n758));
  XNOR2_X1  g557(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(KEYINPUT109), .ZN(new_n760));
  AND2_X1   g559(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n758), .A2(new_n760), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n754), .B1(new_n761), .B2(new_n762), .ZN(G1328gat));
  INV_X1    g562(.A(G36gat), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n757), .A2(new_n764), .A3(new_n693), .ZN(new_n765));
  OR2_X1    g564(.A1(new_n765), .A2(KEYINPUT46), .ZN(new_n766));
  OAI21_X1  g565(.A(G36gat), .B1(new_n753), .B2(new_n646), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n765), .A2(KEYINPUT46), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n766), .A2(new_n767), .A3(new_n768), .ZN(G1329gat));
  INV_X1    g568(.A(G43gat), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n757), .A2(new_n770), .A3(new_n645), .ZN(new_n771));
  OAI21_X1  g570(.A(G43gat), .B1(new_n753), .B2(new_n639), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n771), .A2(new_n772), .A3(KEYINPUT47), .ZN(new_n773));
  OAI21_X1  g572(.A(G43gat), .B1(new_n753), .B2(new_n720), .ZN(new_n774));
  AND2_X1   g573(.A1(new_n771), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n773), .B1(new_n775), .B2(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g575(.A(new_n280), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n755), .A2(new_n756), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n777), .B1(new_n778), .B2(new_n371), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n635), .A2(new_n280), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n779), .B1(new_n753), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(KEYINPUT48), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT48), .ZN(new_n783));
  OAI211_X1 g582(.A(new_n779), .B(new_n783), .C1(new_n753), .C2(new_n780), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n782), .A2(new_n784), .ZN(G1331gat));
  NAND4_X1  g584(.A1(new_n751), .A2(new_n278), .A3(new_n315), .A4(new_n254), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n736), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(new_n690), .ZN(new_n788));
  XNOR2_X1  g587(.A(KEYINPUT111), .B(G57gat), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n788), .B(new_n789), .ZN(G1332gat));
  OR2_X1    g589(.A1(new_n787), .A2(KEYINPUT112), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n787), .A2(KEYINPUT112), .ZN(new_n792));
  AND2_X1   g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n646), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NOR2_X1   g594(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n796));
  XOR2_X1   g595(.A(new_n795), .B(new_n796), .Z(G1333gat));
  NAND3_X1  g596(.A1(new_n791), .A2(new_n719), .A3(new_n792), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(G71gat), .ZN(new_n799));
  INV_X1    g598(.A(G71gat), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT113), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n801), .B1(new_n787), .B2(new_n645), .ZN(new_n802));
  NOR4_X1   g601(.A1(new_n736), .A2(KEYINPUT113), .A3(new_n722), .A4(new_n786), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n800), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n799), .A2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT50), .ZN(new_n806));
  XNOR2_X1  g605(.A(new_n805), .B(new_n806), .ZN(G1334gat));
  NAND2_X1  g606(.A1(new_n793), .A2(new_n635), .ZN(new_n808));
  XNOR2_X1  g607(.A(new_n808), .B(G78gat), .ZN(G1335gat));
  INV_X1    g608(.A(new_n751), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n810), .A2(new_n278), .A3(new_n255), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n740), .A2(new_n811), .ZN(new_n812));
  OAI21_X1  g611(.A(G85gat), .B1(new_n812), .B2(new_n524), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n630), .A2(new_n735), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n315), .B1(new_n654), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n810), .A2(new_n278), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n815), .A2(KEYINPUT51), .A3(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(KEYINPUT51), .B1(new_n815), .B2(new_n816), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n254), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n690), .A2(new_n215), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n813), .B1(new_n820), .B2(new_n821), .ZN(G1336gat));
  OAI21_X1  g621(.A(G92gat), .B1(new_n812), .B2(new_n646), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT52), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n646), .A2(new_n255), .A3(G92gat), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n825), .B1(new_n818), .B2(new_n819), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n823), .A2(new_n824), .A3(new_n826), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n630), .A2(new_n735), .ZN(new_n828));
  AND4_X1   g627(.A1(new_n540), .A2(new_n648), .A3(new_n614), .A4(new_n525), .ZN(new_n829));
  AOI22_X1  g628(.A1(new_n733), .A2(KEYINPUT35), .B1(new_n829), .B2(new_n645), .ZN(new_n830));
  OAI211_X1 g629(.A(new_n738), .B(new_n816), .C1(new_n828), .C2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT51), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n833), .A2(KEYINPUT114), .A3(new_n817), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT114), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n834), .A2(new_n836), .A3(new_n825), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n823), .A2(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n827), .B1(new_n838), .B2(new_n824), .ZN(G1337gat));
  OAI21_X1  g638(.A(G99gat), .B1(new_n812), .B2(new_n720), .ZN(new_n840));
  OR2_X1    g639(.A1(new_n722), .A2(G99gat), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n840), .B1(new_n820), .B2(new_n841), .ZN(G1338gat));
  NOR2_X1   g641(.A1(new_n371), .A2(G106gat), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n834), .A2(new_n836), .A3(new_n254), .A4(new_n843), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n737), .A2(new_n739), .A3(new_n635), .A4(new_n811), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(G106gat), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(KEYINPUT53), .ZN(new_n848));
  OAI211_X1 g647(.A(new_n254), .B(new_n843), .C1(new_n818), .C2(new_n819), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT53), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n849), .A2(new_n846), .A3(new_n850), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n848), .A2(KEYINPUT115), .A3(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT115), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n850), .B1(new_n844), .B2(new_n846), .ZN(new_n854));
  AND3_X1   g653(.A1(new_n849), .A2(new_n846), .A3(new_n850), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n853), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n852), .A2(new_n856), .ZN(G1339gat));
  NAND4_X1  g656(.A1(new_n751), .A2(new_n278), .A3(new_n255), .A4(new_n315), .ZN(new_n858));
  XOR2_X1   g657(.A(KEYINPUT116), .B(KEYINPUT54), .Z(new_n859));
  AOI21_X1  g658(.A(new_n245), .B1(new_n251), .B2(new_n859), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n249), .A2(new_n204), .A3(new_n250), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n242), .A2(new_n861), .A3(KEYINPUT54), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT55), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n860), .A2(new_n862), .A3(KEYINPUT55), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n865), .A2(new_n247), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n660), .B1(new_n659), .B2(new_n661), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n667), .A2(new_n669), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n675), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n677), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n738), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n867), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n254), .A2(new_n871), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n874), .B1(new_n867), .B2(new_n751), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n873), .B1(new_n875), .B2(new_n315), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n858), .B1(new_n876), .B2(new_n278), .ZN(new_n877));
  AND2_X1   g676(.A1(new_n877), .A2(new_n690), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n651), .A2(new_n652), .ZN(new_n879));
  INV_X1    g678(.A(new_n879), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n880), .A2(new_n693), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n878), .A2(new_n810), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(new_n471), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n693), .A2(new_n524), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n722), .A2(new_n635), .ZN(new_n885));
  AND3_X1   g684(.A1(new_n877), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n886), .A2(G113gat), .A3(new_n684), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n883), .A2(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT117), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n888), .B(new_n889), .ZN(G1340gat));
  AND2_X1   g689(.A1(new_n878), .A2(new_n881), .ZN(new_n891));
  AOI21_X1  g690(.A(G120gat), .B1(new_n891), .B2(new_n254), .ZN(new_n892));
  INV_X1    g691(.A(new_n886), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n893), .A2(new_n473), .A3(new_n255), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n892), .A2(new_n894), .ZN(G1341gat));
  NAND3_X1  g694(.A1(new_n891), .A2(new_n479), .A3(new_n278), .ZN(new_n896));
  OAI21_X1  g695(.A(G127gat), .B1(new_n893), .B2(new_n277), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(G1342gat));
  AOI21_X1  g697(.A(new_n481), .B1(new_n886), .B2(new_n738), .ZN(new_n899));
  NOR3_X1   g698(.A1(new_n315), .A2(new_n478), .A3(new_n477), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n878), .A2(new_n881), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n899), .B1(KEYINPUT56), .B2(new_n901), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n901), .A2(KEYINPUT56), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT118), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n901), .A2(KEYINPUT118), .A3(KEYINPUT56), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n902), .B1(new_n905), .B2(new_n906), .ZN(G1343gat));
  NOR2_X1   g706(.A1(new_n719), .A2(new_n371), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n877), .A2(new_n690), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(KEYINPUT119), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n693), .A2(new_n696), .A3(G141gat), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT119), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n877), .A2(new_n912), .A3(new_n690), .A4(new_n908), .ZN(new_n913));
  AND3_X1   g712(.A1(new_n910), .A2(new_n911), .A3(new_n913), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n865), .A2(new_n684), .A3(new_n247), .A4(new_n866), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n738), .B1(new_n915), .B2(new_n874), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n277), .B1(new_n916), .B2(new_n873), .ZN(new_n917));
  AND2_X1   g716(.A1(new_n917), .A2(new_n858), .ZN(new_n918));
  OAI21_X1  g717(.A(KEYINPUT57), .B1(new_n918), .B2(new_n371), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT57), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n877), .A2(new_n920), .A3(new_n635), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n693), .A2(new_n524), .A3(new_n590), .ZN(new_n922));
  NAND4_X1  g721(.A1(new_n919), .A2(new_n684), .A3(new_n921), .A4(new_n922), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(G141gat), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT120), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n914), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT58), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n910), .A2(new_n911), .A3(new_n913), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n927), .B1(new_n928), .B2(KEYINPUT120), .ZN(new_n929));
  NAND4_X1  g728(.A1(new_n919), .A2(new_n810), .A3(new_n921), .A4(new_n922), .ZN(new_n930));
  INV_X1    g729(.A(new_n909), .ZN(new_n931));
  AOI22_X1  g730(.A1(new_n930), .A2(G141gat), .B1(new_n931), .B2(new_n911), .ZN(new_n932));
  OAI22_X1  g731(.A1(new_n926), .A2(new_n929), .B1(new_n927), .B2(new_n932), .ZN(G1344gat));
  NAND3_X1  g732(.A1(new_n910), .A2(new_n646), .A3(new_n913), .ZN(new_n934));
  OR3_X1    g733(.A1(new_n934), .A2(G148gat), .A3(new_n255), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n919), .A2(new_n921), .A3(new_n922), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n936), .A2(new_n255), .ZN(new_n937));
  NOR3_X1   g736(.A1(new_n937), .A2(KEYINPUT59), .A3(new_n328), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT59), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n877), .A2(new_n635), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(KEYINPUT57), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT121), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n942), .B1(new_n316), .B2(new_n684), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n694), .A2(KEYINPUT121), .A3(new_n696), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n917), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n945), .A2(new_n920), .A3(new_n635), .ZN(new_n946));
  NAND4_X1  g745(.A1(new_n941), .A2(new_n254), .A3(new_n922), .A4(new_n946), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n939), .B1(new_n947), .B2(G148gat), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n935), .B1(new_n938), .B2(new_n948), .ZN(G1345gat));
  NAND4_X1  g748(.A1(new_n919), .A2(new_n278), .A3(new_n921), .A4(new_n922), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(G155gat), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n277), .A2(G155gat), .ZN(new_n952));
  NAND4_X1  g751(.A1(new_n910), .A2(new_n646), .A3(new_n913), .A4(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT122), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n951), .A2(KEYINPUT122), .A3(new_n953), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(G1346gat));
  OAI21_X1  g757(.A(G162gat), .B1(new_n936), .B2(new_n315), .ZN(new_n959));
  OR2_X1    g758(.A1(new_n315), .A2(G162gat), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n959), .B1(new_n934), .B2(new_n960), .ZN(G1347gat));
  AND2_X1   g760(.A1(new_n877), .A2(new_n885), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n646), .A2(new_n690), .ZN(new_n963));
  NAND4_X1  g762(.A1(new_n962), .A2(G169gat), .A3(new_n684), .A4(new_n963), .ZN(new_n964));
  AND2_X1   g763(.A1(new_n877), .A2(new_n524), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n880), .A2(new_n646), .ZN(new_n966));
  AND3_X1   g765(.A1(new_n965), .A2(new_n810), .A3(new_n966), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n964), .B1(new_n967), .B2(G169gat), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT123), .ZN(new_n969));
  XNOR2_X1  g768(.A(new_n968), .B(new_n969), .ZN(G1348gat));
  NAND2_X1  g769(.A1(new_n962), .A2(new_n963), .ZN(new_n971));
  OAI21_X1  g770(.A(G176gat), .B1(new_n971), .B2(new_n255), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n255), .A2(G176gat), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n965), .A2(new_n966), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n972), .A2(new_n974), .ZN(G1349gat));
  OAI21_X1  g774(.A(G183gat), .B1(new_n971), .B2(new_n277), .ZN(new_n976));
  NAND4_X1  g775(.A1(new_n965), .A2(new_n382), .A3(new_n278), .A4(new_n966), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  XNOR2_X1  g777(.A(KEYINPUT124), .B(KEYINPUT60), .ZN(new_n979));
  INV_X1    g778(.A(new_n979), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n976), .A2(new_n977), .A3(new_n979), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n981), .A2(new_n982), .ZN(G1350gat));
  AOI21_X1  g782(.A(new_n422), .B1(KEYINPUT126), .B2(KEYINPUT61), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n984), .B1(new_n971), .B2(new_n315), .ZN(new_n985));
  NOR2_X1   g784(.A1(KEYINPUT126), .A2(KEYINPUT61), .ZN(new_n986));
  OR2_X1    g785(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND4_X1  g786(.A1(new_n965), .A2(new_n381), .A3(new_n738), .A4(new_n966), .ZN(new_n988));
  XNOR2_X1  g787(.A(new_n988), .B(KEYINPUT125), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n985), .A2(new_n986), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n987), .A2(new_n989), .A3(new_n990), .ZN(G1351gat));
  NOR3_X1   g790(.A1(new_n719), .A2(new_n371), .A3(new_n646), .ZN(new_n992));
  NOR2_X1   g791(.A1(new_n751), .A2(G197gat), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n965), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  XOR2_X1   g793(.A(new_n994), .B(KEYINPUT127), .Z(new_n995));
  NOR3_X1   g794(.A1(new_n719), .A2(new_n690), .A3(new_n646), .ZN(new_n996));
  NAND3_X1  g795(.A1(new_n941), .A2(new_n946), .A3(new_n996), .ZN(new_n997));
  OAI21_X1  g796(.A(G197gat), .B1(new_n997), .B2(new_n696), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n995), .A2(new_n998), .ZN(G1352gat));
  NOR2_X1   g798(.A1(new_n255), .A2(G204gat), .ZN(new_n1000));
  NAND3_X1  g799(.A1(new_n965), .A2(new_n992), .A3(new_n1000), .ZN(new_n1001));
  XOR2_X1   g800(.A(new_n1001), .B(KEYINPUT62), .Z(new_n1002));
  OAI21_X1  g801(.A(G204gat), .B1(new_n997), .B2(new_n255), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1002), .A2(new_n1003), .ZN(G1353gat));
  NAND2_X1  g803(.A1(new_n965), .A2(new_n992), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n339), .A2(new_n341), .ZN(new_n1006));
  OR3_X1    g805(.A1(new_n1005), .A2(new_n1006), .A3(new_n277), .ZN(new_n1007));
  NAND4_X1  g806(.A1(new_n941), .A2(new_n278), .A3(new_n946), .A4(new_n996), .ZN(new_n1008));
  AND3_X1   g807(.A1(new_n1008), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1009));
  AOI21_X1  g808(.A(KEYINPUT63), .B1(new_n1008), .B2(G211gat), .ZN(new_n1010));
  OAI21_X1  g809(.A(new_n1007), .B1(new_n1009), .B2(new_n1010), .ZN(G1354gat));
  OAI21_X1  g810(.A(G218gat), .B1(new_n997), .B2(new_n315), .ZN(new_n1012));
  NAND2_X1  g811(.A1(new_n738), .A2(new_n337), .ZN(new_n1013));
  OAI21_X1  g812(.A(new_n1012), .B1(new_n1005), .B2(new_n1013), .ZN(G1355gat));
endmodule


