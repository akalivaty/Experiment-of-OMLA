//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 1 1 1 0 1 0 0 1 0 0 1 0 1 0 1 0 1 0 1 0 0 1 1 0 1 1 0 0 1 0 1 0 1 1 1 1 1 1 1 1 1 1 0 1 0 0 1 0 1 0 1 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:01 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n438, new_n439, new_n446, new_n447, new_n448,
    new_n453, new_n457, new_n458, new_n459, new_n460, new_n461, new_n462,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n576, new_n577, new_n578, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n587, new_n588, new_n589,
    new_n590, new_n591, new_n592, new_n594, new_n595, new_n596, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n632, new_n633, new_n636, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n859, new_n860, new_n861, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT65), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT66), .ZN(new_n437));
  OR2_X1    g012(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g013(.A1(new_n436), .A2(new_n437), .ZN(new_n439));
  NAND2_X1  g014(.A1(new_n438), .A2(new_n439), .ZN(G220));
  INV_X1    g015(.A(G96), .ZN(G221));
  INV_X1    g016(.A(G69), .ZN(G235));
  XNOR2_X1  g017(.A(KEYINPUT67), .B(G120), .ZN(G236));
  INV_X1    g018(.A(G57), .ZN(G237));
  INV_X1    g019(.A(G108), .ZN(G238));
  INV_X1    g020(.A(G2072), .ZN(new_n446));
  INV_X1    g021(.A(G2078), .ZN(new_n447));
  NOR2_X1   g022(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g023(.A1(new_n448), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g024(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g025(.A(KEYINPUT68), .B(G452), .Z(G391));
  AND2_X1   g026(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g027(.A1(G7), .A2(G661), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g029(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g030(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR3_X1   g031(.A1(G218), .A2(G221), .A3(G219), .ZN(new_n457));
  NAND3_X1  g032(.A1(new_n438), .A2(new_n439), .A3(new_n457), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT69), .Z(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT2), .ZN(new_n460));
  NOR4_X1   g035(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n461));
  XOR2_X1   g036(.A(new_n461), .B(KEYINPUT70), .Z(new_n462));
  NOR2_X1   g037(.A1(new_n460), .A2(new_n462), .ZN(G325));
  INV_X1    g038(.A(G325), .ZN(G261));
  AOI22_X1  g039(.A1(new_n460), .A2(G2106), .B1(G567), .B2(new_n462), .ZN(G319));
  OR2_X1    g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(G2105), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G137), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  AND3_X1   g045(.A1(new_n470), .A2(KEYINPUT72), .A3(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(KEYINPUT72), .B1(new_n470), .B2(G2104), .ZN(new_n472));
  OAI21_X1  g047(.A(G101), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT71), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g052(.A1(KEYINPUT71), .A2(G113), .A3(G2104), .ZN(new_n478));
  AND2_X1   g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AND2_X1   g054(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n480));
  NOR2_X1   g055(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n481));
  OAI21_X1  g056(.A(G125), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n470), .B1(new_n479), .B2(new_n482), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n474), .A2(new_n483), .ZN(G160));
  AOI21_X1  g059(.A(new_n470), .B1(new_n466), .B2(new_n467), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  XOR2_X1   g061(.A(new_n486), .B(KEYINPUT73), .Z(new_n487));
  NAND2_X1  g062(.A1(new_n468), .A2(G136), .ZN(new_n488));
  NOR2_X1   g063(.A1(G100), .A2(G2105), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(new_n470), .B2(G112), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n487), .B(new_n488), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  XNOR2_X1  g066(.A(new_n491), .B(KEYINPUT74), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  OAI211_X1 g068(.A(G138), .B(new_n470), .C1(new_n480), .C2(new_n481), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n466), .A2(new_n467), .ZN(new_n497));
  NAND2_X1  g072(.A1(G126), .A2(G2105), .ZN(new_n498));
  NAND2_X1  g073(.A1(KEYINPUT4), .A2(G138), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n498), .B1(new_n499), .B2(G2105), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(G114), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G2105), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT75), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT75), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n505), .A2(new_n502), .A3(G2105), .ZN(new_n506));
  OAI21_X1  g081(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n504), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n496), .A2(new_n501), .A3(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(G164));
  NOR2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  XNOR2_X1  g088(.A(KEYINPUT76), .B(G651), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT6), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  XNOR2_X1  g091(.A(KEYINPUT77), .B(G88), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT5), .ZN(new_n518));
  INV_X1    g093(.A(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(KEYINPUT5), .A2(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n516), .A2(new_n517), .A3(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G651), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(KEYINPUT76), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT76), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G651), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n528), .A2(new_n522), .A3(G62), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n516), .A2(G50), .B1(G75), .B2(new_n528), .ZN(new_n530));
  OAI211_X1 g105(.A(new_n523), .B(new_n529), .C1(new_n530), .C2(new_n519), .ZN(G303));
  INV_X1    g106(.A(G303), .ZN(G166));
  INV_X1    g107(.A(KEYINPUT78), .ZN(new_n533));
  INV_X1    g108(.A(new_n521), .ZN(new_n534));
  NOR2_X1   g109(.A1(KEYINPUT5), .A2(G543), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(G63), .A2(G651), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n533), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND4_X1  g113(.A1(new_n522), .A2(KEYINPUT78), .A3(G63), .A4(G651), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n516), .A2(G89), .A3(new_n522), .ZN(new_n541));
  NAND3_X1  g116(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n542), .B(KEYINPUT7), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n540), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(G51), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT79), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n512), .B1(new_n528), .B2(KEYINPUT6), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n548), .B2(new_n519), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n516), .A2(KEYINPUT79), .A3(G543), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n545), .B1(new_n546), .B2(new_n551), .ZN(G286));
  INV_X1    g127(.A(G286), .ZN(G168));
  NAND3_X1  g128(.A1(new_n549), .A2(G52), .A3(new_n550), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n528), .A2(KEYINPUT6), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n536), .B1(new_n555), .B2(new_n513), .ZN(new_n556));
  NAND2_X1  g131(.A1(G77), .A2(G543), .ZN(new_n557));
  INV_X1    g132(.A(G64), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n557), .B1(new_n536), .B2(new_n558), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n556), .A2(G90), .B1(new_n559), .B2(new_n528), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n554), .A2(new_n560), .ZN(G301));
  INV_X1    g136(.A(G301), .ZN(G171));
  NAND3_X1  g137(.A1(new_n549), .A2(G43), .A3(new_n550), .ZN(new_n563));
  OAI21_X1  g138(.A(G56), .B1(new_n534), .B2(new_n535), .ZN(new_n564));
  NAND2_X1  g139(.A1(G68), .A2(G543), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n514), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n566), .B1(new_n556), .B2(G81), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(KEYINPUT80), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT80), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n563), .A2(new_n567), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(G860), .ZN(G153));
  NAND4_X1  g149(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g150(.A1(G1), .A2(G3), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n576), .B(KEYINPUT8), .ZN(new_n577));
  NAND4_X1  g152(.A1(G319), .A2(G483), .A3(G661), .A4(new_n577), .ZN(new_n578));
  XOR2_X1   g153(.A(new_n578), .B(KEYINPUT81), .Z(G188));
  INV_X1    g154(.A(G53), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT82), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n580), .B1(new_n581), .B2(KEYINPUT9), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n516), .A2(G543), .A3(new_n582), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n581), .A2(KEYINPUT9), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n584), .ZN(new_n586));
  NAND4_X1  g161(.A1(new_n516), .A2(G543), .A3(new_n586), .A4(new_n582), .ZN(new_n587));
  NAND2_X1  g162(.A1(G78), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G65), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n536), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n590), .A2(G651), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n516), .A2(G91), .A3(new_n522), .ZN(new_n592));
  NAND4_X1  g167(.A1(new_n585), .A2(new_n587), .A3(new_n591), .A4(new_n592), .ZN(G299));
  NAND2_X1  g168(.A1(new_n556), .A2(G87), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n516), .A2(G49), .A3(G543), .ZN(new_n595));
  OAI21_X1  g170(.A(G651), .B1(new_n522), .B2(G74), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(G288));
  NAND3_X1  g172(.A1(new_n516), .A2(G48), .A3(G543), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n515), .B1(new_n525), .B2(new_n527), .ZN(new_n599));
  OAI211_X1 g174(.A(G86), .B(new_n522), .C1(new_n599), .C2(new_n512), .ZN(new_n600));
  INV_X1    g175(.A(G61), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n601), .B1(new_n520), .B2(new_n521), .ZN(new_n602));
  AND2_X1   g177(.A1(G73), .A2(G543), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n528), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n598), .A2(new_n600), .A3(new_n604), .ZN(G305));
  NAND2_X1  g180(.A1(G72), .A2(G543), .ZN(new_n606));
  INV_X1    g181(.A(G60), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n536), .B2(new_n607), .ZN(new_n608));
  OR2_X1    g183(.A1(new_n608), .A2(KEYINPUT83), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n514), .B1(new_n608), .B2(KEYINPUT83), .ZN(new_n610));
  XNOR2_X1  g185(.A(KEYINPUT84), .B(G85), .ZN(new_n611));
  AOI22_X1  g186(.A1(new_n609), .A2(new_n610), .B1(new_n556), .B2(new_n611), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n549), .A2(G47), .A3(new_n550), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(new_n613), .ZN(G290));
  INV_X1    g189(.A(G868), .ZN(new_n615));
  NOR2_X1   g190(.A1(G301), .A2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT10), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n516), .A2(new_n522), .ZN(new_n618));
  INV_X1    g193(.A(G92), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n556), .A2(KEYINPUT10), .A3(G92), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n549), .A2(G54), .A3(new_n550), .ZN(new_n623));
  NAND2_X1  g198(.A1(G79), .A2(G543), .ZN(new_n624));
  INV_X1    g199(.A(G66), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(new_n536), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(G651), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n622), .A2(new_n623), .A3(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT85), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n616), .B1(new_n629), .B2(new_n615), .ZN(G284));
  AOI21_X1  g205(.A(new_n616), .B1(new_n629), .B2(new_n615), .ZN(G321));
  NOR2_X1   g206(.A1(G286), .A2(new_n615), .ZN(new_n632));
  XOR2_X1   g207(.A(G299), .B(KEYINPUT86), .Z(new_n633));
  AOI21_X1  g208(.A(new_n632), .B1(new_n633), .B2(new_n615), .ZN(G297));
  AOI21_X1  g209(.A(new_n632), .B1(new_n633), .B2(new_n615), .ZN(G280));
  INV_X1    g210(.A(G559), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n629), .B1(new_n636), .B2(G860), .ZN(G148));
  NAND2_X1  g212(.A1(new_n629), .A2(new_n636), .ZN(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n639), .A2(G868), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n573), .A2(new_n615), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(KEYINPUT11), .Z(G282));
  INV_X1    g218(.A(new_n642), .ZN(G323));
  OR2_X1    g219(.A1(new_n471), .A2(new_n472), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n645), .A2(new_n497), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(KEYINPUT12), .Z(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(KEYINPUT13), .Z(new_n648));
  INV_X1    g223(.A(G2100), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n648), .A2(new_n649), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n468), .A2(G135), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n485), .A2(G123), .ZN(new_n653));
  NOR2_X1   g228(.A1(G99), .A2(G2105), .ZN(new_n654));
  OAI21_X1  g229(.A(G2104), .B1(new_n470), .B2(G111), .ZN(new_n655));
  OAI211_X1 g230(.A(new_n652), .B(new_n653), .C1(new_n654), .C2(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(G2096), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n650), .A2(new_n651), .A3(new_n658), .ZN(G156));
  XOR2_X1   g234(.A(G2451), .B(G2454), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT16), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1341), .B(G1348), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G2443), .B(G2446), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2427), .B(G2438), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(G2430), .ZN(new_n667));
  XNOR2_X1  g242(.A(KEYINPUT15), .B(G2435), .ZN(new_n668));
  OR2_X1    g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n667), .A2(new_n668), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n669), .A2(new_n670), .A3(KEYINPUT14), .ZN(new_n671));
  OR2_X1    g246(.A1(new_n665), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n665), .A2(new_n671), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n672), .A2(G14), .A3(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(G401));
  XNOR2_X1  g250(.A(G2084), .B(G2090), .ZN(new_n676));
  XNOR2_X1  g251(.A(G2067), .B(G2678), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT87), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g254(.A1(G2072), .A2(G2078), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n448), .A2(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n676), .B1(new_n679), .B2(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(KEYINPUT89), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n681), .B(KEYINPUT17), .Z(new_n685));
  AOI22_X1  g260(.A1(new_n683), .A2(new_n684), .B1(new_n679), .B2(new_n685), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n686), .B1(new_n684), .B2(new_n683), .ZN(new_n687));
  OR3_X1    g262(.A1(new_n685), .A2(new_n679), .A3(new_n676), .ZN(new_n688));
  NOR3_X1   g263(.A1(new_n678), .A2(new_n676), .A3(new_n681), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT88), .B(KEYINPUT18), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n687), .A2(new_n688), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(new_n657), .ZN(new_n693));
  OR2_X1    g268(.A1(new_n693), .A2(G2100), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(G2100), .ZN(new_n695));
  AND2_X1   g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(G227));
  XOR2_X1   g272(.A(G1971), .B(G1976), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT19), .ZN(new_n699));
  XOR2_X1   g274(.A(G1956), .B(G2474), .Z(new_n700));
  XOR2_X1   g275(.A(G1961), .B(G1966), .Z(new_n701));
  AND2_X1   g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT20), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n700), .A2(new_n701), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n702), .A2(new_n706), .ZN(new_n707));
  MUX2_X1   g282(.A(new_n707), .B(new_n706), .S(new_n699), .Z(new_n708));
  NOR2_X1   g283(.A1(new_n705), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(G1986), .ZN(new_n710));
  XOR2_X1   g285(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(G1986), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n709), .B(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(new_n711), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n713), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g292(.A(G1991), .B(G1996), .ZN(new_n718));
  INV_X1    g293(.A(G1981), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n717), .B(new_n720), .ZN(G229));
  INV_X1    g296(.A(G29), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(G35), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G162), .B2(new_n722), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n724), .A2(KEYINPUT29), .ZN(new_n725));
  INV_X1    g300(.A(G2090), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n724), .A2(KEYINPUT29), .ZN(new_n727));
  AND3_X1   g302(.A1(new_n725), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n726), .B1(new_n725), .B2(new_n727), .ZN(new_n729));
  INV_X1    g304(.A(G16), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n730), .A2(G19), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(new_n573), .B2(new_n730), .ZN(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(G1341), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NOR3_X1   g310(.A1(new_n728), .A2(new_n729), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n722), .A2(G33), .ZN(new_n737));
  AOI22_X1  g312(.A1(new_n497), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n738), .A2(new_n470), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n468), .A2(G139), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT25), .ZN(new_n743));
  NOR3_X1   g318(.A1(new_n739), .A2(new_n741), .A3(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT97), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n737), .B1(new_n746), .B2(new_n722), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(new_n446), .ZN(new_n748));
  INV_X1    g323(.A(G1966), .ZN(new_n749));
  NOR2_X1   g324(.A1(G168), .A2(new_n730), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(new_n730), .B2(G21), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n748), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n730), .A2(G20), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT23), .Z(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(G299), .B2(G16), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(G1956), .Z(new_n756));
  NAND2_X1  g331(.A1(new_n722), .A2(G26), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(KEYINPUT28), .Z(new_n758));
  NAND2_X1  g333(.A1(new_n485), .A2(G128), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT96), .Z(new_n760));
  OR2_X1    g335(.A1(G104), .A2(G2105), .ZN(new_n761));
  INV_X1    g336(.A(G2104), .ZN(new_n762));
  INV_X1    g337(.A(G116), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n762), .B1(new_n763), .B2(G2105), .ZN(new_n764));
  AOI22_X1  g339(.A1(new_n468), .A2(G140), .B1(new_n761), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n760), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n758), .B1(new_n766), .B2(G29), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(G2067), .ZN(new_n768));
  NOR2_X1   g343(.A1(G164), .A2(new_n722), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(G27), .B2(new_n722), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n770), .A2(new_n447), .ZN(new_n771));
  AND2_X1   g346(.A1(new_n722), .A2(G32), .ZN(new_n772));
  XOR2_X1   g347(.A(KEYINPUT98), .B(KEYINPUT26), .Z(new_n773));
  NAND3_X1  g348(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  AOI22_X1  g350(.A1(G129), .A2(new_n485), .B1(new_n468), .B2(G141), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n645), .A2(G105), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n775), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n772), .B1(new_n778), .B2(G29), .ZN(new_n779));
  XNOR2_X1  g354(.A(KEYINPUT27), .B(G1996), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n771), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n779), .A2(new_n780), .ZN(new_n782));
  AND2_X1   g357(.A1(KEYINPUT24), .A2(G34), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n722), .B1(KEYINPUT24), .B2(G34), .ZN(new_n784));
  OAI22_X1  g359(.A1(G160), .A2(new_n722), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  AND2_X1   g360(.A1(new_n785), .A2(G2084), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n785), .A2(G2084), .ZN(new_n787));
  NOR3_X1   g362(.A1(new_n782), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  XOR2_X1   g363(.A(KEYINPUT31), .B(G11), .Z(new_n789));
  INV_X1    g364(.A(G28), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n790), .A2(KEYINPUT30), .ZN(new_n791));
  AOI21_X1  g366(.A(G29), .B1(new_n790), .B2(KEYINPUT30), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n789), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(new_n656), .B2(new_n722), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(new_n770), .B2(new_n447), .ZN(new_n795));
  NAND4_X1  g370(.A1(new_n768), .A2(new_n781), .A3(new_n788), .A4(new_n795), .ZN(new_n796));
  NOR3_X1   g371(.A1(new_n752), .A2(new_n756), .A3(new_n796), .ZN(new_n797));
  NOR2_X1   g372(.A1(G171), .A2(new_n730), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(G5), .B2(new_n730), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  AOI22_X1  g375(.A1(new_n749), .A2(new_n751), .B1(new_n800), .B2(G1961), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G1961), .B2(new_n800), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(new_n734), .B2(new_n733), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n730), .A2(G4), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(new_n629), .B2(new_n730), .ZN(new_n805));
  INV_X1    g380(.A(G1348), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NAND4_X1  g382(.A1(new_n736), .A2(new_n797), .A3(new_n803), .A4(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n730), .A2(G24), .ZN(new_n809));
  INV_X1    g384(.A(G290), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n809), .B1(new_n810), .B2(new_n730), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n811), .A2(G1986), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n811), .A2(G1986), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n814), .A2(KEYINPUT92), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT92), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n812), .A2(new_n816), .A3(new_n813), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n468), .A2(G131), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n485), .A2(G119), .ZN(new_n819));
  NOR2_X1   g394(.A1(G95), .A2(G2105), .ZN(new_n820));
  OAI21_X1  g395(.A(G2104), .B1(new_n470), .B2(G107), .ZN(new_n821));
  OAI211_X1 g396(.A(new_n818), .B(new_n819), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT90), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  MUX2_X1   g399(.A(G25), .B(new_n824), .S(G29), .Z(new_n825));
  XNOR2_X1  g400(.A(KEYINPUT35), .B(G1991), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT91), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n825), .B(new_n827), .Z(new_n828));
  NAND3_X1  g403(.A1(new_n815), .A2(new_n817), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n730), .A2(G6), .ZN(new_n830));
  INV_X1    g405(.A(G305), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n830), .B1(new_n831), .B2(new_n730), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT32), .ZN(new_n833));
  XOR2_X1   g408(.A(KEYINPUT93), .B(G1981), .Z(new_n834));
  OR2_X1    g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n833), .A2(new_n834), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n730), .A2(G22), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(G166), .B2(new_n730), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(G1971), .Z(new_n839));
  NAND2_X1  g414(.A1(new_n730), .A2(G23), .ZN(new_n840));
  INV_X1    g415(.A(G288), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n840), .B1(new_n841), .B2(new_n730), .ZN(new_n842));
  XNOR2_X1  g417(.A(KEYINPUT33), .B(G1976), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT94), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n842), .B(new_n844), .ZN(new_n845));
  NAND4_X1  g420(.A1(new_n835), .A2(new_n836), .A3(new_n839), .A4(new_n845), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n846), .A2(KEYINPUT34), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n829), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(KEYINPUT95), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT95), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n850), .B1(new_n829), .B2(new_n847), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n846), .A2(KEYINPUT34), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(KEYINPUT36), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT36), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n852), .A2(new_n856), .A3(new_n853), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n808), .B1(new_n855), .B2(new_n857), .ZN(G311));
  INV_X1    g433(.A(new_n808), .ZN(new_n859));
  INV_X1    g434(.A(new_n857), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n856), .B1(new_n852), .B2(new_n853), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n859), .B1(new_n860), .B2(new_n861), .ZN(G150));
  NAND3_X1  g437(.A1(new_n549), .A2(G55), .A3(new_n550), .ZN(new_n863));
  NAND2_X1  g438(.A1(G80), .A2(G543), .ZN(new_n864));
  INV_X1    g439(.A(G67), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n864), .B1(new_n536), .B2(new_n865), .ZN(new_n866));
  AOI22_X1  g441(.A1(new_n556), .A2(G93), .B1(new_n866), .B2(new_n528), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n863), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n569), .A2(new_n571), .A3(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT99), .ZN(new_n870));
  AND2_X1   g445(.A1(new_n863), .A2(new_n867), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(new_n568), .ZN(new_n872));
  AND3_X1   g447(.A1(new_n869), .A2(new_n870), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n870), .B1(new_n869), .B2(new_n872), .ZN(new_n874));
  OR3_X1    g449(.A1(new_n873), .A2(new_n874), .A3(KEYINPUT38), .ZN(new_n875));
  AND2_X1   g450(.A1(new_n629), .A2(G559), .ZN(new_n876));
  OAI21_X1  g451(.A(KEYINPUT38), .B1(new_n873), .B2(new_n874), .ZN(new_n877));
  AND3_X1   g452(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n876), .B1(new_n875), .B2(new_n877), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT39), .ZN(new_n880));
  OR3_X1    g455(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(KEYINPUT100), .ZN(new_n882));
  OR2_X1    g457(.A1(new_n878), .A2(new_n879), .ZN(new_n883));
  AOI21_X1  g458(.A(G860), .B1(new_n883), .B2(new_n880), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n868), .A2(G860), .ZN(new_n886));
  XOR2_X1   g461(.A(new_n886), .B(KEYINPUT37), .Z(new_n887));
  NAND2_X1  g462(.A1(new_n885), .A2(new_n887), .ZN(G145));
  XOR2_X1   g463(.A(G160), .B(new_n656), .Z(new_n889));
  XNOR2_X1  g464(.A(new_n492), .B(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n746), .B(G164), .ZN(new_n891));
  INV_X1    g466(.A(new_n766), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n746), .B(new_n510), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(new_n766), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n824), .B(KEYINPUT102), .ZN(new_n897));
  OR2_X1    g472(.A1(new_n897), .A2(new_n647), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n647), .ZN(new_n899));
  AND2_X1   g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n896), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n898), .A2(new_n899), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n902), .A2(new_n893), .A3(new_n895), .ZN(new_n903));
  AOI22_X1  g478(.A1(G130), .A2(new_n485), .B1(new_n468), .B2(G142), .ZN(new_n904));
  OAI21_X1  g479(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT101), .ZN(new_n906));
  INV_X1    g481(.A(G118), .ZN(new_n907));
  AOI22_X1  g482(.A1(new_n905), .A2(new_n906), .B1(new_n907), .B2(G2105), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n908), .B1(new_n906), .B2(new_n905), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n904), .A2(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n778), .B(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n901), .A2(new_n903), .A3(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n911), .B1(new_n901), .B2(new_n903), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n890), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n901), .A2(new_n903), .ZN(new_n916));
  INV_X1    g491(.A(new_n911), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n890), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n918), .A2(new_n919), .A3(new_n912), .ZN(new_n920));
  INV_X1    g495(.A(G37), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n915), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n922), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g498(.A(KEYINPUT107), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT42), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT105), .ZN(new_n926));
  NAND2_X1  g501(.A1(G290), .A2(G288), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  NOR2_X1   g503(.A1(G290), .A2(G288), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n926), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n810), .A2(new_n841), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n931), .A2(KEYINPUT105), .A3(new_n927), .ZN(new_n932));
  XNOR2_X1  g507(.A(G303), .B(new_n831), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n930), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT106), .ZN(new_n935));
  INV_X1    g510(.A(new_n933), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n936), .A2(KEYINPUT105), .A3(new_n927), .A4(new_n931), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n934), .A2(new_n935), .A3(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n935), .B1(new_n934), .B2(new_n937), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n925), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n940), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n942), .A2(KEYINPUT42), .A3(new_n938), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n924), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n563), .A2(new_n570), .A3(new_n567), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n570), .B1(new_n563), .B2(new_n567), .ZN(new_n946));
  NOR3_X1   g521(.A1(new_n945), .A2(new_n871), .A3(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(new_n872), .ZN(new_n948));
  OAI21_X1  g523(.A(KEYINPUT99), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n869), .A2(new_n870), .A3(new_n872), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n639), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(G299), .A2(KEYINPUT103), .ZN(new_n952));
  AND2_X1   g527(.A1(new_n591), .A2(new_n592), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT103), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n953), .A2(new_n954), .A3(new_n587), .A4(new_n585), .ZN(new_n955));
  AOI22_X1  g530(.A1(new_n620), .A2(new_n621), .B1(G651), .B2(new_n626), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n952), .A2(new_n623), .A3(new_n955), .A4(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n628), .A2(KEYINPUT103), .A3(G299), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT41), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n957), .A2(new_n958), .A3(KEYINPUT41), .ZN(new_n962));
  AND2_X1   g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n638), .B1(new_n874), .B2(new_n873), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n951), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT104), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n951), .A2(KEYINPUT104), .A3(new_n963), .A4(new_n964), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n951), .A2(new_n964), .ZN(new_n969));
  INV_X1    g544(.A(new_n959), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n967), .A2(new_n968), .A3(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n941), .A2(new_n943), .A3(new_n924), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n944), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  AND2_X1   g550(.A1(new_n941), .A2(new_n943), .ZN(new_n976));
  NOR3_X1   g551(.A1(new_n976), .A2(new_n972), .A3(new_n924), .ZN(new_n977));
  OAI21_X1  g552(.A(G868), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n868), .A2(new_n615), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(G295));
  NAND2_X1  g555(.A1(new_n978), .A2(new_n979), .ZN(G331));
  INV_X1    g556(.A(KEYINPUT44), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n934), .A2(new_n937), .ZN(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  XNOR2_X1  g559(.A(G286), .B(G301), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n985), .B1(new_n873), .B2(new_n874), .ZN(new_n986));
  XNOR2_X1  g561(.A(G286), .B(G171), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n949), .A2(new_n950), .A3(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n986), .A2(new_n988), .A3(new_n970), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT108), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n986), .A2(new_n988), .ZN(new_n991));
  AOI22_X1  g566(.A1(new_n989), .A2(new_n990), .B1(new_n991), .B2(new_n963), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n986), .A2(new_n988), .A3(new_n970), .A4(KEYINPUT108), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n984), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NOR3_X1   g569(.A1(new_n873), .A2(new_n874), .A3(new_n985), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n987), .B1(new_n949), .B2(new_n950), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n963), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n997), .A2(new_n984), .A3(new_n989), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(new_n921), .ZN(new_n999));
  NOR3_X1   g574(.A1(new_n994), .A2(new_n999), .A3(KEYINPUT43), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT43), .ZN(new_n1001));
  AND2_X1   g576(.A1(new_n998), .A2(new_n921), .ZN(new_n1002));
  AND3_X1   g577(.A1(new_n986), .A2(new_n988), .A3(new_n970), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n961), .A2(new_n962), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1004), .B1(new_n986), .B2(new_n988), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n983), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1001), .B1(new_n1002), .B2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n982), .B1(new_n1000), .B2(new_n1007), .ZN(new_n1008));
  OAI211_X1 g583(.A(KEYINPUT110), .B(KEYINPUT43), .C1(new_n994), .C2(new_n999), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n1006), .A2(new_n998), .A3(new_n1001), .A4(new_n921), .ZN(new_n1010));
  AND2_X1   g585(.A1(new_n1010), .A2(KEYINPUT109), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1010), .A2(KEYINPUT109), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1009), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n989), .A2(new_n990), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1014), .A2(new_n997), .A3(new_n993), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(new_n983), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1001), .B1(new_n1002), .B2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(KEYINPUT44), .B1(new_n1017), .B2(KEYINPUT110), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1008), .B1(new_n1013), .B2(new_n1018), .ZN(G397));
  INV_X1    g594(.A(G1384), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n510), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(KEYINPUT116), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT50), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT116), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n510), .A2(new_n1024), .A3(new_n1020), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1022), .A2(new_n1023), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(G2084), .ZN(new_n1027));
  INV_X1    g602(.A(G125), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1028), .B1(new_n466), .B2(new_n467), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n477), .A2(new_n478), .ZN(new_n1030));
  OAI21_X1  g605(.A(G2105), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1031), .A2(G40), .A3(new_n473), .A4(new_n469), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1032), .B1(new_n1021), .B2(KEYINPUT50), .ZN(new_n1033));
  AND3_X1   g608(.A1(new_n1026), .A2(new_n1027), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT45), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n507), .B1(KEYINPUT75), .B2(new_n503), .ZN(new_n1036));
  AOI22_X1  g611(.A1(new_n1036), .A2(new_n506), .B1(new_n497), .B2(new_n500), .ZN(new_n1037));
  AOI211_X1 g612(.A(KEYINPUT116), .B(G1384), .C1(new_n1037), .C2(new_n496), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1024), .B1(new_n510), .B2(new_n1020), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1035), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(G1384), .B1(new_n1037), .B2(new_n496), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1032), .B1(new_n1041), .B2(KEYINPUT45), .ZN(new_n1042));
  AOI21_X1  g617(.A(G1966), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1043));
  OAI211_X1 g618(.A(KEYINPUT124), .B(G8), .C1(new_n1034), .C2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(G8), .ZN(new_n1045));
  NOR2_X1   g620(.A1(G168), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1044), .A2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(KEYINPUT45), .B1(new_n1022), .B2(new_n1025), .ZN(new_n1049));
  OAI211_X1 g624(.A(G40), .B(G160), .C1(new_n1021), .C2(new_n1035), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n749), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1026), .A2(new_n1027), .A3(new_n1033), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1045), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  AND2_X1   g628(.A1(KEYINPUT124), .A2(KEYINPUT51), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1048), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT51), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1057), .B(G8), .C1(new_n1058), .C2(G286), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1046), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NOR3_X1   g636(.A1(new_n1056), .A2(new_n1061), .A3(KEYINPUT125), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT125), .ZN(new_n1063));
  OAI21_X1  g638(.A(G8), .B1(new_n1034), .B2(new_n1043), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(new_n1047), .ZN(new_n1065));
  AOI22_X1  g640(.A1(new_n1065), .A2(new_n1057), .B1(new_n1058), .B2(new_n1046), .ZN(new_n1066));
  OAI211_X1 g641(.A(new_n1044), .B(new_n1047), .C1(new_n1053), .C2(new_n1054), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1063), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(KEYINPUT62), .B1(new_n1062), .B2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(KEYINPUT125), .B1(new_n1056), .B2(new_n1061), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1066), .A2(new_n1063), .A3(new_n1067), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT62), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1070), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(G303), .A2(G8), .ZN(new_n1074));
  XNOR2_X1  g649(.A(new_n1074), .B(KEYINPUT55), .ZN(new_n1075));
  XOR2_X1   g650(.A(KEYINPUT114), .B(G1971), .Z(new_n1076));
  NAND2_X1  g651(.A1(new_n1021), .A2(new_n1035), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1076), .B1(new_n1042), .B2(new_n1077), .ZN(new_n1078));
  OAI211_X1 g653(.A(G160), .B(G40), .C1(new_n1021), .C2(KEYINPUT50), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1022), .A2(new_n1025), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1079), .B1(new_n1080), .B2(KEYINPUT50), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1078), .B1(new_n1081), .B2(new_n726), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1075), .B1(new_n1082), .B2(new_n1045), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT55), .ZN(new_n1084));
  XNOR2_X1  g659(.A(new_n1074), .B(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1026), .A2(new_n726), .A3(new_n1033), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT115), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1076), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1041), .A2(KEYINPUT45), .ZN(new_n1089));
  OAI211_X1 g664(.A(new_n1087), .B(new_n1088), .C1(new_n1050), .C2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1086), .A2(new_n1090), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1078), .A2(new_n1087), .ZN(new_n1092));
  OAI211_X1 g667(.A(G8), .B(new_n1085), .C1(new_n1091), .C2(new_n1092), .ZN(new_n1093));
  AND2_X1   g668(.A1(new_n1083), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT49), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n719), .B1(new_n604), .B2(KEYINPUT117), .ZN(new_n1096));
  AND2_X1   g671(.A1(G305), .A2(new_n1096), .ZN(new_n1097));
  NOR2_X1   g672(.A1(G305), .A2(new_n1096), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1095), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n604), .A2(KEYINPUT117), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(G1981), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1101), .A2(new_n598), .A3(new_n600), .A4(new_n604), .ZN(new_n1102));
  NAND2_X1  g677(.A1(G305), .A2(new_n1096), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1102), .A2(KEYINPUT49), .A3(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1032), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1022), .A2(new_n1105), .A3(new_n1025), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1099), .A2(new_n1104), .A3(G8), .A4(new_n1106), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n594), .A2(G1976), .A3(new_n595), .A4(new_n596), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1106), .A2(G8), .A3(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(KEYINPUT52), .ZN(new_n1110));
  INV_X1    g685(.A(G1976), .ZN(new_n1111));
  AOI21_X1  g686(.A(KEYINPUT52), .B1(G288), .B2(new_n1111), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1112), .A2(new_n1106), .A3(G8), .A4(new_n1108), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1107), .A2(new_n1110), .A3(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT118), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1107), .A2(new_n1110), .A3(KEYINPUT118), .A4(new_n1113), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1026), .A2(new_n1033), .ZN(new_n1119));
  INV_X1    g694(.A(G1961), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1042), .A2(new_n447), .A3(new_n1077), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT53), .ZN(new_n1122));
  AOI22_X1  g697(.A1(new_n1119), .A2(new_n1120), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1040), .A2(KEYINPUT53), .A3(new_n447), .A4(new_n1042), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  AND4_X1   g700(.A1(G171), .A2(new_n1094), .A3(new_n1118), .A4(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1069), .A2(new_n1073), .A3(new_n1126), .ZN(new_n1127));
  NOR2_X1   g702(.A1(G288), .A2(G1976), .ZN(new_n1128));
  AOI22_X1  g703(.A1(new_n1107), .A2(new_n1128), .B1(new_n719), .B2(new_n831), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1106), .A2(G8), .ZN(new_n1130));
  OAI22_X1  g705(.A1(new_n1093), .A2(new_n1114), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g706(.A(G8), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1132), .A2(new_n1075), .ZN(new_n1133));
  AND4_X1   g708(.A1(KEYINPUT63), .A2(new_n1107), .A3(new_n1113), .A4(new_n1110), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1064), .A2(G286), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1133), .A2(new_n1134), .A3(new_n1135), .A4(new_n1093), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT119), .ZN(new_n1137));
  XNOR2_X1  g712(.A(new_n1136), .B(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1094), .A2(new_n1118), .A3(new_n1135), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT63), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1131), .B1(new_n1138), .B2(new_n1141), .ZN(new_n1142));
  OR2_X1    g717(.A1(new_n1081), .A2(G1956), .ZN(new_n1143));
  NAND2_X1  g718(.A1(G299), .A2(KEYINPUT120), .ZN(new_n1144));
  XNOR2_X1  g719(.A(new_n1144), .B(KEYINPUT57), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1050), .A2(new_n1089), .ZN(new_n1146));
  XNOR2_X1  g721(.A(KEYINPUT121), .B(KEYINPUT56), .ZN(new_n1147));
  XNOR2_X1  g722(.A(new_n1147), .B(G2072), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1143), .A2(new_n1145), .A3(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1145), .B1(new_n1143), .B2(new_n1149), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1106), .A2(G2067), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1152), .B1(new_n806), .B2(new_n1119), .ZN(new_n1153));
  OAI22_X1  g728(.A1(new_n1151), .A2(KEYINPUT122), .B1(new_n628), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT57), .ZN(new_n1155));
  XNOR2_X1  g730(.A(new_n1144), .B(new_n1155), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1081), .A2(G1956), .ZN(new_n1157));
  AND2_X1   g732(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1158));
  OAI211_X1 g733(.A(new_n1156), .B(KEYINPUT122), .C1(new_n1157), .C2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1159), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1150), .B1(new_n1154), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(G1996), .ZN(new_n1162));
  XOR2_X1   g737(.A(KEYINPUT58), .B(G1341), .Z(new_n1163));
  AOI22_X1  g738(.A1(new_n1146), .A2(new_n1162), .B1(new_n1106), .B2(new_n1163), .ZN(new_n1164));
  OR3_X1    g739(.A1(new_n1164), .A2(KEYINPUT59), .A3(new_n572), .ZN(new_n1165));
  OAI21_X1  g740(.A(KEYINPUT59), .B1(new_n1164), .B2(new_n572), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n628), .A2(KEYINPUT60), .ZN(new_n1167));
  AOI22_X1  g742(.A1(new_n1165), .A2(new_n1166), .B1(new_n1153), .B2(new_n1167), .ZN(new_n1168));
  AND2_X1   g743(.A1(new_n1153), .A2(new_n628), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1153), .A2(new_n628), .ZN(new_n1170));
  OAI21_X1  g745(.A(KEYINPUT60), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  NOR3_X1   g746(.A1(new_n1156), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT61), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1168), .A2(new_n1171), .A3(new_n1174), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1156), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1176));
  OR2_X1    g751(.A1(new_n1176), .A2(KEYINPUT123), .ZN(new_n1177));
  AOI21_X1  g752(.A(KEYINPUT61), .B1(new_n1176), .B2(KEYINPUT123), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1172), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1161), .B1(new_n1175), .B2(new_n1179), .ZN(new_n1180));
  XNOR2_X1  g755(.A(G301), .B(KEYINPUT54), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n1122), .A2(G2078), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1181), .B1(new_n1146), .B2(new_n1182), .ZN(new_n1183));
  AOI22_X1  g758(.A1(new_n1125), .A2(new_n1181), .B1(new_n1183), .B2(new_n1123), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1094), .A2(new_n1118), .A3(new_n1184), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n1185), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT126), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1180), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  AOI211_X1 g763(.A(KEYINPUT126), .B(new_n1185), .C1(new_n1070), .C2(new_n1071), .ZN(new_n1189));
  OAI211_X1 g764(.A(new_n1127), .B(new_n1142), .C1(new_n1188), .C2(new_n1189), .ZN(new_n1190));
  NOR2_X1   g765(.A1(new_n1077), .A2(new_n1032), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1191), .A2(new_n1162), .ZN(new_n1192));
  XNOR2_X1  g767(.A(new_n1192), .B(KEYINPUT111), .ZN(new_n1193));
  NOR2_X1   g768(.A1(new_n1193), .A2(new_n778), .ZN(new_n1194));
  XOR2_X1   g769(.A(new_n1191), .B(KEYINPUT112), .Z(new_n1195));
  INV_X1    g770(.A(G2067), .ZN(new_n1196));
  XNOR2_X1  g771(.A(new_n766), .B(new_n1196), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n778), .A2(G1996), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g774(.A(new_n1194), .B1(new_n1195), .B2(new_n1199), .ZN(new_n1200));
  NOR2_X1   g775(.A1(new_n824), .A2(new_n827), .ZN(new_n1201));
  AND2_X1   g776(.A1(new_n824), .A2(new_n827), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n1195), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  AND2_X1   g778(.A1(new_n1200), .A2(new_n1203), .ZN(new_n1204));
  NOR2_X1   g779(.A1(new_n810), .A2(new_n714), .ZN(new_n1205));
  NOR2_X1   g780(.A1(G290), .A2(G1986), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1191), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1204), .A2(new_n1207), .ZN(new_n1208));
  INV_X1    g783(.A(KEYINPUT113), .ZN(new_n1209));
  XNOR2_X1  g784(.A(new_n1208), .B(new_n1209), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1190), .A2(new_n1210), .ZN(new_n1211));
  AND2_X1   g786(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1212));
  NOR2_X1   g787(.A1(new_n766), .A2(G2067), .ZN(new_n1213));
  OAI21_X1  g788(.A(new_n1195), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  INV_X1    g789(.A(new_n1197), .ZN(new_n1215));
  OAI21_X1  g790(.A(new_n1195), .B1(new_n1215), .B2(new_n778), .ZN(new_n1216));
  AND2_X1   g791(.A1(new_n1193), .A2(KEYINPUT46), .ZN(new_n1217));
  NOR2_X1   g792(.A1(new_n1193), .A2(KEYINPUT46), .ZN(new_n1218));
  OAI21_X1  g793(.A(new_n1216), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  XNOR2_X1  g794(.A(new_n1219), .B(KEYINPUT47), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n1206), .A2(new_n1191), .ZN(new_n1221));
  XNOR2_X1  g796(.A(new_n1221), .B(KEYINPUT48), .ZN(new_n1222));
  NAND2_X1  g797(.A1(new_n1204), .A2(new_n1222), .ZN(new_n1223));
  AND3_X1   g798(.A1(new_n1214), .A2(new_n1220), .A3(new_n1223), .ZN(new_n1224));
  NAND2_X1  g799(.A1(new_n1211), .A2(new_n1224), .ZN(G329));
  assign    G231 = 1'b0;
  AND2_X1   g800(.A1(new_n674), .A2(G319), .ZN(new_n1227));
  NAND3_X1  g801(.A1(new_n694), .A2(new_n695), .A3(new_n1227), .ZN(new_n1228));
  OAI21_X1  g802(.A(KEYINPUT127), .B1(G229), .B2(new_n1228), .ZN(new_n1229));
  INV_X1    g803(.A(new_n720), .ZN(new_n1230));
  XNOR2_X1  g804(.A(new_n717), .B(new_n1230), .ZN(new_n1231));
  INV_X1    g805(.A(KEYINPUT127), .ZN(new_n1232));
  NAND4_X1  g806(.A1(new_n1231), .A2(new_n696), .A3(new_n1232), .A4(new_n1227), .ZN(new_n1233));
  NAND2_X1  g807(.A1(new_n1229), .A2(new_n1233), .ZN(new_n1234));
  OAI211_X1 g808(.A(new_n1234), .B(new_n922), .C1(new_n1007), .C2(new_n1000), .ZN(G225));
  INV_X1    g809(.A(G225), .ZN(G308));
endmodule


