

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  BUF_X4 U554 ( .A(n885), .Z(n521) );
  XNOR2_X2 U555 ( .A(n534), .B(KEYINPUT67), .ZN(n885) );
  INV_X2 U556 ( .A(n627), .ZN(n520) );
  NOR2_X1 U557 ( .A1(n538), .A2(n537), .ZN(n539) );
  BUF_X1 U558 ( .A(n710), .Z(n711) );
  INV_X1 U559 ( .A(G2105), .ZN(n533) );
  NOR2_X1 U560 ( .A1(G1384), .A2(n765), .ZN(n732) );
  NOR2_X1 U561 ( .A1(n612), .A2(n611), .ZN(n613) );
  INV_X1 U562 ( .A(n520), .ZN(n675) );
  NOR2_X1 U563 ( .A1(n675), .A2(G2084), .ZN(n669) );
  XOR2_X1 U564 ( .A(KEYINPUT17), .B(n529), .Z(n710) );
  NOR2_X1 U565 ( .A1(G2104), .A2(G2105), .ZN(n529) );
  XNOR2_X1 U566 ( .A(KEYINPUT23), .B(KEYINPUT68), .ZN(n535) );
  NOR2_X1 U567 ( .A1(n748), .A2(n523), .ZN(n749) );
  AND2_X1 U568 ( .A1(n607), .A2(n606), .ZN(n608) );
  AND2_X1 U569 ( .A1(n700), .A2(n527), .ZN(n522) );
  NOR2_X1 U570 ( .A1(n533), .A2(G2104), .ZN(n530) );
  NAND2_X1 U571 ( .A1(n522), .A2(n709), .ZN(n750) );
  XNOR2_X1 U572 ( .A(n685), .B(n684), .ZN(n686) );
  XNOR2_X1 U573 ( .A(n536), .B(n535), .ZN(n537) );
  AND2_X1 U574 ( .A1(n945), .A2(n760), .ZN(n523) );
  AND2_X1 U575 ( .A1(G126), .A2(n716), .ZN(n524) );
  AND2_X1 U576 ( .A1(G114), .A2(n879), .ZN(n525) );
  AND2_X1 U577 ( .A1(n669), .A2(G8), .ZN(n526) );
  OR2_X1 U578 ( .A1(n707), .A2(n699), .ZN(n527) );
  NAND2_X1 U579 ( .A1(n672), .A2(n671), .ZN(n528) );
  INV_X1 U580 ( .A(KEYINPUT26), .ZN(n628) );
  XNOR2_X1 U581 ( .A(n629), .B(n628), .ZN(n631) );
  INV_X1 U582 ( .A(KEYINPUT101), .ZN(n657) );
  XNOR2_X1 U583 ( .A(KEYINPUT29), .B(n653), .ZN(n654) );
  INV_X1 U584 ( .A(KEYINPUT31), .ZN(n665) );
  INV_X1 U585 ( .A(KEYINPUT32), .ZN(n684) );
  NAND2_X1 U586 ( .A1(n528), .A2(n686), .ZN(n701) );
  NOR2_X1 U587 ( .A1(n583), .A2(G651), .ZN(n798) );
  XNOR2_X1 U588 ( .A(n541), .B(KEYINPUT65), .ZN(n602) );
  BUF_X1 U589 ( .A(n602), .Z(G160) );
  AND2_X1 U590 ( .A1(G2105), .A2(G2104), .ZN(n879) );
  NAND2_X1 U591 ( .A1(n879), .A2(G113), .ZN(n540) );
  NAND2_X1 U592 ( .A1(G137), .A2(n710), .ZN(n532) );
  XNOR2_X2 U593 ( .A(n530), .B(KEYINPUT66), .ZN(n716) );
  NAND2_X1 U594 ( .A1(G125), .A2(n716), .ZN(n531) );
  NAND2_X1 U595 ( .A1(n532), .A2(n531), .ZN(n538) );
  NAND2_X1 U596 ( .A1(n533), .A2(G2104), .ZN(n534) );
  NAND2_X1 U597 ( .A1(G101), .A2(n521), .ZN(n536) );
  NAND2_X1 U598 ( .A1(n540), .A2(n539), .ZN(n541) );
  XOR2_X1 U599 ( .A(KEYINPUT0), .B(G543), .Z(n583) );
  NAND2_X1 U600 ( .A1(n798), .A2(G52), .ZN(n545) );
  INV_X1 U601 ( .A(G651), .ZN(n546) );
  NOR2_X1 U602 ( .A1(G543), .A2(n546), .ZN(n542) );
  XOR2_X1 U603 ( .A(KEYINPUT70), .B(n542), .Z(n543) );
  XNOR2_X1 U604 ( .A(KEYINPUT1), .B(n543), .ZN(n791) );
  NAND2_X1 U605 ( .A1(G64), .A2(n791), .ZN(n544) );
  NAND2_X1 U606 ( .A1(n545), .A2(n544), .ZN(n552) );
  NOR2_X1 U607 ( .A1(n583), .A2(n546), .ZN(n794) );
  NAND2_X1 U608 ( .A1(n794), .A2(G77), .ZN(n549) );
  NOR2_X1 U609 ( .A1(G651), .A2(G543), .ZN(n547) );
  XNOR2_X1 U610 ( .A(n547), .B(KEYINPUT64), .ZN(n790) );
  NAND2_X1 U611 ( .A1(G90), .A2(n790), .ZN(n548) );
  NAND2_X1 U612 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U613 ( .A(KEYINPUT9), .B(n550), .Z(n551) );
  NOR2_X1 U614 ( .A1(n552), .A2(n551), .ZN(G171) );
  NAND2_X1 U615 ( .A1(G91), .A2(n790), .ZN(n554) );
  NAND2_X1 U616 ( .A1(G65), .A2(n791), .ZN(n553) );
  NAND2_X1 U617 ( .A1(n554), .A2(n553), .ZN(n557) );
  NAND2_X1 U618 ( .A1(G53), .A2(n798), .ZN(n555) );
  XNOR2_X1 U619 ( .A(KEYINPUT71), .B(n555), .ZN(n556) );
  NOR2_X1 U620 ( .A1(n557), .A2(n556), .ZN(n559) );
  NAND2_X1 U621 ( .A1(n794), .A2(G78), .ZN(n558) );
  NAND2_X1 U622 ( .A1(n559), .A2(n558), .ZN(G299) );
  NAND2_X1 U623 ( .A1(G89), .A2(n790), .ZN(n560) );
  XNOR2_X1 U624 ( .A(n560), .B(KEYINPUT4), .ZN(n562) );
  NAND2_X1 U625 ( .A1(G76), .A2(n794), .ZN(n561) );
  NAND2_X1 U626 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U627 ( .A(n563), .B(KEYINPUT5), .ZN(n569) );
  XNOR2_X1 U628 ( .A(KEYINPUT6), .B(KEYINPUT75), .ZN(n567) );
  NAND2_X1 U629 ( .A1(n798), .A2(G51), .ZN(n565) );
  NAND2_X1 U630 ( .A1(G63), .A2(n791), .ZN(n564) );
  NAND2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(n568) );
  NAND2_X1 U633 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U634 ( .A(KEYINPUT7), .B(n570), .ZN(G168) );
  XOR2_X1 U635 ( .A(G168), .B(KEYINPUT8), .Z(n571) );
  XNOR2_X1 U636 ( .A(KEYINPUT76), .B(n571), .ZN(G286) );
  NAND2_X1 U637 ( .A1(n794), .A2(G75), .ZN(n573) );
  NAND2_X1 U638 ( .A1(G88), .A2(n790), .ZN(n572) );
  NAND2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n577) );
  NAND2_X1 U640 ( .A1(n798), .A2(G50), .ZN(n575) );
  NAND2_X1 U641 ( .A1(G62), .A2(n791), .ZN(n574) );
  NAND2_X1 U642 ( .A1(n575), .A2(n574), .ZN(n576) );
  NOR2_X1 U643 ( .A1(n577), .A2(n576), .ZN(G166) );
  INV_X1 U644 ( .A(G166), .ZN(G303) );
  NAND2_X1 U645 ( .A1(n798), .A2(G49), .ZN(n578) );
  XOR2_X1 U646 ( .A(KEYINPUT81), .B(n578), .Z(n580) );
  NAND2_X1 U647 ( .A1(G651), .A2(G74), .ZN(n579) );
  NAND2_X1 U648 ( .A1(n580), .A2(n579), .ZN(n581) );
  NOR2_X1 U649 ( .A1(n791), .A2(n581), .ZN(n582) );
  XNOR2_X1 U650 ( .A(KEYINPUT82), .B(n582), .ZN(n586) );
  NAND2_X1 U651 ( .A1(n583), .A2(G87), .ZN(n584) );
  XOR2_X1 U652 ( .A(KEYINPUT83), .B(n584), .Z(n585) );
  NAND2_X1 U653 ( .A1(n586), .A2(n585), .ZN(G288) );
  NAND2_X1 U654 ( .A1(G86), .A2(n790), .ZN(n588) );
  NAND2_X1 U655 ( .A1(G61), .A2(n791), .ZN(n587) );
  NAND2_X1 U656 ( .A1(n588), .A2(n587), .ZN(n591) );
  NAND2_X1 U657 ( .A1(n794), .A2(G73), .ZN(n589) );
  XOR2_X1 U658 ( .A(KEYINPUT2), .B(n589), .Z(n590) );
  NOR2_X1 U659 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U660 ( .A(n592), .B(KEYINPUT84), .ZN(n594) );
  NAND2_X1 U661 ( .A1(G48), .A2(n798), .ZN(n593) );
  NAND2_X1 U662 ( .A1(n594), .A2(n593), .ZN(G305) );
  NAND2_X1 U663 ( .A1(n794), .A2(G72), .ZN(n596) );
  NAND2_X1 U664 ( .A1(G85), .A2(n790), .ZN(n595) );
  NAND2_X1 U665 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X1 U666 ( .A(KEYINPUT69), .B(n597), .ZN(n601) );
  NAND2_X1 U667 ( .A1(n791), .A2(G60), .ZN(n599) );
  NAND2_X1 U668 ( .A1(n798), .A2(G47), .ZN(n598) );
  AND2_X1 U669 ( .A1(n599), .A2(n598), .ZN(n600) );
  NAND2_X1 U670 ( .A1(n601), .A2(n600), .ZN(G290) );
  NAND2_X1 U671 ( .A1(n602), .A2(G40), .ZN(n731) );
  INV_X1 U672 ( .A(n731), .ZN(n609) );
  NAND2_X1 U673 ( .A1(G138), .A2(n710), .ZN(n604) );
  NAND2_X1 U674 ( .A1(G102), .A2(n521), .ZN(n603) );
  NAND2_X1 U675 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X1 U676 ( .A(n605), .B(KEYINPUT89), .ZN(n607) );
  NOR2_X1 U677 ( .A1(n524), .A2(n525), .ZN(n606) );
  XNOR2_X1 U678 ( .A(KEYINPUT90), .B(n608), .ZN(n765) );
  NAND2_X1 U679 ( .A1(n609), .A2(n732), .ZN(n627) );
  NAND2_X1 U680 ( .A1(G8), .A2(n627), .ZN(n707) );
  XNOR2_X1 U681 ( .A(KEYINPUT25), .B(G2078), .ZN(n971) );
  NAND2_X1 U682 ( .A1(n520), .A2(n971), .ZN(n610) );
  XNOR2_X1 U683 ( .A(n610), .B(KEYINPUT99), .ZN(n612) );
  NOR2_X1 U684 ( .A1(n520), .A2(G1961), .ZN(n611) );
  XOR2_X1 U685 ( .A(KEYINPUT100), .B(n613), .Z(n662) );
  NAND2_X1 U686 ( .A1(G171), .A2(n662), .ZN(n656) );
  INV_X1 U687 ( .A(G299), .ZN(n947) );
  NAND2_X1 U688 ( .A1(n520), .A2(G2072), .ZN(n614) );
  XNOR2_X1 U689 ( .A(n614), .B(KEYINPUT27), .ZN(n616) );
  INV_X1 U690 ( .A(G1956), .ZN(n920) );
  NOR2_X1 U691 ( .A1(n920), .A2(n520), .ZN(n615) );
  NOR2_X1 U692 ( .A1(n616), .A2(n615), .ZN(n648) );
  NOR2_X1 U693 ( .A1(n947), .A2(n648), .ZN(n617) );
  XOR2_X1 U694 ( .A(n617), .B(KEYINPUT28), .Z(n652) );
  NAND2_X1 U695 ( .A1(n791), .A2(G56), .ZN(n618) );
  XOR2_X1 U696 ( .A(KEYINPUT14), .B(n618), .Z(n624) );
  NAND2_X1 U697 ( .A1(G81), .A2(n790), .ZN(n619) );
  XNOR2_X1 U698 ( .A(n619), .B(KEYINPUT12), .ZN(n621) );
  NAND2_X1 U699 ( .A1(G68), .A2(n794), .ZN(n620) );
  NAND2_X1 U700 ( .A1(n621), .A2(n620), .ZN(n622) );
  XOR2_X1 U701 ( .A(KEYINPUT13), .B(n622), .Z(n623) );
  NOR2_X1 U702 ( .A1(n624), .A2(n623), .ZN(n626) );
  NAND2_X1 U703 ( .A1(n798), .A2(G43), .ZN(n625) );
  NAND2_X1 U704 ( .A1(n626), .A2(n625), .ZN(n965) );
  AND2_X1 U705 ( .A1(n520), .A2(G1996), .ZN(n629) );
  NAND2_X1 U706 ( .A1(n675), .A2(G1341), .ZN(n630) );
  NAND2_X1 U707 ( .A1(n631), .A2(n630), .ZN(n632) );
  NOR2_X1 U708 ( .A1(n965), .A2(n632), .ZN(n644) );
  NAND2_X1 U709 ( .A1(G92), .A2(n790), .ZN(n634) );
  NAND2_X1 U710 ( .A1(G66), .A2(n791), .ZN(n633) );
  NAND2_X1 U711 ( .A1(n634), .A2(n633), .ZN(n639) );
  NAND2_X1 U712 ( .A1(G79), .A2(n794), .ZN(n636) );
  NAND2_X1 U713 ( .A1(G54), .A2(n798), .ZN(n635) );
  NAND2_X1 U714 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U715 ( .A(KEYINPUT74), .B(n637), .ZN(n638) );
  NOR2_X1 U716 ( .A1(n639), .A2(n638), .ZN(n640) );
  XNOR2_X1 U717 ( .A(n640), .B(KEYINPUT15), .ZN(n954) );
  NAND2_X1 U718 ( .A1(G1348), .A2(n675), .ZN(n642) );
  NAND2_X1 U719 ( .A1(n520), .A2(G2067), .ZN(n641) );
  NAND2_X1 U720 ( .A1(n642), .A2(n641), .ZN(n645) );
  NOR2_X1 U721 ( .A1(n954), .A2(n645), .ZN(n643) );
  OR2_X1 U722 ( .A1(n644), .A2(n643), .ZN(n647) );
  NAND2_X1 U723 ( .A1(n954), .A2(n645), .ZN(n646) );
  NAND2_X1 U724 ( .A1(n647), .A2(n646), .ZN(n650) );
  NAND2_X1 U725 ( .A1(n947), .A2(n648), .ZN(n649) );
  NAND2_X1 U726 ( .A1(n650), .A2(n649), .ZN(n651) );
  NAND2_X1 U727 ( .A1(n652), .A2(n651), .ZN(n653) );
  INV_X1 U728 ( .A(n654), .ZN(n655) );
  NAND2_X1 U729 ( .A1(n656), .A2(n655), .ZN(n668) );
  NOR2_X1 U730 ( .A1(G1966), .A2(n707), .ZN(n670) );
  NOR2_X1 U731 ( .A1(n670), .A2(n669), .ZN(n658) );
  XNOR2_X1 U732 ( .A(n658), .B(n657), .ZN(n659) );
  NAND2_X1 U733 ( .A1(n659), .A2(G8), .ZN(n660) );
  XNOR2_X1 U734 ( .A(n660), .B(KEYINPUT30), .ZN(n661) );
  NOR2_X1 U735 ( .A1(n661), .A2(G168), .ZN(n664) );
  NOR2_X1 U736 ( .A1(G171), .A2(n662), .ZN(n663) );
  NOR2_X1 U737 ( .A1(n664), .A2(n663), .ZN(n666) );
  XNOR2_X1 U738 ( .A(n666), .B(n665), .ZN(n667) );
  NAND2_X1 U739 ( .A1(n668), .A2(n667), .ZN(n674) );
  XNOR2_X1 U740 ( .A(n674), .B(KEYINPUT102), .ZN(n672) );
  NOR2_X1 U741 ( .A1(n526), .A2(n670), .ZN(n671) );
  AND2_X1 U742 ( .A1(G286), .A2(G8), .ZN(n673) );
  NAND2_X1 U743 ( .A1(n674), .A2(n673), .ZN(n683) );
  INV_X1 U744 ( .A(G8), .ZN(n681) );
  NOR2_X1 U745 ( .A1(G1971), .A2(n707), .ZN(n677) );
  NOR2_X1 U746 ( .A1(G2090), .A2(n675), .ZN(n676) );
  NOR2_X1 U747 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U748 ( .A1(n678), .A2(G303), .ZN(n679) );
  XOR2_X1 U749 ( .A(KEYINPUT103), .B(n679), .Z(n680) );
  OR2_X1 U750 ( .A1(n681), .A2(n680), .ZN(n682) );
  NAND2_X1 U751 ( .A1(n683), .A2(n682), .ZN(n685) );
  NOR2_X1 U752 ( .A1(G1976), .A2(G288), .ZN(n951) );
  NOR2_X1 U753 ( .A1(G1971), .A2(G303), .ZN(n687) );
  NOR2_X1 U754 ( .A1(n951), .A2(n687), .ZN(n688) );
  NAND2_X1 U755 ( .A1(n701), .A2(n688), .ZN(n689) );
  NAND2_X1 U756 ( .A1(G1976), .A2(G288), .ZN(n957) );
  NAND2_X1 U757 ( .A1(n689), .A2(n957), .ZN(n690) );
  XNOR2_X1 U758 ( .A(n690), .B(KEYINPUT104), .ZN(n691) );
  NOR2_X1 U759 ( .A1(n707), .A2(n691), .ZN(n692) );
  NOR2_X1 U760 ( .A1(KEYINPUT33), .A2(n692), .ZN(n693) );
  XNOR2_X1 U761 ( .A(n693), .B(KEYINPUT105), .ZN(n694) );
  XOR2_X1 U762 ( .A(G1981), .B(G305), .Z(n960) );
  NAND2_X1 U763 ( .A1(n694), .A2(n960), .ZN(n706) );
  INV_X1 U764 ( .A(n706), .ZN(n696) );
  NAND2_X1 U765 ( .A1(KEYINPUT33), .A2(n951), .ZN(n695) );
  NAND2_X1 U766 ( .A1(n696), .A2(n695), .ZN(n700) );
  NOR2_X1 U767 ( .A1(G1981), .A2(G305), .ZN(n697) );
  XOR2_X1 U768 ( .A(n697), .B(KEYINPUT24), .Z(n698) );
  XNOR2_X1 U769 ( .A(KEYINPUT98), .B(n698), .ZN(n699) );
  INV_X1 U770 ( .A(n701), .ZN(n704) );
  NAND2_X1 U771 ( .A1(G166), .A2(G8), .ZN(n702) );
  NOR2_X1 U772 ( .A1(G2090), .A2(n702), .ZN(n703) );
  NOR2_X1 U773 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U774 ( .A1(n706), .A2(n705), .ZN(n708) );
  NAND2_X1 U775 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U776 ( .A1(n711), .A2(G131), .ZN(n712) );
  XOR2_X1 U777 ( .A(KEYINPUT95), .B(n712), .Z(n714) );
  NAND2_X1 U778 ( .A1(n521), .A2(G95), .ZN(n713) );
  NAND2_X1 U779 ( .A1(n714), .A2(n713), .ZN(n715) );
  XOR2_X1 U780 ( .A(KEYINPUT96), .B(n715), .Z(n720) );
  NAND2_X1 U781 ( .A1(n716), .A2(G119), .ZN(n718) );
  NAND2_X1 U782 ( .A1(G107), .A2(n879), .ZN(n717) );
  AND2_X1 U783 ( .A1(n718), .A2(n717), .ZN(n719) );
  NAND2_X1 U784 ( .A1(n720), .A2(n719), .ZN(n870) );
  AND2_X1 U785 ( .A1(n870), .A2(G1991), .ZN(n730) );
  NAND2_X1 U786 ( .A1(G141), .A2(n711), .ZN(n722) );
  NAND2_X1 U787 ( .A1(G117), .A2(n879), .ZN(n721) );
  NAND2_X1 U788 ( .A1(n722), .A2(n721), .ZN(n726) );
  NAND2_X1 U789 ( .A1(G105), .A2(n521), .ZN(n723) );
  XNOR2_X1 U790 ( .A(n723), .B(KEYINPUT38), .ZN(n724) );
  XNOR2_X1 U791 ( .A(n724), .B(KEYINPUT97), .ZN(n725) );
  NOR2_X1 U792 ( .A1(n726), .A2(n725), .ZN(n728) );
  NAND2_X1 U793 ( .A1(G129), .A2(n716), .ZN(n727) );
  NAND2_X1 U794 ( .A1(n728), .A2(n727), .ZN(n892) );
  AND2_X1 U795 ( .A1(n892), .A2(G1996), .ZN(n729) );
  NOR2_X1 U796 ( .A1(n730), .A2(n729), .ZN(n1007) );
  NOR2_X1 U797 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U798 ( .A(KEYINPUT91), .B(n733), .ZN(n734) );
  NOR2_X1 U799 ( .A1(n1007), .A2(n734), .ZN(n753) );
  INV_X1 U800 ( .A(n753), .ZN(n747) );
  INV_X1 U801 ( .A(n734), .ZN(n760) );
  XNOR2_X1 U802 ( .A(G2067), .B(KEYINPUT37), .ZN(n758) );
  NAND2_X1 U803 ( .A1(G116), .A2(n879), .ZN(n736) );
  NAND2_X1 U804 ( .A1(G128), .A2(n716), .ZN(n735) );
  NAND2_X1 U805 ( .A1(n736), .A2(n735), .ZN(n738) );
  XOR2_X1 U806 ( .A(KEYINPUT35), .B(KEYINPUT94), .Z(n737) );
  XNOR2_X1 U807 ( .A(n738), .B(n737), .ZN(n745) );
  NAND2_X1 U808 ( .A1(n521), .A2(G104), .ZN(n739) );
  XNOR2_X1 U809 ( .A(n739), .B(KEYINPUT92), .ZN(n741) );
  NAND2_X1 U810 ( .A1(G140), .A2(n711), .ZN(n740) );
  NAND2_X1 U811 ( .A1(n741), .A2(n740), .ZN(n742) );
  XOR2_X1 U812 ( .A(n742), .B(KEYINPUT34), .Z(n743) );
  XNOR2_X1 U813 ( .A(KEYINPUT93), .B(n743), .ZN(n744) );
  NOR2_X1 U814 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U815 ( .A(KEYINPUT36), .B(n746), .ZN(n895) );
  NOR2_X1 U816 ( .A1(n758), .A2(n895), .ZN(n993) );
  NAND2_X1 U817 ( .A1(n760), .A2(n993), .ZN(n756) );
  NAND2_X1 U818 ( .A1(n747), .A2(n756), .ZN(n748) );
  XNOR2_X1 U819 ( .A(G1986), .B(G290), .ZN(n945) );
  NAND2_X1 U820 ( .A1(n750), .A2(n749), .ZN(n763) );
  NOR2_X1 U821 ( .A1(G1996), .A2(n892), .ZN(n1004) );
  NOR2_X1 U822 ( .A1(G1986), .A2(G290), .ZN(n751) );
  NOR2_X1 U823 ( .A1(G1991), .A2(n870), .ZN(n998) );
  NOR2_X1 U824 ( .A1(n751), .A2(n998), .ZN(n752) );
  NOR2_X1 U825 ( .A1(n753), .A2(n752), .ZN(n754) );
  NOR2_X1 U826 ( .A1(n1004), .A2(n754), .ZN(n755) );
  XNOR2_X1 U827 ( .A(KEYINPUT39), .B(n755), .ZN(n757) );
  NAND2_X1 U828 ( .A1(n757), .A2(n756), .ZN(n759) );
  NAND2_X1 U829 ( .A1(n758), .A2(n895), .ZN(n994) );
  NAND2_X1 U830 ( .A1(n759), .A2(n994), .ZN(n761) );
  NAND2_X1 U831 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U832 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U833 ( .A(n764), .B(KEYINPUT40), .ZN(G329) );
  BUF_X1 U834 ( .A(n765), .Z(G164) );
  AND2_X1 U835 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U836 ( .A(G57), .ZN(G237) );
  INV_X1 U837 ( .A(G132), .ZN(G219) );
  NAND2_X1 U838 ( .A1(G7), .A2(G661), .ZN(n766) );
  XNOR2_X1 U839 ( .A(n766), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U840 ( .A(G223), .ZN(n830) );
  NAND2_X1 U841 ( .A1(n830), .A2(G567), .ZN(n767) );
  XOR2_X1 U842 ( .A(KEYINPUT11), .B(n767), .Z(G234) );
  XNOR2_X1 U843 ( .A(G860), .B(KEYINPUT73), .ZN(n772) );
  OR2_X1 U844 ( .A1(n965), .A2(n772), .ZN(G153) );
  INV_X1 U845 ( .A(G171), .ZN(G301) );
  NAND2_X1 U846 ( .A1(G868), .A2(G301), .ZN(n769) );
  INV_X1 U847 ( .A(G868), .ZN(n811) );
  NAND2_X1 U848 ( .A1(n954), .A2(n811), .ZN(n768) );
  NAND2_X1 U849 ( .A1(n769), .A2(n768), .ZN(G284) );
  NAND2_X1 U850 ( .A1(G868), .A2(G286), .ZN(n771) );
  NAND2_X1 U851 ( .A1(G299), .A2(n811), .ZN(n770) );
  NAND2_X1 U852 ( .A1(n771), .A2(n770), .ZN(G297) );
  NAND2_X1 U853 ( .A1(G559), .A2(n772), .ZN(n773) );
  XOR2_X1 U854 ( .A(KEYINPUT77), .B(n773), .Z(n774) );
  INV_X1 U855 ( .A(n954), .ZN(n898) );
  NAND2_X1 U856 ( .A1(n774), .A2(n898), .ZN(n775) );
  XNOR2_X1 U857 ( .A(n775), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U858 ( .A1(G868), .A2(n965), .ZN(n778) );
  NAND2_X1 U859 ( .A1(G868), .A2(n898), .ZN(n776) );
  NOR2_X1 U860 ( .A1(G559), .A2(n776), .ZN(n777) );
  NOR2_X1 U861 ( .A1(n778), .A2(n777), .ZN(G282) );
  XOR2_X1 U862 ( .A(KEYINPUT18), .B(KEYINPUT78), .Z(n780) );
  NAND2_X1 U863 ( .A1(G123), .A2(n716), .ZN(n779) );
  XNOR2_X1 U864 ( .A(n780), .B(n779), .ZN(n784) );
  NAND2_X1 U865 ( .A1(G135), .A2(n711), .ZN(n782) );
  NAND2_X1 U866 ( .A1(G111), .A2(n879), .ZN(n781) );
  NAND2_X1 U867 ( .A1(n782), .A2(n781), .ZN(n783) );
  NOR2_X1 U868 ( .A1(n784), .A2(n783), .ZN(n786) );
  NAND2_X1 U869 ( .A1(n521), .A2(G99), .ZN(n785) );
  NAND2_X1 U870 ( .A1(n786), .A2(n785), .ZN(n996) );
  XOR2_X1 U871 ( .A(n996), .B(G2096), .Z(n788) );
  XNOR2_X1 U872 ( .A(G2100), .B(KEYINPUT79), .ZN(n787) );
  NAND2_X1 U873 ( .A1(n788), .A2(n787), .ZN(G156) );
  NAND2_X1 U874 ( .A1(n898), .A2(G559), .ZN(n808) );
  XNOR2_X1 U875 ( .A(n965), .B(n808), .ZN(n789) );
  NOR2_X1 U876 ( .A1(n789), .A2(G860), .ZN(n801) );
  NAND2_X1 U877 ( .A1(G93), .A2(n790), .ZN(n793) );
  NAND2_X1 U878 ( .A1(G67), .A2(n791), .ZN(n792) );
  NAND2_X1 U879 ( .A1(n793), .A2(n792), .ZN(n797) );
  NAND2_X1 U880 ( .A1(n794), .A2(G80), .ZN(n795) );
  XOR2_X1 U881 ( .A(KEYINPUT80), .B(n795), .Z(n796) );
  NOR2_X1 U882 ( .A1(n797), .A2(n796), .ZN(n800) );
  NAND2_X1 U883 ( .A1(n798), .A2(G55), .ZN(n799) );
  NAND2_X1 U884 ( .A1(n800), .A2(n799), .ZN(n810) );
  XOR2_X1 U885 ( .A(n801), .B(n810), .Z(G145) );
  XNOR2_X1 U886 ( .A(KEYINPUT19), .B(G303), .ZN(n802) );
  XNOR2_X1 U887 ( .A(n802), .B(G290), .ZN(n805) );
  XNOR2_X1 U888 ( .A(n947), .B(G288), .ZN(n803) );
  XNOR2_X1 U889 ( .A(n803), .B(n810), .ZN(n804) );
  XNOR2_X1 U890 ( .A(n805), .B(n804), .ZN(n806) );
  XNOR2_X1 U891 ( .A(n806), .B(G305), .ZN(n807) );
  XNOR2_X1 U892 ( .A(n965), .B(n807), .ZN(n899) );
  XOR2_X1 U893 ( .A(n899), .B(n808), .Z(n809) );
  NOR2_X1 U894 ( .A1(n811), .A2(n809), .ZN(n813) );
  AND2_X1 U895 ( .A1(n811), .A2(n810), .ZN(n812) );
  NOR2_X1 U896 ( .A1(n813), .A2(n812), .ZN(n814) );
  XNOR2_X1 U897 ( .A(KEYINPUT85), .B(n814), .ZN(G295) );
  NAND2_X1 U898 ( .A1(G2084), .A2(G2078), .ZN(n816) );
  XOR2_X1 U899 ( .A(KEYINPUT20), .B(KEYINPUT86), .Z(n815) );
  XNOR2_X1 U900 ( .A(n816), .B(n815), .ZN(n817) );
  NAND2_X1 U901 ( .A1(G2090), .A2(n817), .ZN(n818) );
  XNOR2_X1 U902 ( .A(KEYINPUT21), .B(n818), .ZN(n819) );
  NAND2_X1 U903 ( .A1(n819), .A2(G2072), .ZN(G158) );
  XOR2_X1 U904 ( .A(KEYINPUT72), .B(G82), .Z(G220) );
  XNOR2_X1 U905 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U906 ( .A1(G220), .A2(G219), .ZN(n821) );
  XNOR2_X1 U907 ( .A(KEYINPUT22), .B(KEYINPUT87), .ZN(n820) );
  XNOR2_X1 U908 ( .A(n821), .B(n820), .ZN(n822) );
  NOR2_X1 U909 ( .A1(n822), .A2(G218), .ZN(n823) );
  NAND2_X1 U910 ( .A1(G96), .A2(n823), .ZN(n836) );
  NAND2_X1 U911 ( .A1(n836), .A2(G2106), .ZN(n827) );
  NAND2_X1 U912 ( .A1(G120), .A2(G108), .ZN(n824) );
  NOR2_X1 U913 ( .A1(G237), .A2(n824), .ZN(n825) );
  NAND2_X1 U914 ( .A1(G69), .A2(n825), .ZN(n837) );
  NAND2_X1 U915 ( .A1(n837), .A2(G567), .ZN(n826) );
  NAND2_X1 U916 ( .A1(n827), .A2(n826), .ZN(n838) );
  NAND2_X1 U917 ( .A1(G661), .A2(G483), .ZN(n828) );
  XNOR2_X1 U918 ( .A(KEYINPUT88), .B(n828), .ZN(n829) );
  NOR2_X1 U919 ( .A1(n838), .A2(n829), .ZN(n834) );
  NAND2_X1 U920 ( .A1(n834), .A2(G36), .ZN(G176) );
  NAND2_X1 U921 ( .A1(G2106), .A2(n830), .ZN(G217) );
  NAND2_X1 U922 ( .A1(G15), .A2(G2), .ZN(n831) );
  XOR2_X1 U923 ( .A(KEYINPUT108), .B(n831), .Z(n832) );
  NAND2_X1 U924 ( .A1(G661), .A2(n832), .ZN(G259) );
  NAND2_X1 U925 ( .A1(G3), .A2(G1), .ZN(n833) );
  NAND2_X1 U926 ( .A1(n834), .A2(n833), .ZN(n835) );
  XOR2_X1 U927 ( .A(KEYINPUT109), .B(n835), .Z(G188) );
  XNOR2_X1 U928 ( .A(G108), .B(KEYINPUT115), .ZN(G238) );
  INV_X1 U930 ( .A(G120), .ZN(G236) );
  INV_X1 U931 ( .A(G96), .ZN(G221) );
  NOR2_X1 U932 ( .A1(n837), .A2(n836), .ZN(G325) );
  INV_X1 U933 ( .A(G325), .ZN(G261) );
  INV_X1 U934 ( .A(n838), .ZN(G319) );
  XOR2_X1 U935 ( .A(G2100), .B(G2096), .Z(n840) );
  XNOR2_X1 U936 ( .A(KEYINPUT42), .B(G2678), .ZN(n839) );
  XNOR2_X1 U937 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U938 ( .A(KEYINPUT43), .B(G2090), .Z(n842) );
  XNOR2_X1 U939 ( .A(G2067), .B(G2072), .ZN(n841) );
  XNOR2_X1 U940 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U941 ( .A(n844), .B(n843), .Z(n846) );
  XNOR2_X1 U942 ( .A(G2084), .B(G2078), .ZN(n845) );
  XNOR2_X1 U943 ( .A(n846), .B(n845), .ZN(G227) );
  XOR2_X1 U944 ( .A(G1986), .B(G1976), .Z(n848) );
  XNOR2_X1 U945 ( .A(G1961), .B(G1956), .ZN(n847) );
  XNOR2_X1 U946 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U947 ( .A(n849), .B(G2474), .Z(n851) );
  XNOR2_X1 U948 ( .A(G1996), .B(G1991), .ZN(n850) );
  XNOR2_X1 U949 ( .A(n851), .B(n850), .ZN(n855) );
  XOR2_X1 U950 ( .A(KEYINPUT41), .B(G1981), .Z(n853) );
  XNOR2_X1 U951 ( .A(G1966), .B(G1971), .ZN(n852) );
  XNOR2_X1 U952 ( .A(n853), .B(n852), .ZN(n854) );
  XNOR2_X1 U953 ( .A(n855), .B(n854), .ZN(G229) );
  NAND2_X1 U954 ( .A1(n716), .A2(G124), .ZN(n856) );
  XNOR2_X1 U955 ( .A(n856), .B(KEYINPUT44), .ZN(n858) );
  NAND2_X1 U956 ( .A1(n879), .A2(G112), .ZN(n857) );
  NAND2_X1 U957 ( .A1(n858), .A2(n857), .ZN(n862) );
  NAND2_X1 U958 ( .A1(G136), .A2(n711), .ZN(n860) );
  NAND2_X1 U959 ( .A1(G100), .A2(n521), .ZN(n859) );
  NAND2_X1 U960 ( .A1(n860), .A2(n859), .ZN(n861) );
  NOR2_X1 U961 ( .A1(n862), .A2(n861), .ZN(G162) );
  NAND2_X1 U962 ( .A1(G118), .A2(n879), .ZN(n864) );
  NAND2_X1 U963 ( .A1(G130), .A2(n716), .ZN(n863) );
  NAND2_X1 U964 ( .A1(n864), .A2(n863), .ZN(n869) );
  NAND2_X1 U965 ( .A1(G142), .A2(n711), .ZN(n866) );
  NAND2_X1 U966 ( .A1(G106), .A2(n521), .ZN(n865) );
  NAND2_X1 U967 ( .A1(n866), .A2(n865), .ZN(n867) );
  XOR2_X1 U968 ( .A(n867), .B(KEYINPUT45), .Z(n868) );
  NOR2_X1 U969 ( .A1(n869), .A2(n868), .ZN(n871) );
  XNOR2_X1 U970 ( .A(n871), .B(n870), .ZN(n878) );
  XOR2_X1 U971 ( .A(KEYINPUT48), .B(KEYINPUT112), .Z(n873) );
  XNOR2_X1 U972 ( .A(KEYINPUT113), .B(KEYINPUT114), .ZN(n872) );
  XNOR2_X1 U973 ( .A(n873), .B(n872), .ZN(n874) );
  XNOR2_X1 U974 ( .A(KEYINPUT46), .B(n874), .ZN(n876) );
  XNOR2_X1 U975 ( .A(n996), .B(KEYINPUT110), .ZN(n875) );
  XNOR2_X1 U976 ( .A(n876), .B(n875), .ZN(n877) );
  XOR2_X1 U977 ( .A(n878), .B(n877), .Z(n890) );
  NAND2_X1 U978 ( .A1(G115), .A2(n879), .ZN(n881) );
  NAND2_X1 U979 ( .A1(G127), .A2(n716), .ZN(n880) );
  NAND2_X1 U980 ( .A1(n881), .A2(n880), .ZN(n882) );
  XNOR2_X1 U981 ( .A(n882), .B(KEYINPUT47), .ZN(n884) );
  NAND2_X1 U982 ( .A1(G139), .A2(n711), .ZN(n883) );
  NAND2_X1 U983 ( .A1(n884), .A2(n883), .ZN(n888) );
  NAND2_X1 U984 ( .A1(G103), .A2(n521), .ZN(n886) );
  XNOR2_X1 U985 ( .A(KEYINPUT111), .B(n886), .ZN(n887) );
  NOR2_X1 U986 ( .A1(n888), .A2(n887), .ZN(n1008) );
  XNOR2_X1 U987 ( .A(G160), .B(n1008), .ZN(n889) );
  XNOR2_X1 U988 ( .A(n890), .B(n889), .ZN(n891) );
  XNOR2_X1 U989 ( .A(G162), .B(n891), .ZN(n894) );
  XOR2_X1 U990 ( .A(G164), .B(n892), .Z(n893) );
  XNOR2_X1 U991 ( .A(n894), .B(n893), .ZN(n896) );
  XOR2_X1 U992 ( .A(n896), .B(n895), .Z(n897) );
  NOR2_X1 U993 ( .A1(G37), .A2(n897), .ZN(G395) );
  XNOR2_X1 U994 ( .A(n898), .B(G286), .ZN(n900) );
  XNOR2_X1 U995 ( .A(n900), .B(n899), .ZN(n901) );
  XNOR2_X1 U996 ( .A(n901), .B(G301), .ZN(n902) );
  NOR2_X1 U997 ( .A1(G37), .A2(n902), .ZN(G397) );
  XNOR2_X1 U998 ( .A(G2451), .B(G2427), .ZN(n912) );
  XOR2_X1 U999 ( .A(G2430), .B(G2443), .Z(n904) );
  XNOR2_X1 U1000 ( .A(KEYINPUT107), .B(G2435), .ZN(n903) );
  XNOR2_X1 U1001 ( .A(n904), .B(n903), .ZN(n908) );
  XOR2_X1 U1002 ( .A(G2438), .B(G2454), .Z(n906) );
  XNOR2_X1 U1003 ( .A(G1341), .B(G1348), .ZN(n905) );
  XNOR2_X1 U1004 ( .A(n906), .B(n905), .ZN(n907) );
  XOR2_X1 U1005 ( .A(n908), .B(n907), .Z(n910) );
  XNOR2_X1 U1006 ( .A(G2446), .B(KEYINPUT106), .ZN(n909) );
  XNOR2_X1 U1007 ( .A(n910), .B(n909), .ZN(n911) );
  XNOR2_X1 U1008 ( .A(n912), .B(n911), .ZN(n913) );
  NAND2_X1 U1009 ( .A1(n913), .A2(G14), .ZN(n919) );
  NAND2_X1 U1010 ( .A1(G319), .A2(n919), .ZN(n916) );
  NOR2_X1 U1011 ( .A1(G227), .A2(G229), .ZN(n914) );
  XNOR2_X1 U1012 ( .A(KEYINPUT49), .B(n914), .ZN(n915) );
  NOR2_X1 U1013 ( .A1(n916), .A2(n915), .ZN(n918) );
  NOR2_X1 U1014 ( .A1(G395), .A2(G397), .ZN(n917) );
  NAND2_X1 U1015 ( .A1(n918), .A2(n917), .ZN(G225) );
  INV_X1 U1016 ( .A(G225), .ZN(G308) );
  INV_X1 U1017 ( .A(G69), .ZN(G235) );
  INV_X1 U1018 ( .A(n919), .ZN(G401) );
  XNOR2_X1 U1019 ( .A(G20), .B(n920), .ZN(n924) );
  XNOR2_X1 U1020 ( .A(G1341), .B(G19), .ZN(n922) );
  XNOR2_X1 U1021 ( .A(G6), .B(G1981), .ZN(n921) );
  NOR2_X1 U1022 ( .A1(n922), .A2(n921), .ZN(n923) );
  NAND2_X1 U1023 ( .A1(n924), .A2(n923), .ZN(n927) );
  XOR2_X1 U1024 ( .A(KEYINPUT59), .B(G1348), .Z(n925) );
  XNOR2_X1 U1025 ( .A(G4), .B(n925), .ZN(n926) );
  NOR2_X1 U1026 ( .A1(n927), .A2(n926), .ZN(n929) );
  XOR2_X1 U1027 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n928) );
  XNOR2_X1 U1028 ( .A(n929), .B(n928), .ZN(n933) );
  XNOR2_X1 U1029 ( .A(G1966), .B(G21), .ZN(n931) );
  XNOR2_X1 U1030 ( .A(G1961), .B(G5), .ZN(n930) );
  NOR2_X1 U1031 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1032 ( .A1(n933), .A2(n932), .ZN(n940) );
  XNOR2_X1 U1033 ( .A(G1971), .B(G22), .ZN(n935) );
  XNOR2_X1 U1034 ( .A(G23), .B(G1976), .ZN(n934) );
  NOR2_X1 U1035 ( .A1(n935), .A2(n934), .ZN(n937) );
  XOR2_X1 U1036 ( .A(G1986), .B(G24), .Z(n936) );
  NAND2_X1 U1037 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1038 ( .A(KEYINPUT58), .B(n938), .ZN(n939) );
  NOR2_X1 U1039 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1040 ( .A(n941), .B(KEYINPUT61), .ZN(n942) );
  XOR2_X1 U1041 ( .A(n942), .B(KEYINPUT126), .Z(n1026) );
  INV_X1 U1042 ( .A(KEYINPUT124), .ZN(n943) );
  NOR2_X1 U1043 ( .A1(n1026), .A2(n943), .ZN(n969) );
  XNOR2_X1 U1044 ( .A(G1971), .B(KEYINPUT122), .ZN(n944) );
  XNOR2_X1 U1045 ( .A(n944), .B(G303), .ZN(n946) );
  NOR2_X1 U1046 ( .A1(n946), .A2(n945), .ZN(n953) );
  XNOR2_X1 U1047 ( .A(n947), .B(G1956), .ZN(n949) );
  XNOR2_X1 U1048 ( .A(G171), .B(G1961), .ZN(n948) );
  NAND2_X1 U1049 ( .A1(n949), .A2(n948), .ZN(n950) );
  NOR2_X1 U1050 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1051 ( .A1(n953), .A2(n952), .ZN(n956) );
  XNOR2_X1 U1052 ( .A(G1348), .B(n954), .ZN(n955) );
  NOR2_X1 U1053 ( .A1(n956), .A2(n955), .ZN(n958) );
  NAND2_X1 U1054 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1055 ( .A(KEYINPUT123), .B(n959), .ZN(n964) );
  XNOR2_X1 U1056 ( .A(G1966), .B(G168), .ZN(n961) );
  NAND2_X1 U1057 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1058 ( .A(n962), .B(KEYINPUT57), .ZN(n963) );
  NAND2_X1 U1059 ( .A1(n964), .A2(n963), .ZN(n967) );
  XNOR2_X1 U1060 ( .A(G1341), .B(n965), .ZN(n966) );
  NOR2_X1 U1061 ( .A1(n967), .A2(n966), .ZN(n1024) );
  NOR2_X1 U1062 ( .A1(KEYINPUT56), .A2(n1024), .ZN(n968) );
  NOR2_X1 U1063 ( .A1(n969), .A2(n968), .ZN(n970) );
  NOR2_X1 U1064 ( .A1(G16), .A2(n970), .ZN(n1033) );
  XOR2_X1 U1065 ( .A(KEYINPUT53), .B(KEYINPUT121), .Z(n984) );
  XNOR2_X1 U1066 ( .A(G27), .B(n971), .ZN(n975) );
  XNOR2_X1 U1067 ( .A(G1996), .B(G32), .ZN(n973) );
  XNOR2_X1 U1068 ( .A(G26), .B(G2067), .ZN(n972) );
  NOR2_X1 U1069 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1070 ( .A1(n975), .A2(n974), .ZN(n978) );
  XOR2_X1 U1071 ( .A(KEYINPUT119), .B(G2072), .Z(n976) );
  XNOR2_X1 U1072 ( .A(G33), .B(n976), .ZN(n977) );
  NOR2_X1 U1073 ( .A1(n978), .A2(n977), .ZN(n979) );
  XOR2_X1 U1074 ( .A(KEYINPUT120), .B(n979), .Z(n981) );
  XNOR2_X1 U1075 ( .A(G1991), .B(G25), .ZN(n980) );
  NOR2_X1 U1076 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1077 ( .A1(n982), .A2(G28), .ZN(n983) );
  XNOR2_X1 U1078 ( .A(n984), .B(n983), .ZN(n989) );
  XNOR2_X1 U1079 ( .A(G2084), .B(KEYINPUT54), .ZN(n985) );
  XNOR2_X1 U1080 ( .A(n985), .B(G34), .ZN(n987) );
  XNOR2_X1 U1081 ( .A(G35), .B(G2090), .ZN(n986) );
  NOR2_X1 U1082 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1083 ( .A1(n989), .A2(n988), .ZN(n990) );
  XOR2_X1 U1084 ( .A(KEYINPUT55), .B(n990), .Z(n991) );
  INV_X1 U1085 ( .A(G29), .ZN(n1020) );
  NAND2_X1 U1086 ( .A1(n991), .A2(n1020), .ZN(n992) );
  NAND2_X1 U1087 ( .A1(G11), .A2(n992), .ZN(n1023) );
  INV_X1 U1088 ( .A(n993), .ZN(n995) );
  NAND2_X1 U1089 ( .A1(n995), .A2(n994), .ZN(n1002) );
  XNOR2_X1 U1090 ( .A(G160), .B(G2084), .ZN(n997) );
  NAND2_X1 U1091 ( .A1(n997), .A2(n996), .ZN(n999) );
  NOR2_X1 U1092 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XOR2_X1 U1093 ( .A(KEYINPUT116), .B(n1000), .Z(n1001) );
  NOR2_X1 U1094 ( .A1(n1002), .A2(n1001), .ZN(n1016) );
  XOR2_X1 U1095 ( .A(G2090), .B(G162), .Z(n1003) );
  NOR2_X1 U1096 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XOR2_X1 U1097 ( .A(KEYINPUT51), .B(n1005), .Z(n1006) );
  NAND2_X1 U1098 ( .A1(n1007), .A2(n1006), .ZN(n1014) );
  XNOR2_X1 U1099 ( .A(G2072), .B(n1008), .ZN(n1010) );
  XNOR2_X1 U1100 ( .A(G164), .B(G2078), .ZN(n1009) );
  NAND2_X1 U1101 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XOR2_X1 U1102 ( .A(KEYINPUT50), .B(n1011), .Z(n1012) );
  XNOR2_X1 U1103 ( .A(KEYINPUT117), .B(n1012), .ZN(n1013) );
  NOR2_X1 U1104 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1105 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1106 ( .A(n1017), .B(KEYINPUT52), .ZN(n1018) );
  XNOR2_X1 U1107 ( .A(n1018), .B(KEYINPUT118), .ZN(n1019) );
  NOR2_X1 U1108 ( .A1(KEYINPUT55), .A2(n1019), .ZN(n1021) );
  NOR2_X1 U1109 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NOR2_X1 U1110 ( .A1(n1023), .A2(n1022), .ZN(n1031) );
  INV_X1 U1111 ( .A(n1024), .ZN(n1025) );
  NAND2_X1 U1112 ( .A1(n1025), .A2(KEYINPUT56), .ZN(n1028) );
  OR2_X1 U1113 ( .A1(KEYINPUT124), .A2(n1026), .ZN(n1027) );
  NAND2_X1 U1114 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1115 ( .A1(n1029), .A2(G16), .ZN(n1030) );
  NAND2_X1 U1116 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NOR2_X1 U1117 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  XOR2_X1 U1118 ( .A(KEYINPUT127), .B(n1034), .Z(n1035) );
  XNOR2_X1 U1119 ( .A(KEYINPUT62), .B(n1035), .ZN(G311) );
  INV_X1 U1120 ( .A(G311), .ZN(G150) );
endmodule

