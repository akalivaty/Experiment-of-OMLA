//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 0 0 1 1 1 0 0 1 1 0 1 1 0 0 0 1 1 0 0 1 0 0 0 0 0 0 1 0 0 0 1 1 1 0 1 1 1 0 1 1 0 1 0 0 1 1 0 0 1 0 0 0 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:33 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n755, new_n756, new_n757, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(new_n187), .B(KEYINPUT70), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT30), .ZN(new_n189));
  XOR2_X1   g003(.A(KEYINPUT0), .B(G128), .Z(new_n190));
  INV_X1    g004(.A(G146), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(KEYINPUT64), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT64), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G146), .ZN(new_n194));
  AOI21_X1  g008(.A(G143), .B1(new_n192), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G143), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n196), .A2(G146), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n190), .B1(new_n195), .B2(new_n197), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n192), .A2(new_n194), .A3(G143), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n196), .A2(G146), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n199), .A2(KEYINPUT0), .A3(G128), .A4(new_n200), .ZN(new_n201));
  AND3_X1   g015(.A1(new_n198), .A2(KEYINPUT65), .A3(new_n201), .ZN(new_n202));
  AOI21_X1  g016(.A(KEYINPUT65), .B1(new_n198), .B2(new_n201), .ZN(new_n203));
  INV_X1    g017(.A(G137), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n204), .A2(G134), .ZN(new_n205));
  INV_X1    g019(.A(G134), .ZN(new_n206));
  OAI21_X1  g020(.A(KEYINPUT11), .B1(new_n206), .B2(G137), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT11), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n208), .A2(new_n204), .A3(G134), .ZN(new_n209));
  AOI211_X1 g023(.A(G131), .B(new_n205), .C1(new_n207), .C2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G131), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n207), .A2(new_n209), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n206), .A2(G137), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n210), .A2(new_n214), .ZN(new_n215));
  NOR3_X1   g029(.A1(new_n202), .A2(new_n203), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n204), .A2(G134), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT66), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n217), .B1(new_n205), .B2(new_n218), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n213), .A2(KEYINPUT66), .ZN(new_n220));
  OAI21_X1  g034(.A(G131), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n205), .B1(new_n207), .B2(new_n209), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(new_n211), .ZN(new_n223));
  AND2_X1   g037(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT1), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n199), .A2(new_n225), .A3(G128), .A4(new_n200), .ZN(new_n226));
  INV_X1    g040(.A(G128), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n227), .B1(new_n199), .B2(KEYINPUT1), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n192), .A2(new_n194), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n197), .B1(new_n229), .B2(new_n196), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n226), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  AND2_X1   g045(.A1(new_n224), .A2(new_n231), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n189), .B1(new_n216), .B2(new_n232), .ZN(new_n233));
  XNOR2_X1  g047(.A(G116), .B(G119), .ZN(new_n234));
  INV_X1    g048(.A(G113), .ZN(new_n235));
  AND2_X1   g049(.A1(new_n235), .A2(KEYINPUT2), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n235), .A2(KEYINPUT2), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n234), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(G119), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G116), .ZN(new_n240));
  INV_X1    g054(.A(G116), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G119), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g057(.A(KEYINPUT2), .B(G113), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n238), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n231), .A2(KEYINPUT67), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT67), .ZN(new_n248));
  OAI211_X1 g062(.A(new_n248), .B(new_n226), .C1(new_n228), .C2(new_n230), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n247), .A2(new_n224), .A3(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n198), .A2(new_n201), .ZN(new_n251));
  OR2_X1    g065(.A1(new_n215), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n250), .A2(KEYINPUT30), .A3(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n233), .A2(new_n246), .A3(new_n253), .ZN(new_n254));
  AND2_X1   g068(.A1(new_n238), .A2(new_n245), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n250), .A2(new_n255), .A3(new_n252), .ZN(new_n256));
  NOR2_X1   g070(.A1(G237), .A2(G953), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G210), .ZN(new_n258));
  XNOR2_X1  g072(.A(new_n258), .B(KEYINPUT27), .ZN(new_n259));
  XNOR2_X1  g073(.A(KEYINPUT26), .B(G101), .ZN(new_n260));
  XNOR2_X1  g074(.A(new_n259), .B(new_n260), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n254), .A2(new_n256), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(KEYINPUT31), .ZN(new_n263));
  XOR2_X1   g077(.A(KEYINPUT68), .B(KEYINPUT31), .Z(new_n264));
  NAND4_X1  g078(.A1(new_n254), .A2(new_n256), .A3(new_n261), .A4(new_n264), .ZN(new_n265));
  AND2_X1   g079(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT69), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n267), .B(new_n246), .C1(new_n216), .C2(new_n232), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(new_n256), .ZN(new_n269));
  INV_X1    g083(.A(new_n203), .ZN(new_n270));
  INV_X1    g084(.A(new_n215), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n198), .A2(KEYINPUT65), .A3(new_n201), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n270), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n224), .A2(new_n231), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n267), .B1(new_n275), .B2(new_n246), .ZN(new_n276));
  OAI21_X1  g090(.A(KEYINPUT28), .B1(new_n269), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT28), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n256), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n261), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n188), .B1(new_n266), .B2(new_n282), .ZN(new_n283));
  AND2_X1   g097(.A1(new_n256), .A2(new_n278), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n250), .A2(new_n252), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(new_n246), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(new_n256), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n284), .B1(new_n287), .B2(KEYINPUT28), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT29), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n281), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(G902), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n203), .A2(new_n215), .ZN(new_n292));
  AOI22_X1  g106(.A1(new_n292), .A2(new_n272), .B1(new_n224), .B2(new_n231), .ZN(new_n293));
  OAI21_X1  g107(.A(KEYINPUT69), .B1(new_n293), .B2(new_n255), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n294), .A2(new_n256), .A3(new_n268), .ZN(new_n295));
  AOI211_X1 g109(.A(new_n281), .B(new_n284), .C1(new_n295), .C2(KEYINPUT28), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n254), .A2(new_n256), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n281), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(new_n289), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n291), .B1(new_n296), .B2(new_n299), .ZN(new_n300));
  AOI22_X1  g114(.A1(new_n283), .A2(KEYINPUT32), .B1(G472), .B2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n188), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n263), .A2(new_n265), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n261), .B1(new_n277), .B2(new_n279), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT32), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT71), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n305), .A2(KEYINPUT71), .A3(new_n306), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n301), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G221), .ZN(new_n312));
  XNOR2_X1  g126(.A(KEYINPUT9), .B(G234), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(G902), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n312), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(G469), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n317), .A2(new_n315), .ZN(new_n318));
  XNOR2_X1  g132(.A(G110), .B(G140), .ZN(new_n319));
  INV_X1    g133(.A(G953), .ZN(new_n320));
  AND2_X1   g134(.A1(new_n320), .A2(G227), .ZN(new_n321));
  XNOR2_X1  g135(.A(new_n319), .B(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT76), .ZN(new_n323));
  XNOR2_X1  g137(.A(G104), .B(G107), .ZN(new_n324));
  INV_X1    g138(.A(G101), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n323), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(G107), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G104), .ZN(new_n328));
  INV_X1    g142(.A(G104), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G107), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n331), .A2(KEYINPUT76), .A3(G101), .ZN(new_n332));
  OAI21_X1  g146(.A(KEYINPUT3), .B1(new_n329), .B2(G107), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT3), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n334), .A2(new_n327), .A3(G104), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n333), .A2(new_n335), .A3(new_n325), .A4(new_n330), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n326), .A2(new_n332), .A3(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(KEYINPUT1), .B1(new_n196), .B2(G146), .ZN(new_n339));
  AOI22_X1  g153(.A1(new_n199), .A2(new_n200), .B1(G128), .B2(new_n339), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n226), .B1(new_n340), .B2(KEYINPUT77), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n199), .A2(new_n200), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n339), .A2(G128), .ZN(new_n343));
  AND3_X1   g157(.A1(new_n342), .A2(KEYINPUT77), .A3(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n338), .B1(new_n341), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT10), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n333), .A2(new_n335), .A3(new_n330), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT4), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n348), .A2(new_n349), .A3(G101), .ZN(new_n350));
  AND3_X1   g164(.A1(new_n198), .A2(new_n350), .A3(new_n201), .ZN(new_n351));
  AND2_X1   g165(.A1(new_n336), .A2(KEYINPUT4), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n348), .A2(G101), .ZN(new_n353));
  AOI21_X1  g167(.A(KEYINPUT75), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  AND4_X1   g168(.A1(KEYINPUT75), .A2(new_n353), .A3(KEYINPUT4), .A4(new_n336), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n351), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n337), .A2(new_n346), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n247), .A2(new_n357), .A3(new_n249), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n347), .A2(new_n356), .A3(new_n215), .A4(new_n358), .ZN(new_n359));
  OAI211_X1 g173(.A(new_n337), .B(new_n226), .C1(new_n230), .C2(new_n228), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n345), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(KEYINPUT12), .B1(new_n361), .B2(new_n271), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT12), .ZN(new_n363));
  AOI211_X1 g177(.A(new_n363), .B(new_n215), .C1(new_n345), .C2(new_n360), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n359), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(new_n322), .ZN(new_n366));
  AND2_X1   g180(.A1(new_n359), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n347), .A2(new_n356), .A3(new_n358), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(new_n271), .ZN(new_n369));
  AOI22_X1  g183(.A1(new_n322), .A2(new_n365), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n318), .B1(new_n370), .B2(G469), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n362), .A2(new_n364), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n359), .A2(new_n366), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n366), .B1(new_n369), .B2(new_n359), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n317), .B(new_n315), .C1(new_n374), .C2(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n316), .B1(new_n371), .B2(new_n376), .ZN(new_n377));
  XNOR2_X1  g191(.A(G125), .B(G140), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(KEYINPUT16), .ZN(new_n379));
  INV_X1    g193(.A(G125), .ZN(new_n380));
  OR3_X1    g194(.A1(new_n380), .A2(KEYINPUT16), .A3(G140), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(new_n191), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n379), .A2(G146), .A3(new_n381), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(G143), .B1(new_n257), .B2(G214), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n257), .A2(G143), .A3(G214), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n390), .A2(KEYINPUT17), .A3(G131), .ZN(new_n391));
  INV_X1    g205(.A(new_n389), .ZN(new_n392));
  OAI21_X1  g206(.A(G131), .B1(new_n392), .B2(new_n387), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n388), .A2(new_n211), .A3(new_n389), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n386), .B(new_n391), .C1(KEYINPUT17), .C2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(KEYINPUT18), .A2(G131), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n388), .A2(new_n389), .A3(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n390), .A2(KEYINPUT18), .A3(G131), .ZN(new_n399));
  INV_X1    g213(.A(new_n229), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(new_n378), .ZN(new_n401));
  INV_X1    g215(.A(new_n378), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(G146), .ZN(new_n403));
  AND3_X1   g217(.A1(new_n401), .A2(new_n403), .A3(KEYINPUT81), .ZN(new_n404));
  AOI21_X1  g218(.A(KEYINPUT81), .B1(new_n401), .B2(new_n403), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n398), .B(new_n399), .C1(new_n404), .C2(new_n405), .ZN(new_n406));
  XNOR2_X1  g220(.A(G113), .B(G122), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n407), .B(new_n329), .ZN(new_n408));
  XOR2_X1   g222(.A(new_n408), .B(KEYINPUT83), .Z(new_n409));
  NAND3_X1  g223(.A1(new_n396), .A2(new_n406), .A3(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n408), .B1(new_n396), .B2(new_n406), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n315), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(G475), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT20), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT73), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n384), .A2(new_n417), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n379), .A2(KEYINPUT73), .A3(new_n381), .A4(G146), .ZN(new_n419));
  AND2_X1   g233(.A1(new_n378), .A2(KEYINPUT19), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n378), .A2(KEYINPUT19), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n400), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n395), .A2(new_n418), .A3(new_n419), .A4(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT82), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n406), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n408), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n424), .B1(new_n406), .B2(new_n423), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n410), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NOR2_X1   g243(.A1(G475), .A2(G902), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n416), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT85), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT84), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n416), .B1(new_n430), .B2(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n434), .B1(new_n433), .B2(new_n430), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n429), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n431), .B1(new_n432), .B2(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n429), .A2(KEYINPUT85), .A3(new_n435), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n415), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n196), .A2(G128), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n227), .A2(G143), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n440), .A2(new_n441), .A3(KEYINPUT88), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(KEYINPUT88), .B1(new_n440), .B2(new_n441), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n206), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n440), .A2(new_n441), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT88), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n448), .A2(G134), .A3(new_n442), .ZN(new_n449));
  XNOR2_X1  g263(.A(G116), .B(G122), .ZN(new_n450));
  AOI22_X1  g264(.A1(new_n445), .A2(new_n449), .B1(new_n327), .B2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT14), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n241), .A2(KEYINPUT14), .A3(G122), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n453), .A2(G107), .A3(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT90), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n453), .A2(KEYINPUT90), .A3(G107), .A4(new_n454), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n451), .A2(new_n459), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n450), .B(new_n327), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n448), .A2(new_n442), .ZN(new_n462));
  AOI21_X1  g276(.A(KEYINPUT89), .B1(new_n462), .B2(new_n206), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT89), .ZN(new_n464));
  AOI211_X1 g278(.A(new_n464), .B(G134), .C1(new_n448), .C2(new_n442), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n461), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT86), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT13), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n467), .B(new_n468), .C1(new_n227), .C2(G143), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(new_n441), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n467), .B1(new_n440), .B2(new_n468), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n227), .A2(G143), .ZN(new_n473));
  AOI22_X1  g287(.A1(new_n472), .A2(KEYINPUT87), .B1(KEYINPUT13), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT87), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n475), .B1(new_n470), .B2(new_n471), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n206), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n460), .B1(new_n466), .B2(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n314), .A2(G217), .A3(new_n320), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n479), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n460), .B(new_n481), .C1(new_n466), .C2(new_n477), .ZN(new_n482));
  AOI21_X1  g296(.A(G902), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(G478), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n485), .A2(KEYINPUT15), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n483), .B1(KEYINPUT15), .B2(new_n485), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(G234), .A2(G237), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n490), .A2(G952), .A3(new_n320), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n490), .A2(G902), .A3(G953), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(KEYINPUT21), .B(G898), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n492), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n489), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n377), .A2(new_n439), .A3(new_n497), .ZN(new_n498));
  OAI21_X1  g312(.A(G214), .B1(G237), .B2(G902), .ZN(new_n499));
  OAI21_X1  g313(.A(G210), .B1(G237), .B2(G902), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n246), .A2(new_n350), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n502), .B1(new_n354), .B2(new_n355), .ZN(new_n503));
  AND2_X1   g317(.A1(new_n234), .A2(KEYINPUT5), .ZN(new_n504));
  OAI21_X1  g318(.A(G113), .B1(new_n240), .B2(KEYINPUT5), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n238), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n506), .A2(new_n337), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  XNOR2_X1  g322(.A(G110), .B(G122), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n503), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n509), .A2(KEYINPUT78), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT75), .ZN(new_n512));
  AND2_X1   g326(.A1(new_n348), .A2(G101), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n336), .A2(KEYINPUT4), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n353), .A2(KEYINPUT75), .A3(KEYINPUT4), .A4(new_n336), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n501), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n511), .B1(new_n517), .B2(new_n507), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n510), .A2(new_n518), .A3(KEYINPUT6), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n251), .A2(G125), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n380), .B(new_n226), .C1(new_n228), .C2(new_n230), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n320), .A2(G224), .ZN(new_n523));
  XNOR2_X1  g337(.A(new_n523), .B(KEYINPUT79), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n522), .B(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT6), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n527), .B(new_n511), .C1(new_n517), .C2(new_n507), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n519), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(KEYINPUT80), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT80), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n519), .A2(new_n526), .A3(new_n531), .A4(new_n528), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n522), .A2(new_n525), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n509), .B(KEYINPUT8), .ZN(new_n535));
  AND2_X1   g349(.A1(new_n506), .A2(new_n337), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n535), .B1(new_n536), .B2(new_n507), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT7), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n522), .A2(new_n538), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n520), .A2(KEYINPUT7), .A3(new_n524), .A4(new_n521), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n534), .A2(new_n537), .A3(new_n539), .A4(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n510), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n315), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n500), .B1(new_n533), .B2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n500), .ZN(new_n546));
  AOI211_X1 g360(.A(new_n546), .B(new_n543), .C1(new_n530), .C2(new_n532), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n499), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n498), .A2(new_n548), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n239), .A2(G128), .ZN(new_n550));
  OR2_X1    g364(.A1(new_n550), .A2(KEYINPUT72), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(KEYINPUT72), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n239), .A2(G128), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(KEYINPUT24), .B(G110), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n227), .A2(KEYINPUT23), .A3(G119), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n553), .B(new_n557), .C1(new_n550), .C2(KEYINPUT23), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n556), .B1(G110), .B2(new_n558), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n559), .A2(new_n418), .A3(new_n419), .A4(new_n401), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n558), .A2(G110), .ZN(new_n561));
  OAI211_X1 g375(.A(new_n385), .B(new_n561), .C1(new_n555), .C2(new_n554), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  XNOR2_X1  g377(.A(KEYINPUT22), .B(G137), .ZN(new_n564));
  INV_X1    g378(.A(G234), .ZN(new_n565));
  NOR3_X1   g379(.A1(new_n312), .A2(new_n565), .A3(G953), .ZN(new_n566));
  XOR2_X1   g380(.A(new_n564), .B(new_n566), .Z(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n563), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n560), .A2(new_n562), .A3(new_n567), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n569), .A2(new_n315), .A3(new_n570), .ZN(new_n571));
  OR2_X1    g385(.A1(new_n571), .A2(KEYINPUT25), .ZN(new_n572));
  OAI21_X1  g386(.A(G217), .B1(new_n565), .B2(G902), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n573), .B1(new_n571), .B2(KEYINPUT25), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n573), .A2(new_n315), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n569), .A2(new_n570), .A3(new_n578), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n579), .B(KEYINPUT74), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n576), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n311), .A2(new_n549), .A3(new_n581), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n582), .B(G101), .ZN(G3));
  INV_X1    g397(.A(KEYINPUT96), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n429), .A2(new_n430), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(KEYINPUT20), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n436), .A2(new_n432), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n586), .A2(new_n587), .A3(new_n438), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(new_n414), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT33), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n590), .B1(new_n478), .B2(new_n479), .ZN(new_n591));
  OAI21_X1  g405(.A(KEYINPUT86), .B1(new_n473), .B2(KEYINPUT13), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n592), .A2(KEYINPUT87), .A3(new_n441), .A4(new_n469), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n593), .B1(new_n468), .B2(new_n440), .ZN(new_n594));
  INV_X1    g408(.A(new_n476), .ZN(new_n595));
  OAI21_X1  g409(.A(G134), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  OAI211_X1 g410(.A(new_n596), .B(new_n461), .C1(new_n463), .C2(new_n465), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT93), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n597), .A2(new_n598), .A3(new_n460), .A4(new_n481), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n482), .A2(KEYINPUT93), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n591), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT94), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n591), .A2(new_n599), .A3(new_n600), .A4(KEYINPUT94), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g419(.A(KEYINPUT33), .B1(new_n480), .B2(new_n482), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n485), .A2(G902), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n605), .A2(KEYINPUT95), .A3(new_n607), .A4(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n484), .A2(new_n485), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n606), .B1(new_n603), .B2(new_n604), .ZN(new_n612));
  AOI21_X1  g426(.A(KEYINPUT95), .B1(new_n612), .B2(new_n608), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n589), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n496), .ZN(new_n616));
  OAI211_X1 g430(.A(new_n499), .B(new_n616), .C1(new_n545), .C2(new_n547), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n584), .B1(new_n615), .B2(new_n618), .ZN(new_n619));
  NOR3_X1   g433(.A1(new_n614), .A2(KEYINPUT96), .A3(new_n617), .ZN(new_n620));
  OR2_X1    g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT92), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n315), .B1(new_n303), .B2(new_n304), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(KEYINPUT91), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n284), .B1(new_n295), .B2(KEYINPUT28), .ZN(new_n625));
  OAI211_X1 g439(.A(new_n263), .B(new_n265), .C1(new_n625), .C2(new_n261), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT91), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n626), .A2(new_n627), .A3(new_n315), .ZN(new_n628));
  AND3_X1   g442(.A1(new_n624), .A2(G472), .A3(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n377), .A2(new_n581), .A3(new_n305), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n622), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  AND3_X1   g445(.A1(new_n377), .A2(new_n581), .A3(new_n305), .ZN(new_n632));
  INV_X1    g446(.A(G472), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n633), .B1(new_n623), .B2(KEYINPUT91), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n628), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n632), .A2(KEYINPUT92), .A3(new_n635), .ZN(new_n636));
  AND3_X1   g450(.A1(new_n621), .A2(new_n631), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(KEYINPUT34), .B(G104), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G6));
  XNOR2_X1  g453(.A(new_n496), .B(KEYINPUT97), .ZN(new_n640));
  OAI211_X1 g454(.A(new_n499), .B(new_n640), .C1(new_n545), .C2(new_n547), .ZN(new_n641));
  AND3_X1   g455(.A1(new_n429), .A2(new_n416), .A3(new_n430), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n414), .B1(new_n642), .B2(new_n431), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(new_n489), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n631), .A2(new_n636), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(G107), .ZN(new_n648));
  XNOR2_X1  g462(.A(KEYINPUT98), .B(KEYINPUT35), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G9));
  AOI21_X1  g464(.A(new_n283), .B1(new_n634), .B2(new_n628), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n568), .A2(KEYINPUT36), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n563), .B(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(new_n578), .ZN(new_n654));
  AND2_X1   g468(.A1(new_n575), .A2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n549), .A2(new_n651), .A3(new_n656), .ZN(new_n657));
  XOR2_X1   g471(.A(KEYINPUT37), .B(G110), .Z(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(KEYINPUT99), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n657), .B(new_n659), .ZN(G12));
  INV_X1    g474(.A(new_n548), .ZN(new_n661));
  OR2_X1    g475(.A1(new_n493), .A2(G900), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n645), .B1(new_n491), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n370), .A2(G469), .ZN(new_n664));
  INV_X1    g478(.A(new_n318), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n664), .A2(new_n376), .A3(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n316), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n668), .A2(new_n655), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n311), .A2(new_n661), .A3(new_n663), .A4(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G128), .ZN(G30));
  INV_X1    g485(.A(new_n489), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n672), .B1(new_n414), .B2(new_n588), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n673), .A2(new_n499), .A3(new_n655), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n662), .A2(new_n491), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(KEYINPUT39), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n377), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n674), .B1(new_n677), .B2(KEYINPUT40), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n533), .A2(new_n544), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(new_n546), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n533), .A2(new_n500), .A3(new_n544), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(KEYINPUT38), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n283), .A2(KEYINPUT32), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n315), .B1(new_n287), .B2(new_n261), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n281), .B1(new_n254), .B2(new_n256), .ZN(new_n686));
  OAI21_X1  g500(.A(G472), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n309), .A2(new_n684), .A3(new_n310), .A4(new_n687), .ZN(new_n688));
  OR2_X1    g502(.A1(new_n677), .A2(KEYINPUT40), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n678), .A2(new_n683), .A3(new_n688), .A4(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G143), .ZN(G45));
  OAI211_X1 g505(.A(new_n589), .B(new_n675), .C1(new_n611), .C2(new_n613), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n311), .A2(new_n693), .A3(new_n661), .A4(new_n669), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G146), .ZN(G48));
  INV_X1    g509(.A(new_n581), .ZN(new_n696));
  AOI211_X1 g510(.A(new_n308), .B(KEYINPUT32), .C1(new_n626), .C2(new_n302), .ZN(new_n697));
  AOI21_X1  g511(.A(KEYINPUT71), .B1(new_n305), .B2(new_n306), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n696), .B1(new_n699), .B2(new_n301), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n315), .B1(new_n374), .B2(new_n375), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(G469), .ZN(new_n702));
  AND3_X1   g516(.A1(new_n702), .A2(new_n667), .A3(new_n376), .ZN(new_n703));
  OAI211_X1 g517(.A(new_n700), .B(new_n703), .C1(new_n619), .C2(new_n620), .ZN(new_n704));
  XNOR2_X1  g518(.A(KEYINPUT41), .B(G113), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n704), .B(new_n705), .ZN(G15));
  NAND3_X1  g520(.A1(new_n700), .A2(new_n646), .A3(new_n703), .ZN(new_n707));
  XNOR2_X1  g521(.A(KEYINPUT100), .B(G116), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n707), .B(new_n708), .ZN(G18));
  NAND3_X1  g523(.A1(new_n656), .A2(new_n439), .A3(new_n497), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n710), .B1(new_n699), .B2(new_n301), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT101), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n702), .A2(new_n667), .A3(new_n376), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n712), .B1(new_n548), .B2(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n682), .A2(new_n703), .A3(KEYINPUT101), .A4(new_n499), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n711), .A2(new_n716), .ZN(new_n717));
  XOR2_X1   g531(.A(KEYINPUT102), .B(G119), .Z(new_n718));
  XNOR2_X1  g532(.A(new_n717), .B(new_n718), .ZN(G21));
  NAND3_X1  g533(.A1(new_n673), .A2(new_n682), .A3(new_n499), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n703), .A2(new_n640), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT103), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n278), .B1(new_n286), .B2(new_n256), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n723), .B1(new_n724), .B2(new_n284), .ZN(new_n725));
  INV_X1    g539(.A(new_n256), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n255), .B1(new_n250), .B2(new_n252), .ZN(new_n727));
  OAI21_X1  g541(.A(KEYINPUT28), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n728), .A2(KEYINPUT103), .A3(new_n279), .ZN(new_n729));
  AND3_X1   g543(.A1(new_n725), .A2(new_n281), .A3(new_n729), .ZN(new_n730));
  OAI211_X1 g544(.A(KEYINPUT104), .B(new_n302), .C1(new_n730), .C2(new_n303), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n623), .A2(G472), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n725), .A2(new_n729), .A3(new_n281), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n266), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g549(.A(KEYINPUT104), .B1(new_n735), .B2(new_n302), .ZN(new_n736));
  NOR3_X1   g550(.A1(new_n733), .A2(new_n696), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n722), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G122), .ZN(G24));
  NOR3_X1   g553(.A1(new_n733), .A2(new_n655), .A3(new_n736), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n716), .A2(new_n740), .A3(new_n693), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G125), .ZN(G27));
  AOI21_X1  g556(.A(new_n696), .B1(new_n301), .B2(new_n307), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n680), .A2(new_n499), .A3(new_n681), .ZN(new_n744));
  OAI21_X1  g558(.A(KEYINPUT105), .B1(new_n744), .B2(new_n668), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n545), .A2(new_n547), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT105), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n746), .A2(new_n377), .A3(new_n747), .A4(new_n499), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n743), .A2(new_n693), .A3(new_n745), .A4(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(KEYINPUT42), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n692), .A2(KEYINPUT42), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n700), .A2(new_n745), .A3(new_n748), .A4(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(new_n211), .ZN(G33));
  NAND2_X1  g568(.A1(new_n311), .A2(new_n581), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n745), .A2(new_n748), .ZN(new_n756));
  INV_X1    g570(.A(new_n663), .ZN(new_n757));
  NOR3_X1   g571(.A1(new_n755), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(new_n206), .ZN(G36));
  OR2_X1    g573(.A1(new_n370), .A2(KEYINPUT45), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n370), .A2(KEYINPUT45), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n760), .A2(G469), .A3(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT106), .ZN(new_n763));
  OR2_X1    g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n762), .A2(new_n763), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n318), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(KEYINPUT46), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT46), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n762), .B(KEYINPUT106), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n768), .B1(new_n769), .B2(new_n318), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n767), .A2(new_n770), .A3(new_n376), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n771), .A2(new_n667), .A3(new_n676), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(new_n611), .ZN(new_n774));
  INV_X1    g588(.A(new_n613), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n589), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(KEYINPUT43), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n651), .A2(new_n655), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT44), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n744), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n776), .A2(KEYINPUT43), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n776), .A2(KEYINPUT43), .ZN(new_n784));
  OAI211_X1 g598(.A(KEYINPUT44), .B(new_n778), .C1(new_n783), .C2(new_n784), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n785), .A2(KEYINPUT107), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n785), .A2(KEYINPUT107), .ZN(new_n787));
  OAI211_X1 g601(.A(new_n773), .B(new_n781), .C1(new_n786), .C2(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G137), .ZN(G39));
  NOR4_X1   g603(.A1(new_n311), .A2(new_n692), .A3(new_n581), .A4(new_n744), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n771), .A2(KEYINPUT47), .A3(new_n667), .ZN(new_n791));
  INV_X1    g605(.A(new_n791), .ZN(new_n792));
  AOI21_X1  g606(.A(KEYINPUT47), .B1(new_n771), .B2(new_n667), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n790), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G140), .ZN(G42));
  INV_X1    g609(.A(new_n683), .ZN(new_n796));
  INV_X1    g610(.A(new_n688), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n581), .A2(new_n499), .A3(new_n667), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n702), .A2(new_n376), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n799), .A2(KEYINPUT49), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n799), .A2(KEYINPUT49), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n798), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n796), .A2(new_n797), .A3(new_n776), .A4(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n740), .A2(new_n693), .A3(new_n745), .A4(new_n748), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n487), .A2(new_n488), .A3(new_n675), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n643), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n746), .A2(new_n499), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(KEYINPUT108), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT108), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n746), .A2(new_n809), .A3(new_n499), .A4(new_n806), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n311), .A2(new_n808), .A3(new_n669), .A4(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n804), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n812), .A2(new_n758), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n311), .A2(new_n581), .A3(new_n745), .A4(new_n748), .ZN(new_n814));
  INV_X1    g628(.A(new_n814), .ZN(new_n815));
  AOI22_X1  g629(.A1(new_n815), .A2(new_n751), .B1(new_n749), .B2(KEYINPUT42), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n439), .A2(new_n489), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n641), .B1(new_n614), .B2(new_n817), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n631), .A2(new_n636), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n582), .A2(new_n657), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n813), .A2(new_n816), .A3(new_n821), .ZN(new_n822));
  AOI22_X1  g636(.A1(new_n711), .A2(new_n716), .B1(new_n722), .B2(new_n737), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n704), .A2(new_n823), .A3(new_n707), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n720), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n377), .A2(new_n655), .A3(new_n675), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n826), .A2(new_n688), .A3(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n741), .A2(new_n694), .A3(new_n670), .A4(new_n828), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n829), .A2(KEYINPUT52), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n829), .A2(KEYINPUT52), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT52), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n833), .B1(new_n741), .B2(new_n670), .ZN(new_n834));
  INV_X1    g648(.A(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n825), .A2(KEYINPUT53), .A3(new_n832), .A4(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT54), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT53), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n804), .B(new_n811), .C1(new_n757), .C2(new_n814), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n753), .A2(new_n839), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n704), .A2(new_n823), .A3(new_n707), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n840), .A2(new_n841), .A3(new_n821), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n741), .A2(new_n670), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n843), .A2(new_n833), .A3(new_n694), .A4(new_n828), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n829), .A2(KEYINPUT52), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n838), .B1(new_n842), .B2(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n836), .A2(new_n837), .A3(new_n847), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n842), .A2(new_n846), .A3(new_n838), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT109), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n850), .B1(new_n822), .B2(new_n824), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n830), .A2(new_n831), .A3(new_n834), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n840), .A2(new_n841), .A3(KEYINPUT109), .A4(new_n821), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n849), .B1(new_n854), .B2(new_n838), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n848), .B1(new_n855), .B2(new_n837), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(KEYINPUT110), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT110), .ZN(new_n858));
  OAI211_X1 g672(.A(new_n858), .B(new_n848), .C1(new_n855), .C2(new_n837), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n744), .A2(new_n713), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n797), .A2(new_n581), .A3(new_n492), .A4(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT112), .ZN(new_n862));
  OR2_X1    g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n861), .A2(new_n862), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n611), .A2(new_n589), .A3(new_n613), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n777), .A2(new_n492), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n867), .A2(new_n740), .A3(new_n860), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n777), .A2(new_n492), .A3(new_n737), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n683), .A2(new_n499), .A3(new_n713), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT50), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n870), .A2(KEYINPUT50), .A3(new_n871), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n869), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(new_n744), .ZN(new_n877));
  INV_X1    g691(.A(new_n793), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n878), .A2(new_n791), .ZN(new_n879));
  INV_X1    g693(.A(new_n799), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n316), .B1(new_n880), .B2(KEYINPUT111), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n881), .B1(KEYINPUT111), .B2(new_n880), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n877), .B(new_n870), .C1(new_n879), .C2(new_n882), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n876), .A2(new_n883), .A3(KEYINPUT51), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n863), .A2(new_n615), .A3(new_n864), .ZN(new_n885));
  INV_X1    g699(.A(G952), .ZN(new_n886));
  AOI211_X1 g700(.A(new_n886), .B(G953), .C1(new_n870), .C2(new_n716), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n867), .A2(new_n743), .A3(new_n860), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(KEYINPUT113), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT48), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT113), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n867), .A2(new_n891), .A3(new_n743), .A4(new_n860), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n889), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n890), .B1(new_n889), .B2(new_n892), .ZN(new_n894));
  OAI211_X1 g708(.A(new_n885), .B(new_n887), .C1(new_n893), .C2(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(KEYINPUT51), .B1(new_n876), .B2(new_n883), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n884), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n857), .A2(new_n859), .A3(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT114), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n857), .A2(KEYINPUT114), .A3(new_n897), .A4(new_n859), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n886), .A2(new_n320), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n803), .B1(new_n900), .B2(new_n903), .ZN(G75));
  NAND2_X1  g718(.A1(new_n519), .A2(new_n528), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n905), .B(new_n526), .ZN(new_n906));
  XNOR2_X1  g720(.A(KEYINPUT115), .B(KEYINPUT55), .ZN(new_n907));
  XOR2_X1   g721(.A(new_n906), .B(new_n907), .Z(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n315), .B1(new_n836), .B2(new_n847), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n910), .A2(G210), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n909), .B1(new_n911), .B2(KEYINPUT56), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n320), .A2(G952), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n911), .A2(KEYINPUT56), .A3(new_n909), .ZN(new_n916));
  OAI21_X1  g730(.A(KEYINPUT116), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(new_n916), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT116), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n918), .A2(new_n919), .A3(new_n912), .A4(new_n914), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n917), .A2(new_n920), .ZN(G51));
  NAND2_X1  g735(.A1(new_n836), .A2(new_n847), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(KEYINPUT54), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n923), .A2(new_n848), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n318), .B(KEYINPUT57), .Z(new_n925));
  OAI22_X1  g739(.A1(new_n924), .A2(new_n925), .B1(new_n375), .B2(new_n374), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n910), .A2(new_n769), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n913), .B1(new_n926), .B2(new_n927), .ZN(G54));
  NAND2_X1  g742(.A1(KEYINPUT58), .A2(G475), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n929), .B(KEYINPUT117), .Z(new_n930));
  AND2_X1   g744(.A1(new_n910), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n914), .B1(new_n931), .B2(new_n429), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n932), .B1(new_n429), .B2(new_n931), .ZN(G60));
  NAND2_X1  g747(.A1(new_n857), .A2(new_n859), .ZN(new_n934));
  XNOR2_X1  g748(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n485), .A2(new_n315), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n935), .B(new_n936), .Z(new_n937));
  INV_X1    g751(.A(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n612), .B1(new_n934), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n612), .A2(new_n938), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n914), .B1(new_n924), .B2(new_n940), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n939), .A2(new_n941), .ZN(G63));
  NAND2_X1  g756(.A1(G217), .A2(G902), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n943), .B(KEYINPUT60), .Z(new_n944));
  NAND2_X1  g758(.A1(new_n922), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(KEYINPUT119), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT119), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n922), .A2(new_n947), .A3(new_n944), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(new_n653), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n569), .A2(new_n570), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n946), .A2(new_n951), .A3(new_n948), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n950), .A2(new_n952), .A3(new_n914), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT61), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n950), .A2(new_n952), .A3(KEYINPUT61), .A4(new_n914), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(new_n956), .ZN(G66));
  INV_X1    g771(.A(G224), .ZN(new_n958));
  OAI21_X1  g772(.A(G953), .B1(new_n495), .B2(new_n958), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT120), .Z(new_n960));
  NAND2_X1  g774(.A1(new_n841), .A2(new_n821), .ZN(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n960), .B1(new_n962), .B2(G953), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n905), .B1(G898), .B2(new_n320), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n963), .B(new_n964), .ZN(G69));
  INV_X1    g779(.A(KEYINPUT124), .ZN(new_n966));
  AND2_X1   g780(.A1(new_n233), .A2(new_n253), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n420), .A2(new_n421), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n967), .B(new_n968), .Z(new_n969));
  INV_X1    g783(.A(new_n969), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n843), .A2(new_n690), .A3(new_n694), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n971), .A2(KEYINPUT62), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n744), .A2(new_n668), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n614), .A2(new_n817), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n700), .A2(new_n676), .A3(new_n973), .A4(new_n974), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n975), .B(KEYINPUT122), .Z(new_n976));
  AND4_X1   g790(.A1(new_n788), .A2(new_n794), .A3(new_n972), .A4(new_n976), .ZN(new_n977));
  AND2_X1   g791(.A1(new_n843), .A2(new_n694), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT62), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n978), .A2(KEYINPUT121), .A3(new_n979), .A4(new_n690), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT121), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n981), .B1(new_n971), .B2(KEYINPUT62), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(KEYINPUT123), .B1(new_n977), .B2(new_n983), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n788), .A2(new_n794), .A3(new_n972), .A4(new_n976), .ZN(new_n985));
  AND2_X1   g799(.A1(new_n980), .A2(new_n982), .ZN(new_n986));
  INV_X1    g800(.A(KEYINPUT123), .ZN(new_n987));
  NOR3_X1   g801(.A1(new_n985), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n984), .A2(new_n988), .ZN(new_n989));
  OAI211_X1 g803(.A(new_n966), .B(new_n970), .C1(new_n989), .C2(G953), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n977), .A2(KEYINPUT123), .A3(new_n983), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n987), .B1(new_n985), .B2(new_n986), .ZN(new_n992));
  AOI21_X1  g806(.A(G953), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  OAI21_X1  g807(.A(KEYINPUT124), .B1(new_n993), .B2(new_n969), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n970), .B1(G900), .B2(G953), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n773), .A2(new_n826), .A3(new_n743), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n753), .A2(new_n758), .ZN(new_n997));
  AND3_X1   g811(.A1(new_n794), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  AND3_X1   g812(.A1(new_n788), .A2(KEYINPUT125), .A3(new_n978), .ZN(new_n999));
  AOI21_X1  g813(.A(KEYINPUT125), .B1(new_n788), .B2(new_n978), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n998), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n995), .B1(new_n1001), .B2(G953), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n990), .A2(new_n994), .A3(new_n1002), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n320), .B1(G227), .B2(G900), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g819(.A(new_n1004), .ZN(new_n1006));
  NAND4_X1  g820(.A1(new_n990), .A2(new_n994), .A3(new_n1006), .A4(new_n1002), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1005), .A2(new_n1007), .ZN(G72));
  NAND2_X1  g822(.A1(G472), .A2(G902), .ZN(new_n1009));
  XOR2_X1   g823(.A(new_n1009), .B(KEYINPUT63), .Z(new_n1010));
  OAI21_X1  g824(.A(new_n1010), .B1(new_n1001), .B2(new_n961), .ZN(new_n1011));
  NAND4_X1  g825(.A1(new_n1011), .A2(new_n256), .A3(new_n281), .A4(new_n254), .ZN(new_n1012));
  INV_X1    g826(.A(new_n262), .ZN(new_n1013));
  NOR2_X1   g827(.A1(new_n1013), .A2(KEYINPUT127), .ZN(new_n1014));
  XOR2_X1   g828(.A(new_n1014), .B(new_n298), .Z(new_n1015));
  NAND2_X1  g829(.A1(new_n1015), .A2(new_n1010), .ZN(new_n1016));
  OAI211_X1 g830(.A(new_n1012), .B(new_n914), .C1(new_n855), .C2(new_n1016), .ZN(new_n1017));
  INV_X1    g831(.A(new_n1010), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1018), .B1(new_n989), .B2(new_n962), .ZN(new_n1019));
  INV_X1    g833(.A(KEYINPUT126), .ZN(new_n1020));
  OR2_X1    g834(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g835(.A(new_n686), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n1022), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n1017), .B1(new_n1021), .B2(new_n1023), .ZN(G57));
endmodule


