//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 1 1 0 1 0 1 1 1 0 0 1 1 1 1 1 0 1 0 0 1 0 1 1 1 1 1 0 1 1 0 1 1 0 0 1 1 0 0 1 1 1 0 0 1 1 0 0 0 1 1 1 1 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:29 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n510, new_n511,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n543, new_n544,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n564, new_n565, new_n566, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n595,
    new_n596, new_n599, new_n600, new_n601, new_n603, new_n604, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1186, new_n1187;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT65), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(G125), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  OAI211_X1 g043(.A(G137), .B(new_n463), .C1(new_n464), .C2(new_n465), .ZN(new_n469));
  AND2_X1   g044(.A1(new_n463), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G101), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n468), .A2(new_n472), .ZN(G160));
  OR2_X1    g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n463), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n463), .A2(G112), .ZN(new_n478));
  OAI21_X1  g053(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n479));
  AOI21_X1  g054(.A(G2105), .B1(new_n474), .B2(new_n475), .ZN(new_n480));
  AND3_X1   g055(.A1(new_n480), .A2(KEYINPUT67), .A3(G136), .ZN(new_n481));
  AOI21_X1  g056(.A(KEYINPUT67), .B1(new_n480), .B2(G136), .ZN(new_n482));
  OAI221_X1 g057(.A(new_n477), .B1(new_n478), .B2(new_n479), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT68), .ZN(G162));
  OAI211_X1 g059(.A(G126), .B(G2105), .C1(new_n464), .C2(new_n465), .ZN(new_n485));
  INV_X1    g060(.A(G114), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(G138), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n491), .B1(new_n464), .B2(new_n465), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n491), .B(new_n494), .C1(new_n465), .C2(new_n464), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n489), .B1(new_n493), .B2(new_n495), .ZN(G164));
  OR2_X1    g071(.A1(KEYINPUT5), .A2(G543), .ZN(new_n497));
  NAND2_X1  g072(.A1(KEYINPUT5), .A2(G543), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI22_X1  g074(.A1(new_n499), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n500));
  INV_X1    g075(.A(G651), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  XNOR2_X1  g077(.A(KEYINPUT6), .B(G651), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n499), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(G88), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n503), .A2(G543), .ZN(new_n506));
  INV_X1    g081(.A(G50), .ZN(new_n507));
  OAI22_X1  g082(.A1(new_n504), .A2(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n502), .A2(new_n508), .ZN(G166));
  NAND3_X1  g084(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n510));
  XNOR2_X1  g085(.A(new_n510), .B(KEYINPUT7), .ZN(new_n511));
  INV_X1    g086(.A(G51), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n511), .B1(new_n506), .B2(new_n512), .ZN(new_n513));
  AND2_X1   g088(.A1(new_n497), .A2(new_n498), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n503), .A2(G89), .ZN(new_n515));
  NAND2_X1  g090(.A1(G63), .A2(G651), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  OR2_X1    g092(.A1(new_n513), .A2(new_n517), .ZN(G286));
  INV_X1    g093(.A(G286), .ZN(G168));
  INV_X1    g094(.A(KEYINPUT69), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n499), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n521), .A2(new_n501), .ZN(new_n522));
  INV_X1    g097(.A(G90), .ZN(new_n523));
  INV_X1    g098(.A(G52), .ZN(new_n524));
  OAI22_X1  g099(.A1(new_n504), .A2(new_n523), .B1(new_n506), .B2(new_n524), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n520), .B1(new_n522), .B2(new_n525), .ZN(new_n526));
  OR2_X1    g101(.A1(KEYINPUT6), .A2(G651), .ZN(new_n527));
  NAND2_X1  g102(.A1(KEYINPUT6), .A2(G651), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n527), .A2(new_n528), .B1(new_n497), .B2(new_n498), .ZN(new_n529));
  INV_X1    g104(.A(G543), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n530), .B1(new_n527), .B2(new_n528), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n529), .A2(G90), .B1(new_n531), .B2(G52), .ZN(new_n532));
  OAI211_X1 g107(.A(new_n532), .B(KEYINPUT69), .C1(new_n501), .C2(new_n521), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n526), .A2(new_n533), .ZN(G171));
  AOI22_X1  g109(.A1(new_n499), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n535), .A2(new_n501), .ZN(new_n536));
  INV_X1    g111(.A(G81), .ZN(new_n537));
  INV_X1    g112(.A(G43), .ZN(new_n538));
  OAI22_X1  g113(.A1(new_n504), .A2(new_n537), .B1(new_n506), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G860), .ZN(G153));
  NAND4_X1  g116(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g117(.A1(G1), .A2(G3), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT8), .ZN(new_n544));
  NAND4_X1  g119(.A1(G319), .A2(G483), .A3(G661), .A4(new_n544), .ZN(G188));
  INV_X1    g120(.A(G53), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT70), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT9), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NOR2_X1   g124(.A1(KEYINPUT70), .A2(KEYINPUT9), .ZN(new_n550));
  OAI22_X1  g125(.A1(new_n506), .A2(new_n546), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  OAI211_X1 g126(.A(new_n531), .B(G53), .C1(new_n547), .C2(new_n548), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n499), .A2(G65), .ZN(new_n554));
  INV_X1    g129(.A(G78), .ZN(new_n555));
  OAI21_X1  g130(.A(KEYINPUT71), .B1(new_n555), .B2(new_n530), .ZN(new_n556));
  OR3_X1    g131(.A1(new_n555), .A2(new_n530), .A3(KEYINPUT71), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n554), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G651), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n529), .A2(G91), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n553), .A2(new_n559), .A3(new_n560), .ZN(G299));
  INV_X1    g136(.A(G171), .ZN(G301));
  INV_X1    g137(.A(G166), .ZN(G303));
  NAND2_X1  g138(.A1(new_n529), .A2(G87), .ZN(new_n564));
  OAI21_X1  g139(.A(G651), .B1(new_n499), .B2(G74), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n531), .A2(G49), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(G288));
  AOI22_X1  g142(.A1(new_n529), .A2(G86), .B1(new_n531), .B2(G48), .ZN(new_n568));
  NAND2_X1  g143(.A1(G73), .A2(G543), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT72), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n569), .B(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(G61), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n572), .B1(new_n497), .B2(new_n498), .ZN(new_n573));
  OAI21_X1  g148(.A(G651), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n568), .A2(new_n574), .ZN(G305));
  AOI22_X1  g150(.A1(new_n499), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n576), .A2(new_n501), .ZN(new_n577));
  XNOR2_X1  g152(.A(KEYINPUT73), .B(G85), .ZN(new_n578));
  INV_X1    g153(.A(G47), .ZN(new_n579));
  OAI22_X1  g154(.A1(new_n504), .A2(new_n578), .B1(new_n506), .B2(new_n579), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(G290));
  AOI22_X1  g157(.A1(new_n499), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n583));
  INV_X1    g158(.A(G54), .ZN(new_n584));
  OAI22_X1  g159(.A1(new_n583), .A2(new_n501), .B1(new_n584), .B2(new_n506), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT74), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  OAI221_X1 g162(.A(KEYINPUT74), .B1(new_n506), .B2(new_n584), .C1(new_n583), .C2(new_n501), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AND3_X1   g164(.A1(new_n499), .A2(new_n503), .A3(G92), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n590), .B(KEYINPUT10), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  MUX2_X1   g167(.A(new_n592), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g168(.A(new_n592), .B(G301), .S(G868), .Z(G321));
  NAND2_X1  g169(.A1(G286), .A2(G868), .ZN(new_n595));
  INV_X1    g170(.A(G299), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n596), .B2(G868), .ZN(G297));
  OAI21_X1  g172(.A(new_n595), .B1(new_n596), .B2(G868), .ZN(G280));
  NOR2_X1   g173(.A1(new_n592), .A2(G559), .ZN(new_n599));
  INV_X1    g174(.A(new_n592), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n599), .B1(G860), .B2(new_n600), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n601), .B(KEYINPUT75), .ZN(G148));
  NOR3_X1   g177(.A1(new_n536), .A2(new_n539), .A3(G868), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n599), .B(KEYINPUT76), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n603), .B1(new_n604), .B2(G868), .ZN(G323));
  XNOR2_X1  g180(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XNOR2_X1  g181(.A(KEYINPUT3), .B(G2104), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n607), .A2(new_n470), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT12), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT13), .ZN(new_n610));
  INV_X1    g185(.A(G2100), .ZN(new_n611));
  OR2_X1    g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n610), .A2(new_n611), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n480), .A2(G135), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n476), .A2(G123), .ZN(new_n615));
  OR2_X1    g190(.A1(G99), .A2(G2105), .ZN(new_n616));
  OAI211_X1 g191(.A(new_n616), .B(G2104), .C1(G111), .C2(new_n463), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n614), .A2(new_n615), .A3(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(G2096), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n618), .B(new_n619), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n612), .A2(new_n613), .A3(new_n620), .ZN(G156));
  XOR2_X1   g196(.A(G2451), .B(G2454), .Z(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT16), .ZN(new_n623));
  XNOR2_X1  g198(.A(G1341), .B(G1348), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n623), .B(new_n624), .ZN(new_n625));
  INV_X1    g200(.A(KEYINPUT14), .ZN(new_n626));
  XNOR2_X1  g201(.A(G2427), .B(G2438), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2430), .ZN(new_n628));
  XNOR2_X1  g203(.A(KEYINPUT15), .B(G2435), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n626), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n630), .B1(new_n629), .B2(new_n628), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n625), .B(new_n631), .Z(new_n632));
  XNOR2_X1  g207(.A(G2443), .B(G2446), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n632), .A2(new_n633), .ZN(new_n635));
  AND3_X1   g210(.A1(new_n634), .A2(G14), .A3(new_n635), .ZN(G401));
  INV_X1    g211(.A(KEYINPUT18), .ZN(new_n637));
  XOR2_X1   g212(.A(G2084), .B(G2090), .Z(new_n638));
  XNOR2_X1  g213(.A(G2067), .B(G2678), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n640), .A2(KEYINPUT17), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n638), .A2(new_n639), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n637), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(new_n611), .ZN(new_n644));
  XOR2_X1   g219(.A(G2072), .B(G2078), .Z(new_n645));
  AOI21_X1  g220(.A(new_n645), .B1(new_n640), .B2(KEYINPUT18), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(new_n619), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n644), .B(new_n647), .ZN(G227));
  XNOR2_X1  g223(.A(G1956), .B(G2474), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT77), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1961), .B(G1966), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1971), .B(G1976), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT19), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n656), .B(KEYINPUT20), .Z(new_n657));
  NOR2_X1   g232(.A1(new_n650), .A2(new_n652), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n659), .A2(new_n655), .A3(new_n653), .ZN(new_n660));
  OAI211_X1 g235(.A(new_n657), .B(new_n660), .C1(new_n655), .C2(new_n659), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1991), .B(G1996), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G1981), .B(G1986), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT78), .ZN(new_n665));
  XNOR2_X1  g240(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n663), .B(new_n667), .ZN(G229));
  INV_X1    g243(.A(G16), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n669), .A2(G21), .ZN(new_n670));
  OAI21_X1  g245(.A(new_n670), .B1(G168), .B2(new_n669), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(KEYINPUT90), .Z(new_n672));
  INV_X1    g247(.A(G1966), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n674), .B(KEYINPUT91), .Z(new_n675));
  NAND3_X1  g250(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n676));
  INV_X1    g251(.A(KEYINPUT25), .ZN(new_n677));
  OR2_X1    g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n676), .A2(new_n677), .ZN(new_n679));
  AOI22_X1  g254(.A1(new_n678), .A2(new_n679), .B1(new_n480), .B2(G139), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT85), .ZN(new_n681));
  AOI22_X1  g256(.A1(new_n607), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n682));
  OR2_X1    g257(.A1(new_n682), .A2(new_n463), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  MUX2_X1   g259(.A(G33), .B(new_n684), .S(G29), .Z(new_n685));
  NOR2_X1   g260(.A1(new_n685), .A2(G2072), .ZN(new_n686));
  AND2_X1   g261(.A1(new_n685), .A2(G2072), .ZN(new_n687));
  AOI211_X1 g262(.A(new_n686), .B(new_n687), .C1(new_n673), .C2(new_n672), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n669), .A2(G5), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n689), .B1(G171), .B2(new_n669), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(G1961), .ZN(new_n691));
  INV_X1    g266(.A(G29), .ZN(new_n692));
  INV_X1    g267(.A(G34), .ZN(new_n693));
  AND2_X1   g268(.A1(new_n693), .A2(KEYINPUT24), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n693), .A2(KEYINPUT24), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n692), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n696), .B1(G160), .B2(new_n692), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(G2084), .Z(new_n698));
  XOR2_X1   g273(.A(KEYINPUT92), .B(G28), .Z(new_n699));
  AOI21_X1  g274(.A(G29), .B1(new_n699), .B2(KEYINPUT30), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(KEYINPUT30), .B2(new_n699), .ZN(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT31), .B(G11), .ZN(new_n702));
  OAI211_X1 g277(.A(new_n701), .B(new_n702), .C1(new_n618), .C2(new_n692), .ZN(new_n703));
  NOR2_X1   g278(.A1(G27), .A2(G29), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n704), .B1(G164), .B2(G29), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n703), .B1(G2078), .B2(new_n705), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n698), .B(new_n706), .C1(G2078), .C2(new_n705), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n691), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n675), .A2(new_n688), .A3(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT27), .B(G1996), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n692), .A2(G32), .ZN(new_n712));
  NAND3_X1  g287(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT86), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(KEYINPUT26), .Z(new_n715));
  NAND2_X1  g290(.A1(new_n480), .A2(G141), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n476), .A2(G129), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n470), .A2(G105), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n716), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n715), .A2(new_n719), .ZN(new_n720));
  OR2_X1    g295(.A1(new_n720), .A2(KEYINPUT87), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n720), .A2(KEYINPUT87), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n712), .B1(new_n724), .B2(new_n692), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT88), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n709), .B1(new_n711), .B2(new_n726), .ZN(new_n727));
  OAI21_X1  g302(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n728));
  INV_X1    g303(.A(G107), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n728), .B1(new_n729), .B2(G2105), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT80), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(G131), .B2(new_n480), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n476), .A2(G119), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT79), .ZN(new_n734));
  AND2_X1   g309(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n735), .A2(G29), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G25), .B2(G29), .ZN(new_n737));
  XOR2_X1   g312(.A(KEYINPUT35), .B(G1991), .Z(new_n738));
  AND2_X1   g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n737), .A2(new_n738), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n669), .A2(G24), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(new_n581), .B2(new_n669), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(G1986), .ZN(new_n743));
  NOR3_X1   g318(.A1(new_n739), .A2(new_n740), .A3(new_n743), .ZN(new_n744));
  MUX2_X1   g319(.A(G6), .B(G305), .S(G16), .Z(new_n745));
  XOR2_X1   g320(.A(KEYINPUT32), .B(G1981), .Z(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT81), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n745), .B(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n669), .A2(G22), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G166), .B2(new_n669), .ZN(new_n750));
  INV_X1    g325(.A(G1971), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n669), .A2(G23), .ZN(new_n753));
  INV_X1    g328(.A(G288), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n753), .B1(new_n754), .B2(new_n669), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT33), .B(G1976), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT82), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n755), .B(new_n757), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n748), .A2(new_n752), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n759), .A2(KEYINPUT34), .ZN(new_n760));
  OR2_X1    g335(.A1(new_n759), .A2(KEYINPUT34), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n744), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT36), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n692), .A2(G35), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G162), .B2(new_n692), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT29), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n766), .A2(G2090), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT93), .Z(new_n768));
  NAND3_X1  g343(.A1(new_n727), .A2(new_n763), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n669), .A2(G20), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT23), .Z(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(G299), .B2(G16), .ZN(new_n772));
  INV_X1    g347(.A(G1956), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(new_n766), .B2(G2090), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT94), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n600), .A2(G16), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G4), .B2(G16), .ZN(new_n778));
  INV_X1    g353(.A(G1348), .ZN(new_n779));
  OR2_X1    g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n778), .A2(new_n779), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n669), .A2(G19), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(new_n540), .B2(new_n669), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(G1341), .Z(new_n784));
  NAND2_X1  g359(.A1(new_n692), .A2(G26), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT83), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT28), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n480), .A2(G140), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n476), .A2(G128), .ZN(new_n789));
  OR2_X1    g364(.A1(G104), .A2(G2105), .ZN(new_n790));
  OAI211_X1 g365(.A(new_n790), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n788), .A2(new_n789), .A3(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(new_n792), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n787), .B1(new_n793), .B2(new_n692), .ZN(new_n794));
  INV_X1    g369(.A(G2067), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND4_X1  g371(.A1(new_n780), .A2(new_n781), .A3(new_n784), .A4(new_n796), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT84), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n726), .A2(new_n711), .ZN(new_n799));
  AND2_X1   g374(.A1(new_n799), .A2(KEYINPUT89), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n799), .A2(KEYINPUT89), .ZN(new_n801));
  OAI211_X1 g376(.A(new_n776), .B(new_n798), .C1(new_n800), .C2(new_n801), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n769), .A2(new_n802), .ZN(G311));
  INV_X1    g378(.A(G311), .ZN(G150));
  NAND2_X1  g379(.A1(new_n600), .A2(G559), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(KEYINPUT38), .Z(new_n806));
  AOI22_X1  g381(.A1(new_n499), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n807), .A2(new_n501), .ZN(new_n808));
  XNOR2_X1  g383(.A(KEYINPUT95), .B(G93), .ZN(new_n809));
  INV_X1    g384(.A(G55), .ZN(new_n810));
  OAI22_X1  g385(.A1(new_n504), .A2(new_n809), .B1(new_n506), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n808), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n540), .A2(new_n812), .ZN(new_n813));
  OAI22_X1  g388(.A1(new_n536), .A2(new_n539), .B1(new_n808), .B2(new_n811), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n806), .B(new_n815), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n816), .A2(KEYINPUT39), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(KEYINPUT39), .ZN(new_n818));
  XOR2_X1   g393(.A(KEYINPUT96), .B(G860), .Z(new_n819));
  NAND3_X1  g394(.A1(new_n817), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n812), .A2(new_n819), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT37), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n820), .A2(new_n822), .ZN(G145));
  NAND2_X1  g398(.A1(new_n493), .A2(new_n495), .ZN(new_n824));
  AND2_X1   g399(.A1(new_n485), .A2(new_n488), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n723), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n721), .A2(G164), .A3(new_n722), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(new_n735), .ZN(new_n830));
  INV_X1    g405(.A(new_n735), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n827), .A2(new_n831), .A3(new_n828), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n480), .A2(G142), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n476), .A2(G130), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n463), .A2(G118), .ZN(new_n836));
  OAI21_X1  g411(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n837));
  OAI211_X1 g412(.A(new_n834), .B(new_n835), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT99), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(new_n609), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n684), .A2(KEYINPUT98), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT98), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n681), .A2(new_n842), .A3(new_n683), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n841), .A2(new_n793), .A3(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n793), .B1(new_n841), .B2(new_n843), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n840), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n846), .ZN(new_n848));
  INV_X1    g423(.A(new_n840), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n848), .A2(new_n844), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n833), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(G160), .B(KEYINPUT97), .ZN(new_n853));
  XNOR2_X1  g428(.A(G162), .B(new_n853), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n854), .B(new_n618), .Z(new_n855));
  NAND4_X1  g430(.A1(new_n830), .A2(new_n847), .A3(new_n850), .A4(new_n832), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n852), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  XOR2_X1   g432(.A(new_n857), .B(KEYINPUT102), .Z(new_n858));
  AOI211_X1 g433(.A(KEYINPUT100), .B(new_n855), .C1(new_n856), .C2(new_n852), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT100), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n852), .A2(new_n856), .ZN(new_n861));
  INV_X1    g436(.A(new_n855), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n860), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  OR2_X1    g438(.A1(new_n859), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(KEYINPUT101), .B(G37), .ZN(new_n865));
  NAND4_X1  g440(.A1(new_n858), .A2(new_n864), .A3(KEYINPUT40), .A4(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT40), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n865), .B1(new_n859), .B2(new_n863), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n857), .B(KEYINPUT102), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n867), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  AND2_X1   g445(.A1(new_n866), .A2(new_n870), .ZN(G395));
  INV_X1    g446(.A(G868), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n872), .B1(new_n808), .B2(new_n811), .ZN(new_n873));
  AND2_X1   g448(.A1(new_n813), .A2(new_n814), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n604), .B(new_n874), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n596), .A2(new_n589), .A3(new_n591), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n596), .B1(new_n589), .B2(new_n591), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n875), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n592), .A2(G299), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT41), .ZN(new_n882));
  AND3_X1   g457(.A1(new_n881), .A2(new_n882), .A3(new_n876), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n882), .B1(new_n881), .B2(new_n876), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n880), .B1(new_n885), .B2(new_n875), .ZN(new_n886));
  XNOR2_X1  g461(.A(G166), .B(G288), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n581), .B(G305), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n887), .B(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(KEYINPUT42), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n886), .B(new_n890), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n873), .B1(new_n891), .B2(new_n872), .ZN(G295));
  OAI21_X1  g467(.A(new_n873), .B1(new_n891), .B2(new_n872), .ZN(G331));
  INV_X1    g468(.A(KEYINPUT43), .ZN(new_n894));
  AOI21_X1  g469(.A(G286), .B1(new_n526), .B2(new_n533), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n526), .A2(new_n533), .A3(G286), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n874), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT103), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n897), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n815), .B1(new_n901), .B2(new_n895), .ZN(new_n902));
  NAND4_X1  g477(.A1(new_n874), .A2(new_n896), .A3(KEYINPUT103), .A4(new_n897), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n900), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(KEYINPUT41), .B1(new_n877), .B2(new_n878), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n881), .A2(new_n882), .A3(new_n876), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n905), .A2(KEYINPUT104), .A3(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT104), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n884), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n904), .A2(new_n907), .A3(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n879), .A2(new_n902), .A3(new_n898), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n889), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n900), .A2(new_n903), .A3(new_n879), .A4(new_n902), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n898), .A2(new_n902), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n916), .B1(new_n883), .B2(new_n884), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n915), .A2(new_n917), .A3(new_n889), .ZN(new_n918));
  AND2_X1   g493(.A1(new_n918), .A2(new_n865), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT105), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n914), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n889), .B1(new_n910), .B2(new_n911), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n918), .A2(new_n865), .ZN(new_n923));
  OAI21_X1  g498(.A(KEYINPUT105), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n894), .B1(new_n921), .B2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(G37), .ZN(new_n926));
  AND2_X1   g501(.A1(new_n918), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n915), .A2(new_n917), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(new_n913), .ZN(new_n929));
  AOI21_X1  g504(.A(KEYINPUT43), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g505(.A(KEYINPUT44), .B1(new_n925), .B2(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n914), .A2(new_n919), .A3(new_n894), .ZN(new_n932));
  AND2_X1   g507(.A1(new_n927), .A2(new_n929), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n932), .B1(new_n933), .B2(new_n894), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT106), .ZN(new_n937));
  AND3_X1   g512(.A1(new_n931), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n937), .B1(new_n931), .B2(new_n936), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n938), .A2(new_n939), .ZN(G397));
  AOI21_X1  g515(.A(G1384), .B1(new_n824), .B2(new_n825), .ZN(new_n941));
  OAI21_X1  g516(.A(KEYINPUT110), .B1(new_n941), .B2(KEYINPUT45), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n466), .A2(new_n467), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(G2105), .ZN(new_n944));
  AND2_X1   g519(.A1(new_n469), .A2(new_n471), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n944), .A2(new_n945), .A3(G40), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n946), .B1(new_n941), .B2(KEYINPUT45), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT110), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT45), .ZN(new_n949));
  OAI211_X1 g524(.A(new_n948), .B(new_n949), .C1(G164), .C2(G1384), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n942), .A2(new_n947), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(KEYINPUT111), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT111), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n942), .A2(new_n947), .A3(new_n953), .A4(new_n950), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n952), .A2(new_n751), .A3(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT112), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n952), .A2(KEYINPUT112), .A3(new_n751), .A4(new_n954), .ZN(new_n958));
  INV_X1    g533(.A(G40), .ZN(new_n959));
  NOR3_X1   g534(.A1(new_n468), .A2(new_n472), .A3(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT50), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n960), .B1(new_n941), .B2(new_n961), .ZN(new_n962));
  NOR3_X1   g537(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(G2090), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n957), .A2(new_n958), .A3(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(G8), .ZN(new_n968));
  NOR2_X1   g543(.A1(G166), .A2(new_n968), .ZN(new_n969));
  XNOR2_X1  g544(.A(KEYINPUT113), .B(KEYINPUT55), .ZN(new_n970));
  OR2_X1    g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT113), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n969), .B1(new_n972), .B2(KEYINPUT55), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n968), .B1(new_n941), .B2(new_n960), .ZN(new_n975));
  INV_X1    g550(.A(G1981), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n976), .B1(new_n574), .B2(KEYINPUT114), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(G305), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n568), .B(new_n574), .C1(KEYINPUT114), .C2(new_n976), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT49), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n975), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n980), .A2(new_n981), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT115), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n980), .A2(KEYINPUT115), .A3(new_n981), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n982), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n754), .A2(G1976), .ZN(new_n988));
  INV_X1    g563(.A(G1976), .ZN(new_n989));
  AOI21_X1  g564(.A(KEYINPUT52), .B1(G288), .B2(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n975), .A2(new_n988), .A3(new_n990), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n975), .A2(new_n988), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT52), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n991), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n987), .A2(new_n994), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n967), .A2(G8), .A3(new_n974), .A4(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n754), .A2(new_n989), .ZN(new_n997));
  OAI22_X1  g572(.A1(new_n987), .A2(new_n997), .B1(G1981), .B2(G305), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(new_n975), .ZN(new_n999));
  AND2_X1   g574(.A1(new_n996), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(G286), .A2(G8), .ZN(new_n1001));
  XOR2_X1   g576(.A(new_n1001), .B(KEYINPUT122), .Z(new_n1002));
  OAI21_X1  g577(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1003));
  INV_X1    g578(.A(G1384), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n826), .A2(new_n961), .A3(new_n1004), .ZN(new_n1005));
  XOR2_X1   g580(.A(KEYINPUT118), .B(G2084), .Z(new_n1006));
  NAND4_X1  g581(.A1(new_n1003), .A2(new_n1005), .A3(new_n960), .A4(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n949), .B1(G164), .B2(G1384), .ZN(new_n1009));
  AOI21_X1  g584(.A(G1966), .B1(new_n947), .B2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1002), .A2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(G8), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1013));
  AOI21_X1  g588(.A(KEYINPUT123), .B1(new_n1013), .B2(new_n1002), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT51), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1012), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT123), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n826), .A2(KEYINPUT45), .A3(new_n1004), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1009), .A2(new_n960), .A3(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(new_n673), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n968), .B1(new_n1020), .B2(new_n1007), .ZN(new_n1021));
  XNOR2_X1  g596(.A(new_n1001), .B(KEYINPUT122), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1017), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1013), .A2(new_n1002), .A3(KEYINPUT123), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1023), .A2(KEYINPUT51), .A3(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(G2078), .B1(new_n952), .B2(new_n954), .ZN(new_n1026));
  OR2_X1    g601(.A1(new_n1026), .A2(KEYINPUT53), .ZN(new_n1027));
  OAI21_X1  g602(.A(KEYINPUT121), .B1(new_n962), .B2(new_n963), .ZN(new_n1028));
  INV_X1    g603(.A(G1961), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT121), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1003), .A2(new_n1005), .A3(new_n1030), .A4(new_n960), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1028), .A2(new_n1029), .A3(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(KEYINPUT125), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT125), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1028), .A2(new_n1034), .A3(new_n1029), .A4(new_n1031), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT54), .ZN(new_n1036));
  NAND2_X1  g611(.A1(G171), .A2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n526), .A2(new_n533), .A3(KEYINPUT54), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(G2078), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1009), .A2(KEYINPUT53), .A3(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n960), .A2(KEYINPUT126), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT126), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n946), .A2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1018), .A2(new_n1042), .A3(new_n1044), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1041), .A2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1039), .A2(new_n1046), .ZN(new_n1047));
  AND3_X1   g622(.A1(new_n1033), .A2(new_n1035), .A3(new_n1047), .ZN(new_n1048));
  AOI22_X1  g623(.A1(new_n1016), .A2(new_n1025), .B1(new_n1027), .B2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n967), .A2(G8), .A3(new_n974), .ZN(new_n1050));
  OAI211_X1 g625(.A(KEYINPUT116), .B(new_n960), .C1(new_n941), .C2(new_n961), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(new_n1005), .ZN(new_n1052));
  AOI21_X1  g627(.A(KEYINPUT116), .B1(new_n1003), .B2(new_n960), .ZN(new_n1053));
  OR3_X1    g628(.A1(new_n1052), .A2(new_n1053), .A3(G2090), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n955), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(G8), .ZN(new_n1056));
  INV_X1    g631(.A(new_n974), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT117), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1058), .B1(new_n987), .B2(new_n994), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n993), .B1(new_n975), .B2(new_n988), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1060), .B1(new_n992), .B2(new_n990), .ZN(new_n1061));
  AOI21_X1  g636(.A(KEYINPUT115), .B1(new_n980), .B2(new_n981), .ZN(new_n1062));
  AOI211_X1 g637(.A(new_n984), .B(KEYINPUT49), .C1(new_n978), .C2(new_n979), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n1061), .B(KEYINPUT117), .C1(new_n1064), .C2(new_n982), .ZN(new_n1065));
  AOI22_X1  g640(.A1(new_n1056), .A2(new_n1057), .B1(new_n1059), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT124), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n947), .A2(KEYINPUT53), .A3(new_n1040), .A4(new_n1009), .ZN(new_n1068));
  AND3_X1   g643(.A1(new_n1032), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1067), .B1(new_n1032), .B2(new_n1068), .ZN(new_n1070));
  OAI22_X1  g645(.A1(new_n1069), .A2(new_n1070), .B1(KEYINPUT53), .B2(new_n1026), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(new_n1039), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1049), .A2(new_n1050), .A3(new_n1066), .A4(new_n1072), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n773), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT119), .ZN(new_n1075));
  AOI21_X1  g650(.A(KEYINPUT57), .B1(new_n553), .B2(new_n1075), .ZN(new_n1076));
  XNOR2_X1  g651(.A(new_n1076), .B(G299), .ZN(new_n1077));
  XNOR2_X1  g652(.A(KEYINPUT56), .B(G2072), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n942), .A2(new_n947), .A3(new_n950), .A4(new_n1078), .ZN(new_n1079));
  AND3_X1   g654(.A1(new_n1074), .A2(new_n1077), .A3(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1028), .A2(new_n779), .A3(new_n1031), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT120), .ZN(new_n1082));
  INV_X1    g657(.A(new_n495), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n494), .B1(new_n607), .B2(new_n491), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1004), .B1(new_n1085), .B2(new_n489), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1082), .B1(new_n1086), .B2(new_n946), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n941), .A2(new_n960), .A3(KEYINPUT120), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(new_n795), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1081), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(new_n600), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1074), .A2(new_n1079), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1077), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1080), .B1(new_n1092), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT61), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1077), .B1(new_n1074), .B2(new_n1079), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1097), .B1(new_n1080), .B2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1074), .A2(new_n1077), .A3(new_n1079), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1095), .A2(KEYINPUT61), .A3(new_n1100), .ZN(new_n1101));
  AND2_X1   g676(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1081), .A2(KEYINPUT60), .A3(new_n1090), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(new_n600), .ZN(new_n1104));
  AOI21_X1  g679(.A(KEYINPUT60), .B1(new_n1081), .B2(new_n1090), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(G1996), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n942), .A2(new_n947), .A3(new_n1107), .A4(new_n950), .ZN(new_n1108));
  XOR2_X1   g683(.A(KEYINPUT58), .B(G1341), .Z(new_n1109));
  NAND3_X1  g684(.A1(new_n1087), .A2(new_n1088), .A3(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(new_n540), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT59), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1081), .A2(KEYINPUT60), .A3(new_n592), .A4(new_n1090), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1111), .A2(KEYINPUT59), .A3(new_n540), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1114), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1106), .A2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1096), .B1(new_n1102), .B2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1000), .B1(new_n1073), .B2(new_n1119), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1013), .A2(G286), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1066), .A2(new_n1050), .A3(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT63), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n995), .A2(KEYINPUT63), .A3(new_n1121), .ZN(new_n1124));
  AOI22_X1  g699(.A1(new_n955), .A2(new_n956), .B1(new_n965), .B2(new_n964), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n968), .B1(new_n1125), .B2(new_n958), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1124), .B1(new_n1126), .B2(new_n974), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n967), .A2(G8), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(new_n1057), .ZN(new_n1129));
  AOI22_X1  g704(.A1(new_n1122), .A2(new_n1123), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(KEYINPUT127), .B1(new_n1120), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1016), .A2(new_n1025), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1027), .A2(new_n1048), .ZN(new_n1136));
  AND3_X1   g711(.A1(new_n1135), .A2(new_n1072), .A3(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1096), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT60), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1091), .A2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1140), .A2(new_n600), .A3(new_n1103), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1141), .A2(new_n1115), .A3(new_n1116), .A4(new_n1114), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1138), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  AND2_X1   g719(.A1(new_n1066), .A2(new_n1050), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1137), .A2(new_n1144), .A3(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT127), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1134), .A2(new_n1146), .A3(new_n1147), .A4(new_n1000), .ZN(new_n1148));
  XOR2_X1   g723(.A(new_n1135), .B(KEYINPUT62), .Z(new_n1149));
  NAND4_X1  g724(.A1(new_n1149), .A2(G171), .A3(new_n1145), .A4(new_n1071), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1131), .A2(new_n1148), .A3(new_n1150), .ZN(new_n1151));
  OR3_X1    g726(.A1(new_n1009), .A2(KEYINPUT107), .A3(new_n946), .ZN(new_n1152));
  OAI21_X1  g727(.A(KEYINPUT107), .B1(new_n1009), .B2(new_n946), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1154), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n724), .A2(new_n1107), .ZN(new_n1156));
  XNOR2_X1  g731(.A(new_n792), .B(G2067), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1155), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n724), .A2(new_n1155), .A3(new_n1107), .ZN(new_n1159));
  AND2_X1   g734(.A1(new_n1159), .A2(KEYINPUT108), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1159), .A2(KEYINPUT108), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1158), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT109), .ZN(new_n1163));
  XNOR2_X1  g738(.A(new_n1162), .B(new_n1163), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n735), .A2(new_n738), .ZN(new_n1165));
  AND2_X1   g740(.A1(new_n735), .A2(new_n738), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1155), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1164), .A2(new_n1167), .ZN(new_n1168));
  XOR2_X1   g743(.A(new_n581), .B(G1986), .Z(new_n1169));
  AOI21_X1  g744(.A(new_n1168), .B1(new_n1155), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1151), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1155), .A2(new_n1107), .ZN(new_n1172));
  XNOR2_X1  g747(.A(new_n1172), .B(KEYINPUT46), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1155), .B1(new_n723), .B2(new_n1157), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  XNOR2_X1  g750(.A(new_n1175), .B(KEYINPUT47), .ZN(new_n1176));
  NOR3_X1   g751(.A1(new_n1154), .A2(G1986), .A3(G290), .ZN(new_n1177));
  XNOR2_X1  g752(.A(new_n1177), .B(KEYINPUT48), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1176), .B1(new_n1168), .B2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n793), .A2(new_n795), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1154), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1179), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1171), .A2(new_n1183), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g759(.A1(new_n858), .A2(new_n864), .A3(new_n865), .ZN(new_n1186));
  NOR4_X1   g760(.A1(G229), .A2(new_n461), .A3(G401), .A4(G227), .ZN(new_n1187));
  AND3_X1   g761(.A1(new_n1186), .A2(new_n934), .A3(new_n1187), .ZN(G308));
  NAND3_X1  g762(.A1(new_n1186), .A2(new_n934), .A3(new_n1187), .ZN(G225));
endmodule


