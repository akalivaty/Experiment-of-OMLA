//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 1 0 1 1 0 0 0 0 1 1 0 0 0 0 1 0 0 0 0 1 1 1 1 1 1 1 0 0 0 0 1 0 0 1 0 1 0 1 1 0 0 1 0 1 0 1 1 0 1 1 0 0 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:50 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n713,
    new_n714, new_n715, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n972, new_n973, new_n974, new_n975, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020;
  INV_X1    g000(.A(G224), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(G953), .ZN(new_n188));
  AND2_X1   g002(.A1(KEYINPUT0), .A2(G128), .ZN(new_n189));
  NOR2_X1   g003(.A1(KEYINPUT0), .A2(G128), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT64), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(KEYINPUT64), .A2(G146), .ZN(new_n195));
  AOI21_X1  g009(.A(G143), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G143), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n197), .A2(G146), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n191), .B1(new_n196), .B2(new_n198), .ZN(new_n199));
  OAI21_X1  g013(.A(KEYINPUT65), .B1(new_n193), .B2(G143), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT65), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n201), .A2(new_n197), .A3(G146), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n194), .A2(G143), .A3(new_n195), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n203), .A2(new_n204), .A3(new_n189), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n199), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT72), .ZN(new_n207));
  INV_X1    g021(.A(G125), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(KEYINPUT72), .A2(G125), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n206), .A2(KEYINPUT88), .A3(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G128), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n213), .A2(KEYINPUT1), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n203), .A2(new_n204), .A3(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(new_n211), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n213), .B1(new_n204), .B2(KEYINPUT1), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n196), .A2(new_n198), .ZN(new_n218));
  OAI211_X1 g032(.A(new_n215), .B(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n212), .A2(new_n219), .ZN(new_n220));
  AOI21_X1  g034(.A(KEYINPUT88), .B1(new_n206), .B2(new_n211), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n188), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(new_n221), .ZN(new_n223));
  INV_X1    g037(.A(new_n188), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n223), .A2(new_n224), .A3(new_n219), .A4(new_n212), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n222), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G104), .ZN(new_n227));
  OAI21_X1  g041(.A(KEYINPUT3), .B1(new_n227), .B2(G107), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n229));
  INV_X1    g043(.A(G107), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n229), .A2(new_n230), .A3(G104), .ZN(new_n231));
  AND2_X1   g045(.A1(new_n228), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G101), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(KEYINPUT82), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT82), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G101), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n227), .A2(G107), .ZN(new_n237));
  AND3_X1   g051(.A1(new_n234), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT83), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n232), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n228), .A2(new_n231), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n234), .A2(new_n236), .A3(new_n237), .ZN(new_n242));
  OAI21_X1  g056(.A(KEYINPUT83), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n240), .A2(new_n243), .ZN(new_n244));
  XOR2_X1   g058(.A(KEYINPUT2), .B(G113), .Z(new_n245));
  INV_X1    g059(.A(G119), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(KEYINPUT67), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT67), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G119), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n247), .A2(new_n249), .A3(G116), .ZN(new_n250));
  INV_X1    g064(.A(G116), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G119), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n245), .A2(new_n250), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n230), .A2(G104), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(new_n237), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G101), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n250), .A2(KEYINPUT5), .A3(new_n252), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT5), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n247), .A2(new_n249), .A3(new_n258), .A4(G116), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n257), .A2(G113), .A3(new_n259), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n244), .A2(new_n253), .A3(new_n256), .A4(new_n260), .ZN(new_n261));
  XOR2_X1   g075(.A(G110), .B(G122), .Z(new_n262));
  XNOR2_X1  g076(.A(new_n262), .B(KEYINPUT86), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n228), .A2(new_n231), .A3(new_n237), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G101), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(KEYINPUT4), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n266), .B1(new_n240), .B2(new_n243), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT4), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n264), .A2(new_n268), .A3(G101), .ZN(new_n269));
  INV_X1    g083(.A(new_n253), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n245), .B1(new_n250), .B2(new_n252), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n269), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n261), .B(new_n263), .C1(new_n267), .C2(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n239), .B1(new_n232), .B2(new_n238), .ZN(new_n274));
  NOR3_X1   g088(.A1(new_n241), .A2(new_n242), .A3(KEYINPUT83), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n256), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n260), .A2(new_n253), .ZN(new_n277));
  OAI22_X1  g091(.A1(new_n267), .A2(new_n272), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n263), .B(KEYINPUT87), .ZN(new_n279));
  AOI22_X1  g093(.A1(new_n273), .A2(KEYINPUT6), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  AND3_X1   g094(.A1(new_n278), .A2(KEYINPUT6), .A3(new_n279), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n226), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(G902), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n244), .A2(new_n253), .A3(new_n256), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT89), .ZN(new_n285));
  AND3_X1   g099(.A1(new_n259), .A2(new_n285), .A3(G113), .ZN(new_n286));
  INV_X1    g100(.A(new_n257), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n285), .B1(new_n259), .B2(G113), .ZN(new_n288));
  NOR3_X1   g102(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  AND2_X1   g103(.A1(new_n259), .A2(G113), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n270), .B1(new_n257), .B2(new_n290), .ZN(new_n291));
  AOI22_X1  g105(.A1(new_n240), .A2(new_n243), .B1(G101), .B2(new_n255), .ZN(new_n292));
  OAI22_X1  g106(.A1(new_n284), .A2(new_n289), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  XNOR2_X1  g107(.A(new_n263), .B(KEYINPUT8), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT7), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n188), .A2(new_n296), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n223), .A2(new_n219), .A3(new_n212), .A4(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n206), .A2(new_n211), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(new_n219), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n300), .B1(new_n296), .B2(new_n188), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n295), .A2(new_n273), .A3(new_n298), .A4(new_n301), .ZN(new_n302));
  OAI21_X1  g116(.A(G210), .B1(G237), .B2(G902), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n282), .A2(new_n283), .A3(new_n302), .A4(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT90), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  AND2_X1   g120(.A1(new_n302), .A2(new_n283), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n307), .A2(KEYINPUT90), .A3(new_n282), .A4(new_n303), .ZN(new_n308));
  INV_X1    g122(.A(new_n303), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n273), .A2(KEYINPUT6), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n278), .A2(new_n279), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n278), .A2(KEYINPUT6), .A3(new_n279), .ZN(new_n313));
  AOI22_X1  g127(.A1(new_n312), .A2(new_n313), .B1(new_n222), .B2(new_n225), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n302), .A2(new_n283), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n309), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n306), .A2(new_n308), .A3(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(G214), .B1(G237), .B2(G902), .ZN(new_n318));
  XNOR2_X1  g132(.A(new_n318), .B(KEYINPUT85), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n317), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  XNOR2_X1  g136(.A(KEYINPUT9), .B(G234), .ZN(new_n323));
  OAI21_X1  g137(.A(G221), .B1(new_n323), .B2(G902), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(G469), .ZN(new_n326));
  INV_X1    g140(.A(G953), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G227), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n328), .B(KEYINPUT80), .ZN(new_n329));
  XOR2_X1   g143(.A(G110), .B(G140), .Z(new_n330));
  XNOR2_X1  g144(.A(new_n329), .B(new_n330), .ZN(new_n331));
  AND2_X1   g145(.A1(KEYINPUT64), .A2(G146), .ZN(new_n332));
  NOR2_X1   g146(.A1(KEYINPUT64), .A2(G146), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AOI22_X1  g148(.A1(new_n334), .A2(G143), .B1(new_n200), .B2(new_n202), .ZN(new_n335));
  INV_X1    g149(.A(new_n198), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n213), .B1(new_n336), .B2(KEYINPUT1), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n215), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n244), .A2(new_n338), .A3(new_n256), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT10), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  AND3_X1   g155(.A1(new_n199), .A2(new_n269), .A3(new_n205), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n274), .A2(new_n275), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n342), .B1(new_n343), .B2(new_n266), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT11), .ZN(new_n345));
  INV_X1    g159(.A(G134), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n345), .B1(new_n346), .B2(G137), .ZN(new_n347));
  INV_X1    g161(.A(G137), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n348), .A2(KEYINPUT11), .A3(G134), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n346), .A2(G137), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n347), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(G131), .ZN(new_n352));
  INV_X1    g166(.A(G131), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n347), .A2(new_n349), .A3(new_n353), .A4(new_n350), .ZN(new_n354));
  AND2_X1   g168(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n215), .B1(new_n217), .B2(new_n218), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n292), .A2(KEYINPUT10), .A3(new_n356), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n341), .A2(new_n344), .A3(new_n355), .A4(new_n357), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n339), .B1(new_n356), .B2(new_n292), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n352), .A2(new_n354), .ZN(new_n360));
  AND3_X1   g174(.A1(new_n359), .A2(KEYINPUT12), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(KEYINPUT12), .B1(new_n359), .B2(new_n360), .ZN(new_n362));
  OAI211_X1 g176(.A(new_n331), .B(new_n358), .C1(new_n361), .C2(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n341), .A2(new_n344), .A3(new_n357), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(new_n360), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n331), .B1(new_n365), .B2(new_n358), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT84), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n363), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  AOI211_X1 g182(.A(KEYINPUT84), .B(new_n331), .C1(new_n365), .C2(new_n358), .ZN(new_n369));
  OAI211_X1 g183(.A(new_n326), .B(new_n283), .C1(new_n368), .C2(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n358), .B1(new_n361), .B2(new_n362), .ZN(new_n371));
  XNOR2_X1  g185(.A(new_n331), .B(KEYINPUT81), .ZN(new_n372));
  AND2_X1   g186(.A1(new_n358), .A2(new_n331), .ZN(new_n373));
  AOI22_X1  g187(.A1(new_n371), .A2(new_n372), .B1(new_n365), .B2(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(G469), .B1(new_n374), .B2(G902), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n325), .B1(new_n370), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(KEYINPUT18), .A2(G131), .ZN(new_n377));
  INV_X1    g191(.A(G237), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n378), .A2(new_n327), .A3(G214), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(new_n197), .ZN(new_n380));
  NOR2_X1   g194(.A1(G237), .A2(G953), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n381), .A2(G143), .A3(G214), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT92), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n377), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n380), .A2(KEYINPUT92), .A3(new_n382), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  OR2_X1    g201(.A1(KEYINPUT71), .A2(G140), .ZN(new_n388));
  NAND2_X1  g202(.A1(KEYINPUT71), .A2(G140), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n388), .A2(G125), .A3(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n209), .A2(G140), .A3(new_n210), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  OAI21_X1  g207(.A(G146), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  XNOR2_X1  g208(.A(G125), .B(G140), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n334), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(new_n382), .ZN(new_n398));
  AOI21_X1  g212(.A(G143), .B1(new_n381), .B2(G214), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n377), .B(KEYINPUT93), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n387), .A2(new_n397), .A3(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(KEYINPUT19), .B1(new_n391), .B2(new_n393), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT19), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n395), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n404), .A2(new_n334), .A3(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n390), .A2(new_n392), .A3(KEYINPUT16), .ZN(new_n408));
  NOR2_X1   g222(.A1(KEYINPUT16), .A2(G140), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n211), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n408), .A2(G146), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n407), .A2(new_n411), .ZN(new_n412));
  OAI21_X1  g226(.A(G131), .B1(new_n398), .B2(new_n399), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT94), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n400), .A2(new_n353), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n383), .A2(KEYINPUT94), .A3(G131), .ZN(new_n417));
  AND3_X1   g231(.A1(new_n415), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n403), .B1(new_n412), .B2(new_n418), .ZN(new_n419));
  XNOR2_X1  g233(.A(G113), .B(G122), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n420), .B(new_n227), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT17), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n415), .A2(new_n416), .A3(new_n424), .A4(new_n417), .ZN(new_n425));
  AOI21_X1  g239(.A(KEYINPUT94), .B1(new_n383), .B2(G131), .ZN(new_n426));
  AOI211_X1 g240(.A(new_n414), .B(new_n353), .C1(new_n380), .C2(new_n382), .ZN(new_n427));
  OAI21_X1  g241(.A(KEYINPUT17), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n425), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n411), .A2(KEYINPUT73), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n408), .A2(new_n410), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n193), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT73), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n408), .A2(new_n433), .A3(G146), .A4(new_n410), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n430), .A2(new_n432), .A3(new_n434), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n421), .B(new_n403), .C1(new_n429), .C2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n423), .A2(new_n436), .ZN(new_n437));
  NOR2_X1   g251(.A1(G475), .A2(G902), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n438), .B(KEYINPUT95), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n437), .A2(new_n440), .ZN(new_n441));
  XOR2_X1   g255(.A(KEYINPUT91), .B(KEYINPUT20), .Z(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT20), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n437), .A2(new_n445), .A3(new_n440), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n403), .B1(new_n429), .B2(new_n435), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(new_n422), .ZN(new_n448));
  AOI21_X1  g262(.A(G902), .B1(new_n448), .B2(new_n436), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  AOI22_X1  g264(.A1(new_n444), .A2(new_n446), .B1(new_n450), .B2(G475), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT98), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n197), .A2(G128), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n213), .A2(G143), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n453), .A2(new_n454), .A3(new_n346), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n346), .B1(new_n453), .B2(new_n454), .ZN(new_n457));
  XOR2_X1   g271(.A(G116), .B(G122), .Z(new_n458));
  OAI22_X1  g272(.A1(new_n456), .A2(new_n457), .B1(G107), .B2(new_n458), .ZN(new_n459));
  XNOR2_X1  g273(.A(G116), .B(G122), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT14), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(G122), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n463), .A2(G116), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n230), .B1(new_n464), .B2(KEYINPUT14), .ZN(new_n465));
  AOI21_X1  g279(.A(KEYINPUT96), .B1(new_n462), .B2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n462), .A2(KEYINPUT96), .A3(new_n465), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n459), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n458), .A2(G107), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n460), .A2(new_n230), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n455), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n197), .A2(G128), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT13), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n473), .B1(new_n474), .B2(new_n453), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n197), .A2(KEYINPUT13), .A3(G128), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n346), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n472), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(G217), .ZN(new_n479));
  NOR3_X1   g293(.A1(new_n323), .A2(new_n479), .A3(G953), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  NOR3_X1   g295(.A1(new_n469), .A2(new_n478), .A3(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n459), .ZN(new_n483));
  INV_X1    g297(.A(new_n468), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n483), .B1(new_n484), .B2(new_n466), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n475), .A2(new_n476), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(G134), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n487), .B(new_n455), .C1(new_n471), .C2(new_n470), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n480), .B1(new_n485), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n283), .B1(new_n482), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(KEYINPUT97), .ZN(new_n491));
  INV_X1    g305(.A(G478), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n492), .A2(KEYINPUT15), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT97), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n494), .B(new_n283), .C1(new_n482), .C2(new_n489), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n491), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  OR2_X1    g310(.A1(new_n490), .A2(new_n493), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(G234), .A2(G237), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n500), .A2(G952), .A3(new_n327), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n500), .A2(G902), .A3(G953), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  XNOR2_X1  g318(.A(KEYINPUT21), .B(G898), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n502), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n451), .A2(new_n452), .A3(new_n499), .A4(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n442), .B1(new_n437), .B2(new_n440), .ZN(new_n509));
  AOI211_X1 g323(.A(KEYINPUT20), .B(new_n439), .C1(new_n423), .C2(new_n436), .ZN(new_n510));
  INV_X1    g324(.A(G475), .ZN(new_n511));
  OAI22_X1  g325(.A1(new_n509), .A2(new_n510), .B1(new_n511), .B2(new_n449), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n496), .A2(new_n497), .A3(new_n507), .ZN(new_n513));
  OAI21_X1  g327(.A(KEYINPUT98), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n508), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n322), .A2(new_n376), .A3(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT28), .ZN(new_n518));
  OAI21_X1  g332(.A(KEYINPUT68), .B1(new_n355), .B2(new_n206), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT68), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n360), .A2(new_n520), .A3(new_n199), .A4(new_n205), .ZN(new_n521));
  INV_X1    g335(.A(new_n350), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n346), .A2(G137), .ZN(new_n523));
  OAI21_X1  g337(.A(G131), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  AND2_X1   g338(.A1(new_n524), .A2(new_n354), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n356), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n519), .A2(new_n521), .A3(new_n526), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n270), .A2(new_n271), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n519), .A2(new_n526), .A3(new_n528), .A4(new_n521), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n518), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n355), .A2(new_n206), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(KEYINPUT28), .B1(new_n534), .B2(new_n526), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  XOR2_X1   g350(.A(KEYINPUT26), .B(G101), .Z(new_n537));
  NAND2_X1  g351(.A1(new_n381), .A2(G210), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n537), .B(new_n538), .ZN(new_n539));
  XNOR2_X1  g353(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n539), .B(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n536), .A2(KEYINPUT29), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n283), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT66), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n545), .B1(new_n355), .B2(new_n206), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n360), .A2(KEYINPUT66), .A3(new_n199), .A4(new_n205), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n546), .A2(new_n526), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(new_n529), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n518), .B1(new_n549), .B2(new_n531), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n542), .B1(new_n550), .B2(new_n535), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT30), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n548), .A2(new_n552), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n519), .A2(new_n526), .A3(KEYINPUT30), .A4(new_n521), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n553), .A2(new_n529), .A3(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n555), .A2(new_n531), .A3(new_n541), .ZN(new_n556));
  AOI21_X1  g370(.A(KEYINPUT29), .B1(new_n551), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(G472), .B1(new_n544), .B2(new_n557), .ZN(new_n558));
  AND2_X1   g372(.A1(new_n542), .A2(new_n531), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n555), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(KEYINPUT31), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n541), .B1(new_n550), .B2(new_n535), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT31), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n555), .A2(new_n563), .A3(new_n559), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n561), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT32), .ZN(new_n566));
  NOR2_X1   g380(.A1(G472), .A2(G902), .ZN(new_n567));
  AND3_X1   g381(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n566), .B1(new_n565), .B2(new_n567), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n558), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT23), .ZN(new_n571));
  XNOR2_X1  g385(.A(KEYINPUT67), .B(G119), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n571), .B1(new_n572), .B2(G128), .ZN(new_n573));
  XNOR2_X1  g387(.A(KEYINPUT74), .B(G110), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n246), .A2(G128), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n575), .B1(new_n572), .B2(G128), .ZN(new_n576));
  OAI211_X1 g390(.A(new_n573), .B(new_n574), .C1(new_n576), .C2(new_n571), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(KEYINPUT75), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n247), .A2(new_n249), .A3(G128), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n579), .B1(new_n246), .B2(G128), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(KEYINPUT23), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT75), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n581), .A2(new_n582), .A3(new_n573), .A4(new_n574), .ZN(new_n583));
  XOR2_X1   g397(.A(KEYINPUT24), .B(G110), .Z(new_n584));
  OR2_X1    g398(.A1(new_n576), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n578), .A2(new_n583), .A3(new_n585), .ZN(new_n586));
  AND2_X1   g400(.A1(new_n411), .A2(new_n396), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n573), .B1(new_n576), .B2(new_n571), .ZN(new_n589));
  AOI22_X1  g403(.A1(new_n589), .A2(G110), .B1(new_n576), .B2(new_n584), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n435), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT77), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n327), .A2(G221), .A3(G234), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n594), .B(KEYINPUT76), .ZN(new_n595));
  XNOR2_X1  g409(.A(KEYINPUT22), .B(G137), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n595), .B(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n592), .A2(new_n593), .A3(new_n597), .ZN(new_n598));
  AOI22_X1  g412(.A1(new_n586), .A2(new_n587), .B1(new_n435), .B2(new_n590), .ZN(new_n599));
  INV_X1    g413(.A(new_n597), .ZN(new_n600));
  OAI21_X1  g414(.A(KEYINPUT77), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  AOI22_X1  g415(.A1(new_n598), .A2(new_n601), .B1(new_n599), .B2(new_n600), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(G234), .ZN(new_n604));
  AOI21_X1  g418(.A(G902), .B1(new_n604), .B2(G217), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n605), .B(KEYINPUT79), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(G902), .B1(new_n599), .B2(new_n600), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n593), .B1(new_n592), .B2(new_n597), .ZN(new_n609));
  NOR3_X1   g423(.A1(new_n599), .A2(KEYINPUT77), .A3(new_n600), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n608), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT25), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n598), .A2(new_n601), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n614), .A2(KEYINPUT25), .A3(new_n608), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n613), .A2(KEYINPUT78), .A3(new_n615), .ZN(new_n616));
  OAI21_X1  g430(.A(G217), .B1(new_n604), .B2(G902), .ZN(new_n617));
  XOR2_X1   g431(.A(new_n617), .B(KEYINPUT70), .Z(new_n618));
  AOI21_X1  g432(.A(KEYINPUT25), .B1(new_n614), .B2(new_n608), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT78), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n607), .B1(new_n616), .B2(new_n621), .ZN(new_n622));
  AND2_X1   g436(.A1(new_n570), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n517), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n234), .A2(new_n236), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(G3));
  NAND2_X1  g440(.A1(new_n565), .A2(new_n283), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(G472), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n565), .A2(new_n567), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  AND3_X1   g445(.A1(new_n631), .A2(new_n622), .A3(new_n376), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n492), .A2(G902), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n481), .B1(new_n469), .B2(new_n478), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n485), .A2(new_n488), .A3(new_n480), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT33), .ZN(new_n636));
  AND3_X1   g450(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n636), .B1(new_n634), .B2(new_n635), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n633), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(KEYINPUT100), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n491), .A2(new_n492), .A3(new_n495), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT100), .ZN(new_n642));
  OAI211_X1 g456(.A(new_n642), .B(new_n633), .C1(new_n637), .C2(new_n638), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n640), .A2(new_n641), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n512), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n304), .A2(KEYINPUT99), .A3(new_n320), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n646), .A2(new_n320), .A3(new_n316), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n307), .A2(new_n282), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n648), .A2(KEYINPUT99), .A3(new_n320), .A4(new_n309), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n645), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n632), .A2(new_n507), .A3(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT34), .B(G104), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G6));
  NOR2_X1   g467(.A1(new_n441), .A2(new_n443), .ZN(new_n654));
  OR2_X1    g468(.A1(new_n654), .A2(new_n509), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n450), .A2(G475), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n655), .A2(new_n656), .A3(new_n498), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n657), .B1(new_n647), .B2(new_n649), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n632), .A2(new_n507), .A3(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT35), .B(G107), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G9));
  NAND2_X1  g475(.A1(new_n616), .A2(new_n621), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n597), .A2(KEYINPUT36), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n599), .B(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n664), .A2(new_n606), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n631), .A2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n517), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT37), .B(G110), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G12));
  OR2_X1    g486(.A1(new_n503), .A2(G900), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(new_n501), .ZN(new_n674));
  AND2_X1   g488(.A1(new_n376), .A2(new_n674), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n658), .A2(new_n675), .A3(new_n570), .A4(new_n667), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G128), .ZN(G30));
  INV_X1    g491(.A(KEYINPUT38), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n317), .B(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n665), .B1(new_n616), .B2(new_n621), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n512), .A2(new_n498), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n629), .A2(KEYINPUT32), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n541), .B1(new_n555), .B2(new_n531), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n530), .A2(new_n531), .A3(new_n541), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(new_n283), .ZN(new_n688));
  OAI21_X1  g502(.A(G472), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n682), .B1(new_n685), .B2(new_n689), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n680), .A2(new_n320), .A3(new_n681), .A4(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n370), .A2(new_n375), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(KEYINPUT101), .B(KEYINPUT39), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n674), .B(new_n694), .ZN(new_n695));
  NOR3_X1   g509(.A1(new_n693), .A2(new_n325), .A3(new_n695), .ZN(new_n696));
  OR2_X1    g510(.A1(new_n696), .A2(KEYINPUT40), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(KEYINPUT40), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n691), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(new_n197), .ZN(G45));
  NAND4_X1  g514(.A1(new_n675), .A2(new_n570), .A3(new_n650), .A4(new_n667), .ZN(new_n701));
  XNOR2_X1  g515(.A(KEYINPUT102), .B(G146), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(G48));
  OAI21_X1  g517(.A(new_n283), .B1(new_n368), .B2(new_n369), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(G469), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n705), .A2(new_n324), .A3(new_n370), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n706), .A2(new_n506), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n623), .A2(new_n650), .A3(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(KEYINPUT41), .B(G113), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n708), .B(new_n709), .ZN(G15));
  NAND3_X1  g524(.A1(new_n623), .A2(new_n658), .A3(new_n707), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G116), .ZN(G18));
  AND3_X1   g526(.A1(new_n667), .A2(new_n570), .A3(new_n515), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n706), .B1(new_n647), .B2(new_n649), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G119), .ZN(G21));
  OAI21_X1  g530(.A(new_n541), .B1(new_n532), .B2(new_n535), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n561), .A2(new_n564), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(new_n567), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(KEYINPUT103), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT103), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n718), .A2(new_n721), .A3(new_n567), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n628), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  OR2_X1    g537(.A1(new_n622), .A2(KEYINPUT104), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n622), .A2(KEYINPUT104), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n723), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n647), .A2(new_n649), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n727), .A2(new_n512), .A3(new_n498), .ZN(new_n728));
  NOR3_X1   g542(.A1(new_n728), .A2(new_n506), .A3(new_n706), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n726), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G122), .ZN(G24));
  NOR2_X1   g545(.A1(new_n723), .A2(new_n681), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n512), .A2(new_n644), .A3(new_n674), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT105), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n512), .A2(new_n644), .A3(KEYINPUT105), .A4(new_n674), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n714), .A2(new_n732), .A3(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G125), .ZN(G27));
  OR2_X1    g554(.A1(new_n685), .A2(KEYINPUT108), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n685), .A2(KEYINPUT108), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n741), .A2(new_n558), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n724), .A2(new_n725), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  AND3_X1   g559(.A1(new_n306), .A2(new_n308), .A3(new_n316), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n746), .A2(new_n324), .A3(new_n692), .A4(new_n320), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n747), .A2(new_n737), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(KEYINPUT42), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n745), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n748), .A2(KEYINPUT106), .A3(new_n623), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT106), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n306), .A2(new_n320), .A3(new_n308), .A4(new_n316), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n753), .A2(new_n325), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n754), .A2(new_n692), .A3(new_n735), .A4(new_n736), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n570), .A2(new_n622), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n752), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT42), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n751), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(KEYINPUT107), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT107), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n751), .A2(new_n757), .A3(new_n761), .A4(new_n758), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n750), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(new_n353), .ZN(G33));
  AND4_X1   g578(.A1(new_n656), .A2(new_n655), .A3(new_n498), .A4(new_n674), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n570), .A2(new_n765), .A3(new_n622), .ZN(new_n766));
  OR2_X1    g580(.A1(new_n766), .A2(new_n747), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G134), .ZN(G36));
  NAND2_X1  g582(.A1(new_n451), .A2(new_n644), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT43), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n771), .A2(new_n630), .A3(new_n667), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(KEYINPUT44), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n371), .A2(new_n372), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n373), .A2(new_n365), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT45), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n374), .A2(KEYINPUT45), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n778), .A2(G469), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(G469), .A2(G902), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT46), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n780), .A2(KEYINPUT46), .A3(new_n781), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n784), .A2(new_n370), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(new_n324), .ZN(new_n787));
  NOR3_X1   g601(.A1(new_n787), .A2(new_n695), .A3(new_n753), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n773), .A2(new_n788), .ZN(new_n789));
  XOR2_X1   g603(.A(KEYINPUT109), .B(G137), .Z(new_n790));
  XNOR2_X1  g604(.A(new_n789), .B(new_n790), .ZN(G39));
  INV_X1    g605(.A(KEYINPUT47), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n787), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n786), .A2(KEYINPUT47), .A3(new_n324), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NOR4_X1   g609(.A1(new_n570), .A2(new_n622), .A3(new_n733), .A4(new_n753), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G140), .ZN(G42));
  NAND2_X1  g612(.A1(new_n705), .A2(new_n370), .ZN(new_n799));
  OR2_X1    g613(.A1(new_n799), .A2(KEYINPUT115), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(KEYINPUT115), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n800), .A2(new_n325), .A3(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n793), .A2(new_n794), .A3(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT118), .ZN(new_n804));
  OR2_X1    g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n771), .A2(new_n502), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n726), .A2(new_n806), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n807), .A2(new_n753), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n803), .A2(new_n804), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n805), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(new_n799), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n679), .A2(new_n324), .A3(new_n319), .A4(new_n811), .ZN(new_n812));
  AND2_X1   g626(.A1(KEYINPUT116), .A2(KEYINPUT50), .ZN(new_n813));
  NOR2_X1   g627(.A1(KEYINPUT116), .A2(KEYINPUT50), .ZN(new_n814));
  OAI22_X1  g628(.A1(new_n807), .A2(new_n812), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  OR2_X1    g629(.A1(new_n807), .A2(new_n812), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n815), .B1(new_n816), .B2(new_n814), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n799), .A2(new_n325), .A3(new_n753), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n806), .A2(new_n818), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n685), .A2(new_n689), .ZN(new_n820));
  AND4_X1   g634(.A1(new_n622), .A2(new_n820), .A3(new_n818), .A4(new_n502), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n512), .A2(new_n644), .ZN(new_n822));
  AOI22_X1  g636(.A1(new_n819), .A2(new_n732), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n810), .A2(KEYINPUT51), .A3(new_n817), .A4(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n726), .A2(new_n714), .A3(new_n806), .ZN(new_n825));
  XOR2_X1   g639(.A(new_n825), .B(KEYINPUT119), .Z(new_n826));
  NAND3_X1  g640(.A1(new_n819), .A2(new_n744), .A3(new_n743), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(KEYINPUT48), .ZN(new_n828));
  INV_X1    g642(.A(G952), .ZN(new_n829));
  INV_X1    g643(.A(new_n645), .ZN(new_n830));
  AOI211_X1 g644(.A(new_n829), .B(G953), .C1(new_n821), .C2(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n824), .A2(new_n826), .A3(new_n828), .A4(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n803), .A2(new_n808), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n817), .A2(new_n823), .A3(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT51), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  OR2_X1    g650(.A1(new_n836), .A2(KEYINPUT117), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(KEYINPUT117), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n832), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(new_n750), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n756), .A2(new_n747), .A3(new_n737), .ZN(new_n841));
  AOI21_X1  g655(.A(KEYINPUT42), .B1(new_n841), .B2(KEYINPUT106), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n761), .B1(new_n842), .B2(new_n757), .ZN(new_n843));
  AND4_X1   g657(.A1(new_n761), .A2(new_n751), .A3(new_n757), .A4(new_n758), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n840), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n645), .A2(KEYINPUT111), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n451), .A2(new_n498), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT111), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n512), .A2(new_n644), .A3(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n846), .A2(new_n847), .A3(new_n849), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n322), .A2(new_n850), .A3(new_n507), .ZN(new_n851));
  AOI22_X1  g665(.A1(new_n632), .A2(new_n851), .B1(new_n713), .B2(new_n714), .ZN(new_n852));
  OAI211_X1 g666(.A(new_n623), .B(new_n707), .C1(new_n650), .C2(new_n658), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n517), .B1(new_n669), .B2(new_n623), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n852), .A2(new_n730), .A3(new_n853), .A4(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n667), .A2(new_n628), .A3(new_n722), .A4(new_n720), .ZN(new_n856));
  OAI21_X1  g670(.A(KEYINPUT112), .B1(new_n856), .B2(new_n755), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT112), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n748), .A2(new_n858), .A3(new_n732), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n655), .A2(new_n656), .A3(new_n499), .A4(new_n674), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n861), .A2(new_n753), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n862), .A2(new_n570), .A3(new_n667), .A4(new_n376), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n860), .A2(new_n767), .A3(new_n863), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n855), .A2(new_n864), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n690), .A2(new_n727), .A3(new_n681), .A4(new_n675), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n739), .A2(new_n866), .A3(new_n676), .A4(new_n701), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT52), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n867), .B(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n845), .A2(new_n865), .A3(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT53), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT54), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n739), .A2(new_n676), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n874), .A2(new_n868), .A3(new_n701), .A4(new_n866), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n867), .A2(KEYINPUT52), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n739), .A2(new_n676), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(KEYINPUT52), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n875), .A2(new_n876), .A3(new_n878), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n879), .A2(KEYINPUT53), .A3(new_n845), .A4(new_n865), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n872), .A2(new_n873), .A3(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT113), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n875), .A2(new_n876), .A3(new_n878), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n632), .A2(new_n851), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n884), .A2(new_n853), .A3(new_n715), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n516), .B1(new_n756), .B2(new_n668), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n886), .B1(new_n726), .B2(new_n729), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n863), .B1(new_n747), .B2(new_n766), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n888), .B1(new_n857), .B2(new_n859), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n885), .A2(new_n887), .A3(new_n889), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n883), .A2(new_n763), .A3(new_n890), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n882), .B1(new_n891), .B2(KEYINPUT53), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n763), .A2(new_n890), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(new_n879), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n894), .A2(KEYINPUT113), .A3(new_n871), .ZN(new_n895));
  OAI21_X1  g709(.A(KEYINPUT114), .B1(new_n870), .B2(new_n871), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT114), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n893), .A2(new_n897), .A3(KEYINPUT53), .A4(new_n869), .ZN(new_n898));
  AOI22_X1  g712(.A1(new_n892), .A2(new_n895), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n839), .B(new_n881), .C1(new_n873), .C2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n829), .A2(new_n327), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n769), .A2(new_n325), .A3(new_n319), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT49), .ZN(new_n904));
  OAI211_X1 g718(.A(new_n744), .B(new_n903), .C1(new_n904), .C2(new_n811), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n905), .B(KEYINPUT110), .Z(new_n906));
  NAND2_X1  g720(.A1(new_n811), .A2(new_n904), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n906), .A2(new_n820), .A3(new_n679), .A4(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n902), .A2(new_n908), .ZN(G75));
  OR3_X1    g723(.A1(new_n327), .A2(KEYINPUT120), .A3(G952), .ZN(new_n910));
  OAI21_X1  g724(.A(KEYINPUT120), .B1(new_n327), .B2(G952), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT121), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n280), .A2(new_n281), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(new_n226), .ZN(new_n916));
  INV_X1    g730(.A(G210), .ZN(new_n917));
  AOI211_X1 g731(.A(new_n917), .B(new_n283), .C1(new_n872), .C2(new_n880), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n918), .A2(KEYINPUT55), .A3(KEYINPUT56), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT55), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n283), .B1(new_n872), .B2(new_n880), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n921), .A2(G210), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT56), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n920), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n916), .B1(new_n919), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(KEYINPUT55), .B1(new_n918), .B2(KEYINPUT56), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n922), .A2(new_n920), .A3(new_n923), .ZN(new_n927));
  INV_X1    g741(.A(new_n916), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n914), .B1(new_n925), .B2(new_n929), .ZN(G51));
  AOI211_X1 g744(.A(new_n283), .B(new_n780), .C1(new_n872), .C2(new_n880), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n781), .B(KEYINPUT57), .Z(new_n932));
  AND3_X1   g746(.A1(new_n872), .A2(new_n873), .A3(new_n880), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n873), .B1(new_n872), .B2(new_n880), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n932), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n368), .A2(new_n369), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n931), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(KEYINPUT122), .B1(new_n938), .B2(new_n912), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT122), .ZN(new_n940));
  INV_X1    g754(.A(new_n912), .ZN(new_n941));
  AOI21_X1  g755(.A(KEYINPUT53), .B1(new_n893), .B2(new_n869), .ZN(new_n942));
  NOR4_X1   g756(.A1(new_n883), .A2(new_n763), .A3(new_n890), .A4(new_n871), .ZN(new_n943));
  OAI21_X1  g757(.A(KEYINPUT54), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(new_n881), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n936), .B1(new_n945), .B2(new_n932), .ZN(new_n946));
  OAI211_X1 g760(.A(new_n940), .B(new_n941), .C1(new_n946), .C2(new_n931), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n939), .A2(new_n947), .ZN(G54));
  NAND3_X1  g762(.A1(new_n921), .A2(KEYINPUT58), .A3(G475), .ZN(new_n949));
  OR2_X1    g763(.A1(new_n949), .A2(new_n437), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n437), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n912), .B1(new_n950), .B2(new_n951), .ZN(G60));
  OR2_X1    g766(.A1(new_n637), .A2(new_n638), .ZN(new_n953));
  NAND2_X1  g767(.A1(G478), .A2(G902), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT59), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(KEYINPUT123), .B1(new_n945), .B2(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT123), .ZN(new_n959));
  AOI211_X1 g773(.A(new_n959), .B(new_n956), .C1(new_n944), .C2(new_n881), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n913), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n881), .B1(new_n899), .B2(new_n873), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n953), .B1(new_n962), .B2(new_n955), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n961), .A2(new_n963), .ZN(G63));
  NAND2_X1  g778(.A1(G217), .A2(G902), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(KEYINPUT60), .Z(new_n966));
  OAI21_X1  g780(.A(new_n966), .B1(new_n942), .B2(new_n943), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n914), .B1(new_n967), .B2(new_n603), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n968), .B1(new_n664), .B2(new_n967), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT61), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n969), .B(new_n970), .ZN(G66));
  OAI21_X1  g785(.A(G953), .B1(new_n505), .B2(new_n187), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n855), .B(KEYINPUT124), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n972), .B1(new_n973), .B2(G953), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n915), .B1(G898), .B2(new_n327), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n974), .B(new_n975), .ZN(G69));
  AOI22_X1  g790(.A1(new_n788), .A2(new_n773), .B1(new_n795), .B2(new_n796), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n850), .B(KEYINPUT125), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n756), .A2(new_n753), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n978), .A2(new_n696), .A3(new_n979), .ZN(new_n980));
  AND2_X1   g794(.A1(new_n977), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n739), .A2(new_n676), .A3(new_n701), .ZN(new_n982));
  OAI21_X1  g796(.A(KEYINPUT62), .B1(new_n699), .B2(new_n982), .ZN(new_n983));
  OR3_X1    g797(.A1(new_n699), .A2(KEYINPUT62), .A3(new_n982), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n981), .A2(KEYINPUT126), .A3(new_n983), .A4(new_n984), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n984), .A2(new_n977), .A3(new_n983), .A4(new_n980), .ZN(new_n986));
  INV_X1    g800(.A(KEYINPUT126), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n985), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n989), .A2(new_n327), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT127), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n553), .A2(new_n554), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n404), .A2(new_n406), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n992), .B(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(new_n994), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n990), .A2(new_n991), .A3(new_n995), .ZN(new_n996));
  OR4_X1    g810(.A1(new_n695), .A2(new_n745), .A3(new_n728), .A4(new_n787), .ZN(new_n997));
  INV_X1    g811(.A(new_n982), .ZN(new_n998));
  NAND4_X1  g812(.A1(new_n977), .A2(new_n997), .A3(new_n767), .A4(new_n998), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n999), .A2(new_n763), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n1000), .A2(new_n327), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n995), .B1(G900), .B2(G953), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g817(.A(G953), .B1(new_n985), .B2(new_n988), .ZN(new_n1004));
  OAI21_X1  g818(.A(KEYINPUT127), .B1(new_n1004), .B2(new_n994), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n996), .A2(new_n1003), .A3(new_n1005), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n327), .B1(G227), .B2(G900), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g822(.A(new_n1007), .ZN(new_n1009));
  NAND4_X1  g823(.A1(new_n996), .A2(new_n1005), .A3(new_n1009), .A4(new_n1003), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1008), .A2(new_n1010), .ZN(G72));
  NAND2_X1  g825(.A1(G472), .A2(G902), .ZN(new_n1012));
  XOR2_X1   g826(.A(new_n1012), .B(KEYINPUT63), .Z(new_n1013));
  NAND2_X1  g827(.A1(new_n556), .A2(new_n1013), .ZN(new_n1014));
  NOR3_X1   g828(.A1(new_n899), .A2(new_n686), .A3(new_n1014), .ZN(new_n1015));
  INV_X1    g829(.A(new_n686), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n985), .A2(new_n988), .A3(new_n973), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1016), .B1(new_n1017), .B2(new_n1013), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1000), .A2(new_n973), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n556), .B1(new_n1019), .B2(new_n1013), .ZN(new_n1020));
  NOR4_X1   g834(.A1(new_n1015), .A2(new_n912), .A3(new_n1018), .A4(new_n1020), .ZN(G57));
endmodule


