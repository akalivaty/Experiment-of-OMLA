//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 0 0 1 1 0 1 1 1 0 0 1 1 0 1 1 1 0 0 0 0 1 1 0 1 1 1 0 1 0 1 1 1 1 1 1 1 0 0 1 1 1 1 1 1 0 1 1 1 1 0 0 0 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:19 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n570, new_n572, new_n573,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n586, new_n587, new_n588, new_n590,
    new_n591, new_n592, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n630,
    new_n633, new_n634, new_n636, new_n637, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1191, new_n1192, new_n1193, new_n1195, new_n1196, new_n1197;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT64), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(G567), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  INV_X1    g031(.A(new_n451), .ZN(new_n457));
  AOI21_X1  g032(.A(new_n456), .B1(new_n457), .B2(G2106), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  NAND3_X1  g034(.A1(new_n459), .A2(G101), .A3(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(KEYINPUT65), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT65), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2105), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  OAI211_X1 g040(.A(new_n461), .B(new_n463), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G137), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n460), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT68), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  OAI211_X1 g045(.A(KEYINPUT68), .B(new_n460), .C1(new_n466), .C2(new_n467), .ZN(new_n471));
  AND2_X1   g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n461), .A2(new_n463), .ZN(new_n473));
  INV_X1    g048(.A(G125), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT3), .ZN(new_n475));
  INV_X1    g050(.A(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n474), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(G113), .A2(G2104), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(KEYINPUT66), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT66), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n482), .A2(G113), .A3(G2104), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n473), .B1(new_n479), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(KEYINPUT67), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT67), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(new_n473), .C1(new_n479), .C2(new_n484), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n472), .A2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G160));
  NOR2_X1   g066(.A1(new_n464), .A2(new_n465), .ZN(new_n492));
  XNOR2_X1  g067(.A(KEYINPUT65), .B(G2105), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G124), .ZN(new_n495));
  OAI221_X1 g070(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n493), .C2(G112), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n492), .A2(G2105), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(G136), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT69), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n498), .A2(KEYINPUT69), .A3(G136), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n497), .B1(new_n501), .B2(new_n502), .ZN(G162));
  INV_X1    g078(.A(G138), .ZN(new_n504));
  OAI21_X1  g079(.A(KEYINPUT4), .B1(new_n466), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n477), .A2(new_n478), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT4), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n506), .A2(new_n493), .A3(new_n507), .A4(G138), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g084(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n510));
  INV_X1    g085(.A(G114), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n510), .B1(new_n511), .B2(G2105), .ZN(new_n512));
  AND2_X1   g087(.A1(G126), .A2(G2105), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n513), .B1(new_n464), .B2(new_n465), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT70), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n506), .A2(KEYINPUT70), .A3(new_n513), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n512), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n509), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(new_n519), .ZN(G164));
  INV_X1    g095(.A(KEYINPUT5), .ZN(new_n521));
  INV_X1    g096(.A(G543), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(KEYINPUT5), .A2(G543), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(KEYINPUT6), .A2(G651), .ZN(new_n526));
  AND2_X1   g101(.A1(KEYINPUT6), .A2(G651), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(new_n528), .ZN(new_n529));
  OAI21_X1  g104(.A(G543), .B1(new_n527), .B2(new_n526), .ZN(new_n530));
  INV_X1    g105(.A(new_n530), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n529), .A2(G88), .B1(G50), .B2(new_n531), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n525), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n533));
  INV_X1    g108(.A(G651), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT71), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NOR3_X1   g112(.A1(new_n533), .A2(KEYINPUT71), .A3(new_n534), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n532), .B1(new_n537), .B2(new_n538), .ZN(G303));
  INV_X1    g114(.A(G303), .ZN(G166));
  NOR2_X1   g115(.A1(new_n527), .A2(new_n526), .ZN(new_n541));
  INV_X1    g116(.A(G89), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(G63), .A2(G651), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n525), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n531), .A2(G51), .ZN(new_n547));
  NAND3_X1  g122(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT7), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n546), .A2(new_n547), .A3(new_n549), .ZN(G286));
  INV_X1    g125(.A(G286), .ZN(G168));
  INV_X1    g126(.A(G90), .ZN(new_n552));
  INV_X1    g127(.A(G52), .ZN(new_n553));
  OAI22_X1  g128(.A1(new_n528), .A2(new_n552), .B1(new_n553), .B2(new_n530), .ZN(new_n554));
  AND2_X1   g129(.A1(new_n523), .A2(new_n524), .ZN(new_n555));
  INV_X1    g130(.A(G64), .ZN(new_n556));
  INV_X1    g131(.A(G77), .ZN(new_n557));
  OAI22_X1  g132(.A1(new_n555), .A2(new_n556), .B1(new_n557), .B2(new_n522), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT72), .ZN(new_n559));
  AOI21_X1  g134(.A(new_n534), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  OAI221_X1 g135(.A(KEYINPUT72), .B1(new_n557), .B2(new_n522), .C1(new_n555), .C2(new_n556), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n554), .B1(new_n560), .B2(new_n561), .ZN(G171));
  NAND2_X1  g137(.A1(new_n531), .A2(G43), .ZN(new_n563));
  INV_X1    g138(.A(G81), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n564), .B2(new_n528), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n525), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n566), .A2(new_n534), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G860), .ZN(G153));
  AND3_X1   g144(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G36), .ZN(G176));
  NAND2_X1  g146(.A1(G1), .A2(G3), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT8), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n570), .A2(new_n573), .ZN(G188));
  OAI211_X1 g149(.A(G53), .B(G543), .C1(new_n527), .C2(new_n526), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n575), .B(KEYINPUT9), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n525), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n578));
  INV_X1    g153(.A(G91), .ZN(new_n579));
  OAI22_X1  g154(.A1(new_n578), .A2(new_n534), .B1(new_n528), .B2(new_n579), .ZN(new_n580));
  NOR3_X1   g155(.A1(new_n577), .A2(new_n580), .A3(KEYINPUT73), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT73), .ZN(new_n582));
  INV_X1    g157(.A(new_n580), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n582), .B1(new_n583), .B2(new_n576), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n581), .A2(new_n584), .ZN(G299));
  NAND2_X1  g160(.A1(new_n558), .A2(new_n559), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n586), .A2(G651), .A3(new_n561), .ZN(new_n587));
  INV_X1    g162(.A(new_n554), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(G301));
  NAND2_X1  g164(.A1(new_n529), .A2(G87), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n531), .A2(G49), .ZN(new_n591));
  OAI21_X1  g166(.A(G651), .B1(new_n525), .B2(G74), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(G288));
  INV_X1    g168(.A(G61), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n594), .B1(new_n523), .B2(new_n524), .ZN(new_n595));
  AND2_X1   g170(.A1(G73), .A2(G543), .ZN(new_n596));
  OAI21_X1  g171(.A(G651), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n597), .A2(KEYINPUT74), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT74), .ZN(new_n599));
  OAI211_X1 g174(.A(new_n599), .B(G651), .C1(new_n595), .C2(new_n596), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(G86), .ZN(new_n602));
  INV_X1    g177(.A(G48), .ZN(new_n603));
  OAI22_X1  g178(.A1(new_n528), .A2(new_n602), .B1(new_n603), .B2(new_n530), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n601), .A2(new_n605), .ZN(G305));
  AOI22_X1  g181(.A1(new_n525), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n607), .A2(new_n534), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT75), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n608), .B(new_n609), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n529), .A2(G85), .B1(G47), .B2(new_n531), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(G290));
  INV_X1    g187(.A(G868), .ZN(new_n613));
  NOR2_X1   g188(.A1(G171), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(G79), .A2(G543), .ZN(new_n615));
  INV_X1    g190(.A(G66), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n555), .B2(new_n616), .ZN(new_n617));
  OR2_X1    g192(.A1(new_n530), .A2(KEYINPUT76), .ZN(new_n618));
  INV_X1    g193(.A(G54), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n619), .B1(new_n530), .B2(KEYINPUT76), .ZN(new_n620));
  AOI22_X1  g195(.A1(G651), .A2(new_n617), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n529), .A2(G92), .ZN(new_n622));
  INV_X1    g197(.A(KEYINPUT10), .ZN(new_n623));
  NOR2_X1   g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AOI21_X1  g199(.A(KEYINPUT10), .B1(new_n529), .B2(G92), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n621), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n614), .B1(new_n613), .B2(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT77), .ZN(G284));
  XNOR2_X1  g203(.A(new_n627), .B(KEYINPUT78), .ZN(G321));
  NAND2_X1  g204(.A1(G299), .A2(new_n613), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n630), .B1(new_n613), .B2(G168), .ZN(G297));
  OAI21_X1  g206(.A(new_n630), .B1(new_n613), .B2(G168), .ZN(G280));
  INV_X1    g207(.A(new_n626), .ZN(new_n633));
  INV_X1    g208(.A(G559), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n633), .B1(new_n634), .B2(G860), .ZN(G148));
  NAND2_X1  g210(.A1(new_n633), .A2(new_n634), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(G868), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n637), .B1(G868), .B2(new_n568), .ZN(G323));
  XNOR2_X1  g213(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g214(.A1(new_n498), .A2(G2104), .ZN(new_n640));
  XOR2_X1   g215(.A(KEYINPUT79), .B(KEYINPUT12), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(KEYINPUT13), .B(G2100), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n494), .A2(G123), .ZN(new_n645));
  OAI221_X1 g220(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n493), .C2(G111), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n498), .A2(G135), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n645), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n648), .A2(KEYINPUT80), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n648), .A2(KEYINPUT80), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  AND2_X1   g227(.A1(new_n652), .A2(G2096), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n652), .A2(G2096), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n644), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n655), .B(KEYINPUT81), .Z(G156));
  XOR2_X1   g231(.A(KEYINPUT82), .B(KEYINPUT14), .Z(new_n657));
  XNOR2_X1  g232(.A(KEYINPUT15), .B(G2435), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(G2438), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2427), .B(G2430), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n657), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n661), .B1(new_n659), .B2(new_n660), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2451), .B(G2454), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT16), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1341), .B(G1348), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n662), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G2443), .B(G2446), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n669), .A2(G14), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n667), .A2(new_n668), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n670), .A2(new_n671), .ZN(G401));
  XNOR2_X1  g247(.A(G2067), .B(G2678), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT83), .ZN(new_n674));
  XOR2_X1   g249(.A(G2084), .B(G2090), .Z(new_n675));
  NAND2_X1  g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G2072), .B(G2078), .Z(new_n677));
  NOR2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT18), .ZN(new_n679));
  OR2_X1    g254(.A1(new_n674), .A2(new_n675), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n677), .B(KEYINPUT17), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n680), .A2(new_n676), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n677), .B(KEYINPUT84), .ZN(new_n683));
  OAI211_X1 g258(.A(new_n679), .B(new_n682), .C1(new_n680), .C2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(G2100), .ZN(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT85), .B(G2096), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(G227));
  XNOR2_X1  g262(.A(G1971), .B(G1976), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT86), .B(KEYINPUT19), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1956), .B(G2474), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1961), .B(G1966), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT20), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n690), .A2(KEYINPUT87), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n691), .A2(new_n692), .ZN(new_n697));
  INV_X1    g272(.A(new_n693), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n697), .B1(new_n690), .B2(new_n698), .ZN(new_n699));
  OR2_X1    g274(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n696), .A2(new_n699), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n695), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(G1991), .B(G1996), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(G1981), .B(G1986), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(G229));
  NOR2_X1   g283(.A1(G16), .A2(G22), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(G166), .B2(G16), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(G1971), .Z(new_n711));
  NOR2_X1   g286(.A1(G16), .A2(G23), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(KEYINPUT90), .Z(new_n713));
  INV_X1    g288(.A(G16), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n713), .B1(G288), .B2(new_n714), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT33), .B(G1976), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(G305), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n718), .A2(new_n714), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(G6), .B2(new_n714), .ZN(new_n720));
  XOR2_X1   g295(.A(KEYINPUT32), .B(G1981), .Z(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT89), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n717), .B1(new_n720), .B2(new_n722), .ZN(new_n723));
  OR2_X1    g298(.A1(new_n720), .A2(new_n722), .ZN(new_n724));
  AND3_X1   g299(.A1(new_n711), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(KEYINPUT34), .ZN(new_n726));
  OR2_X1    g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n725), .A2(new_n726), .ZN(new_n728));
  MUX2_X1   g303(.A(G24), .B(G290), .S(G16), .Z(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(G1986), .Z(new_n730));
  INV_X1    g305(.A(G29), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(G25), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n494), .A2(G119), .ZN(new_n733));
  OAI221_X1 g308(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n493), .C2(G107), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n498), .A2(G131), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n733), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n732), .B1(new_n737), .B2(new_n731), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT88), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT35), .B(G1991), .Z(new_n740));
  XOR2_X1   g315(.A(new_n739), .B(new_n740), .Z(new_n741));
  NAND4_X1  g316(.A1(new_n727), .A2(new_n728), .A3(new_n730), .A4(new_n741), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT36), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n652), .A2(G29), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT99), .ZN(new_n745));
  NOR2_X1   g320(.A1(G16), .A2(G19), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(new_n568), .B2(G16), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT93), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n745), .B1(G1341), .B2(new_n748), .ZN(new_n749));
  NOR2_X1   g324(.A1(G171), .A2(new_n714), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(G5), .B2(new_n714), .ZN(new_n751));
  INV_X1    g326(.A(G1961), .ZN(new_n752));
  INV_X1    g327(.A(G2084), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n731), .B1(KEYINPUT24), .B2(G34), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(KEYINPUT24), .B2(G34), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(new_n490), .B2(G29), .ZN(new_n756));
  OAI22_X1  g331(.A1(new_n751), .A2(new_n752), .B1(new_n753), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n748), .A2(G1341), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n714), .A2(G21), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G168), .B2(new_n714), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n731), .A2(G26), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT28), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n494), .A2(G128), .ZN(new_n763));
  OAI221_X1 g338(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n493), .C2(G116), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n498), .A2(G140), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n763), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(new_n766), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n762), .B1(new_n767), .B2(new_n731), .ZN(new_n768));
  XNOR2_X1  g343(.A(KEYINPUT94), .B(G2067), .ZN(new_n769));
  OAI22_X1  g344(.A1(new_n760), .A2(G1966), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(new_n768), .B2(new_n769), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n751), .A2(new_n752), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n731), .A2(G27), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G164), .B2(new_n731), .ZN(new_n774));
  INV_X1    g349(.A(G2078), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NAND4_X1  g351(.A1(new_n758), .A2(new_n771), .A3(new_n772), .A4(new_n776), .ZN(new_n777));
  NOR3_X1   g352(.A1(new_n749), .A2(new_n757), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(G299), .A2(G16), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n714), .A2(G20), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT23), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(G1956), .ZN(new_n783));
  NOR2_X1   g358(.A1(G4), .A2(G16), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT91), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(new_n626), .B2(new_n714), .ZN(new_n786));
  XOR2_X1   g361(.A(KEYINPUT92), .B(G1348), .Z(new_n787));
  NOR2_X1   g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  AND2_X1   g363(.A1(new_n786), .A2(new_n787), .ZN(new_n789));
  AND2_X1   g364(.A1(new_n756), .A2(new_n753), .ZN(new_n790));
  NOR4_X1   g365(.A1(new_n783), .A2(new_n788), .A3(new_n789), .A4(new_n790), .ZN(new_n791));
  NOR2_X1   g366(.A1(G29), .A2(G33), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT95), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n493), .A2(G103), .A3(G2104), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT25), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(G139), .B2(new_n498), .ZN(new_n796));
  AOI22_X1  g371(.A1(new_n506), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n797), .A2(new_n493), .ZN(new_n798));
  INV_X1    g373(.A(KEYINPUT96), .ZN(new_n799));
  OR2_X1    g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n798), .A2(new_n799), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n796), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(KEYINPUT97), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND4_X1  g379(.A1(new_n796), .A2(KEYINPUT97), .A3(new_n800), .A4(new_n801), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n793), .B1(new_n806), .B2(new_n731), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(G2072), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n731), .A2(G35), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(G162), .B2(new_n731), .ZN(new_n810));
  XOR2_X1   g385(.A(new_n810), .B(KEYINPUT29), .Z(new_n811));
  INV_X1    g386(.A(G2090), .ZN(new_n812));
  AND2_X1   g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n731), .A2(G32), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n494), .A2(G129), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT98), .ZN(new_n816));
  AND3_X1   g391(.A1(new_n459), .A2(G105), .A3(G2104), .ZN(new_n817));
  NAND3_X1  g392(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT26), .ZN(new_n819));
  AOI211_X1 g394(.A(new_n817), .B(new_n819), .C1(G141), .C2(new_n498), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n816), .A2(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(new_n821), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n814), .B1(new_n822), .B2(new_n731), .ZN(new_n823));
  XOR2_X1   g398(.A(KEYINPUT27), .B(G1996), .Z(new_n824));
  OR2_X1    g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n823), .A2(new_n824), .ZN(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT31), .B(G11), .ZN(new_n827));
  XOR2_X1   g402(.A(KEYINPUT30), .B(G28), .Z(new_n828));
  OAI21_X1  g403(.A(new_n827), .B1(new_n828), .B2(G29), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n829), .B1(new_n760), .B2(G1966), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n825), .A2(new_n826), .A3(new_n830), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n811), .A2(new_n812), .ZN(new_n832));
  NOR3_X1   g407(.A1(new_n813), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  AND4_X1   g408(.A1(new_n778), .A2(new_n791), .A3(new_n808), .A4(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n743), .A2(new_n834), .ZN(G150));
  INV_X1    g410(.A(G150), .ZN(G311));
  AOI22_X1  g411(.A1(new_n525), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n837));
  OR2_X1    g412(.A1(new_n837), .A2(new_n534), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n529), .A2(G93), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT100), .ZN(new_n840));
  OAI211_X1 g415(.A(G55), .B(G543), .C1(new_n527), .C2(new_n526), .ZN(new_n841));
  NAND4_X1  g416(.A1(new_n838), .A2(new_n839), .A3(new_n840), .A4(new_n841), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n837), .A2(new_n534), .ZN(new_n843));
  INV_X1    g418(.A(G93), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n841), .B1(new_n528), .B2(new_n844), .ZN(new_n845));
  OAI21_X1  g420(.A(KEYINPUT100), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n842), .A2(new_n568), .A3(new_n846), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n838), .A2(new_n841), .A3(new_n839), .ZN(new_n848));
  OAI221_X1 g423(.A(new_n563), .B1(new_n528), .B2(new_n564), .C1(new_n534), .C2(new_n566), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n848), .A2(new_n849), .A3(KEYINPUT100), .ZN(new_n850));
  AND2_X1   g425(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT38), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n626), .A2(new_n634), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT39), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n856), .B(KEYINPUT101), .Z(new_n857));
  AOI21_X1  g432(.A(G860), .B1(new_n854), .B2(new_n855), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n848), .A2(G860), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n860), .B(KEYINPUT37), .Z(new_n861));
  NAND2_X1  g436(.A1(new_n859), .A2(new_n861), .ZN(G145));
  INV_X1    g437(.A(KEYINPUT103), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n806), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n804), .A2(KEYINPUT103), .A3(new_n805), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n822), .A2(new_n767), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n821), .A2(new_n766), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n866), .A2(new_n519), .A3(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n519), .B1(new_n866), .B2(new_n867), .ZN(new_n870));
  OAI211_X1 g445(.A(new_n864), .B(new_n865), .C1(new_n869), .C2(new_n870), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n806), .A2(new_n863), .ZN(new_n872));
  INV_X1    g447(.A(new_n870), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n872), .A2(new_n873), .A3(new_n868), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(KEYINPUT104), .B(KEYINPUT105), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n494), .A2(G130), .ZN(new_n878));
  OAI221_X1 g453(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n493), .C2(G118), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n498), .A2(G142), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  OR2_X1    g456(.A1(new_n642), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n881), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n882), .A2(new_n736), .A3(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n736), .B1(new_n882), .B2(new_n883), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n877), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n886), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n888), .A2(new_n876), .A3(new_n884), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n875), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT106), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n871), .A2(new_n874), .A3(new_n890), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  AND3_X1   g470(.A1(new_n649), .A2(KEYINPUT102), .A3(new_n650), .ZN(new_n896));
  AOI21_X1  g471(.A(KEYINPUT102), .B1(new_n649), .B2(new_n650), .ZN(new_n897));
  OR3_X1    g472(.A1(new_n896), .A2(new_n897), .A3(G160), .ZN(new_n898));
  OAI21_X1  g473(.A(G160), .B1(new_n896), .B2(new_n897), .ZN(new_n899));
  AND3_X1   g474(.A1(new_n898), .A2(G162), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(G162), .B1(new_n898), .B2(new_n899), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n890), .B1(new_n871), .B2(new_n874), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n902), .B1(new_n903), .B2(KEYINPUT106), .ZN(new_n904));
  AOI21_X1  g479(.A(G37), .B1(new_n895), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT107), .ZN(new_n906));
  INV_X1    g481(.A(new_n894), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n907), .A2(new_n903), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n906), .B1(new_n908), .B2(new_n902), .ZN(new_n909));
  AND4_X1   g484(.A1(new_n906), .A2(new_n892), .A3(new_n894), .A4(new_n902), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n905), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(KEYINPUT108), .B(KEYINPUT40), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n911), .B(new_n912), .ZN(G395));
  NAND2_X1  g488(.A1(new_n848), .A2(new_n613), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n851), .B(new_n636), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n626), .B1(new_n581), .B2(new_n584), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n622), .B(new_n623), .ZN(new_n917));
  OAI21_X1  g492(.A(KEYINPUT73), .B1(new_n577), .B2(new_n580), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n583), .A2(new_n582), .A3(new_n576), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n917), .A2(new_n918), .A3(new_n919), .A4(new_n621), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n916), .A2(new_n920), .A3(KEYINPUT109), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT109), .ZN(new_n922));
  NAND3_X1  g497(.A1(G299), .A2(new_n922), .A3(new_n633), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  OR2_X1    g499(.A1(new_n915), .A2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT110), .ZN(new_n926));
  OR2_X1    g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n921), .A2(KEYINPUT41), .A3(new_n923), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT41), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n916), .A2(new_n920), .A3(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n915), .A2(new_n928), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n925), .A2(new_n926), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n927), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(G288), .ZN(new_n934));
  XNOR2_X1  g509(.A(G290), .B(new_n934), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n718), .B(G303), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n935), .B(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n937), .B(KEYINPUT42), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n933), .B(new_n938), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n914), .B1(new_n939), .B2(new_n613), .ZN(G295));
  OAI21_X1  g515(.A(new_n914), .B1(new_n939), .B2(new_n613), .ZN(G331));
  INV_X1    g516(.A(KEYINPUT44), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT115), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT112), .ZN(new_n944));
  NAND3_X1  g519(.A1(G301), .A2(new_n944), .A3(G168), .ZN(new_n945));
  OAI21_X1  g520(.A(KEYINPUT112), .B1(G171), .B2(G286), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n587), .A2(G286), .A3(new_n588), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT113), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(G171), .A2(KEYINPUT113), .A3(G286), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n947), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n851), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n947), .A2(new_n952), .A3(new_n851), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n916), .A2(new_n920), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(KEYINPUT41), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n955), .A2(new_n956), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(KEYINPUT41), .B1(new_n921), .B2(new_n923), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n943), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  AND3_X1   g536(.A1(new_n947), .A2(new_n952), .A3(new_n851), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n851), .B1(new_n947), .B2(new_n952), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n924), .A2(new_n929), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n964), .A2(KEYINPUT115), .A3(new_n965), .A4(new_n958), .ZN(new_n966));
  OAI211_X1 g541(.A(new_n923), .B(new_n921), .C1(new_n962), .C2(new_n963), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n961), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(new_n937), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n928), .A2(new_n955), .A3(new_n930), .A4(new_n956), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n937), .A2(new_n971), .A3(new_n967), .ZN(new_n972));
  INV_X1    g547(.A(G37), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n970), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(KEYINPUT43), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n937), .B1(new_n967), .B2(new_n971), .ZN(new_n978));
  XOR2_X1   g553(.A(KEYINPUT111), .B(KEYINPUT43), .Z(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  OR3_X1    g555(.A1(new_n974), .A2(new_n978), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n942), .B1(new_n977), .B2(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n970), .A2(new_n975), .A3(new_n979), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(KEYINPUT116), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT116), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n970), .A2(new_n985), .A3(new_n975), .A4(new_n979), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n980), .B1(new_n974), .B2(new_n978), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(KEYINPUT114), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT114), .ZN(new_n989));
  OAI211_X1 g564(.A(new_n989), .B(new_n980), .C1(new_n974), .C2(new_n978), .ZN(new_n990));
  AOI22_X1  g565(.A1(new_n984), .A2(new_n986), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n982), .B1(new_n991), .B2(new_n942), .ZN(G397));
  NAND4_X1  g567(.A1(new_n489), .A2(G40), .A3(new_n470), .A4(new_n471), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT117), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n472), .A2(KEYINPUT117), .A3(G40), .A4(new_n489), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(G1384), .B1(new_n509), .B2(new_n518), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n998), .A2(KEYINPUT45), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(G2067), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n767), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n766), .A2(G2067), .ZN(new_n1004));
  AND2_X1   g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n822), .A2(G1996), .ZN(new_n1006));
  INV_X1    g581(.A(G1996), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n821), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1005), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n737), .A2(new_n740), .ZN(new_n1011));
  OR2_X1    g586(.A1(new_n737), .A2(new_n740), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1010), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g588(.A(G290), .B(G1986), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1001), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT118), .ZN(new_n1016));
  AND3_X1   g591(.A1(new_n998), .A2(new_n1016), .A3(KEYINPUT45), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1016), .B1(new_n998), .B2(KEYINPUT45), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(new_n999), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n1019), .A2(new_n997), .A3(new_n775), .A4(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT53), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g598(.A(new_n998), .B(KEYINPUT50), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n997), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(new_n752), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n999), .B1(new_n995), .B2(new_n996), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT45), .ZN(new_n1028));
  AOI211_X1 g603(.A(new_n1028), .B(G1384), .C1(new_n509), .C2(new_n518), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1027), .A2(KEYINPUT53), .A3(new_n775), .A4(new_n1030), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1023), .A2(G301), .A3(new_n1026), .A4(new_n1031), .ZN(new_n1032));
  AND2_X1   g607(.A1(new_n1032), .A2(KEYINPUT54), .ZN(new_n1033));
  AOI22_X1  g608(.A1(new_n1021), .A2(new_n1022), .B1(new_n752), .B2(new_n1025), .ZN(new_n1034));
  XOR2_X1   g609(.A(KEYINPUT125), .B(G2078), .Z(new_n1035));
  AND4_X1   g610(.A1(KEYINPUT53), .A2(new_n485), .A3(G40), .A4(new_n1035), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n1019), .A2(new_n472), .A3(new_n1020), .A4(new_n1036), .ZN(new_n1037));
  AOI211_X1 g612(.A(KEYINPUT126), .B(G301), .C1(new_n1034), .C2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT126), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1023), .A2(new_n1026), .A3(new_n1037), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1039), .B1(new_n1040), .B2(G171), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1033), .B1(new_n1038), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT54), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1040), .A2(G171), .ZN(new_n1044));
  AOI21_X1  g619(.A(G301), .B1(new_n1034), .B2(new_n1031), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1043), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n997), .A2(new_n753), .A3(new_n1024), .ZN(new_n1047));
  AOI211_X1 g622(.A(new_n1029), .B(new_n999), .C1(new_n995), .C2(new_n996), .ZN(new_n1048));
  OAI211_X1 g623(.A(G168), .B(new_n1047), .C1(new_n1048), .C2(G1966), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(G8), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n997), .A2(new_n1020), .A3(new_n1030), .ZN(new_n1051));
  INV_X1    g626(.A(G1966), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(G168), .B1(new_n1053), .B2(new_n1047), .ZN(new_n1054));
  OAI21_X1  g629(.A(KEYINPUT51), .B1(new_n1050), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT51), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1049), .A2(new_n1056), .A3(G8), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT52), .ZN(new_n1059));
  INV_X1    g634(.A(G1384), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n519), .A2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1061), .B1(new_n995), .B2(new_n996), .ZN(new_n1062));
  INV_X1    g637(.A(G8), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(G1976), .ZN(new_n1065));
  NOR2_X1   g640(.A1(G288), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1059), .B1(new_n1064), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT49), .ZN(new_n1069));
  INV_X1    g644(.A(G1981), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n601), .A2(new_n1070), .A3(new_n605), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1070), .B1(new_n601), .B2(new_n605), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1069), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1073), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1075), .A2(KEYINPUT49), .A3(new_n1071), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1077));
  NOR3_X1   g652(.A1(new_n1077), .A2(new_n1063), .A3(new_n1062), .ZN(new_n1078));
  XNOR2_X1  g653(.A(KEYINPUT119), .B(G1976), .ZN(new_n1079));
  NAND2_X1  g654(.A1(G288), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(new_n1059), .ZN(new_n1081));
  NOR4_X1   g656(.A1(new_n1062), .A2(new_n1063), .A3(new_n1066), .A4(new_n1081), .ZN(new_n1082));
  NOR3_X1   g657(.A1(new_n1068), .A2(new_n1078), .A3(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(G1971), .B1(new_n1027), .B2(new_n1019), .ZN(new_n1084));
  AND3_X1   g659(.A1(new_n997), .A2(new_n812), .A3(new_n1024), .ZN(new_n1085));
  OAI21_X1  g660(.A(G8), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(G303), .A2(G8), .ZN(new_n1087));
  XNOR2_X1  g662(.A(new_n1087), .B(KEYINPUT55), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1088), .ZN(new_n1090));
  OAI211_X1 g665(.A(new_n1090), .B(G8), .C1(new_n1084), .C2(new_n1085), .ZN(new_n1091));
  AND3_X1   g666(.A1(new_n1083), .A2(new_n1089), .A3(new_n1091), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1042), .A2(new_n1046), .A3(new_n1058), .A4(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n997), .A2(new_n998), .ZN(new_n1094));
  XOR2_X1   g669(.A(KEYINPUT58), .B(G1341), .Z(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1027), .A2(new_n1007), .A3(new_n1019), .ZN(new_n1097));
  AND2_X1   g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g673(.A(KEYINPUT124), .B1(new_n1098), .B2(new_n849), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT59), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n849), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT124), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1099), .A2(new_n1100), .A3(new_n1103), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1105));
  AOI211_X1 g680(.A(KEYINPUT124), .B(new_n849), .C1(new_n1096), .C2(new_n1097), .ZN(new_n1106));
  OAI21_X1  g681(.A(KEYINPUT59), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1104), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT60), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT123), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n997), .A2(new_n1110), .A3(new_n1002), .A4(new_n998), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1061), .A2(KEYINPUT50), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT50), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n998), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1115), .B1(new_n996), .B2(new_n995), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1111), .B1(new_n1116), .B2(G1348), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1110), .B1(new_n1062), .B2(new_n1002), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1109), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(KEYINPUT123), .B1(new_n1094), .B2(G2067), .ZN(new_n1120));
  INV_X1    g695(.A(G1348), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1025), .A2(new_n1121), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1120), .A2(KEYINPUT60), .A3(new_n1111), .A4(new_n1122), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1119), .A2(new_n633), .A3(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1117), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1125), .A2(KEYINPUT60), .A3(new_n626), .A4(new_n1120), .ZN(new_n1126));
  AND2_X1   g701(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  XNOR2_X1  g702(.A(KEYINPUT56), .B(G2072), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1027), .A2(new_n1019), .A3(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(KEYINPUT122), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT122), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1027), .A2(new_n1131), .A3(new_n1019), .A4(new_n1128), .ZN(new_n1132));
  INV_X1    g707(.A(G1956), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1025), .A2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1130), .A2(new_n1132), .A3(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n583), .A2(new_n576), .ZN(new_n1136));
  AOI21_X1  g711(.A(KEYINPUT57), .B1(new_n576), .B2(KEYINPUT121), .ZN(new_n1137));
  XOR2_X1   g712(.A(new_n1136), .B(new_n1137), .Z(new_n1138));
  NAND2_X1  g713(.A1(new_n1135), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1138), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1130), .A2(new_n1140), .A3(new_n1132), .A4(new_n1134), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT61), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1139), .A2(KEYINPUT61), .A3(new_n1141), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1108), .A2(new_n1127), .A3(new_n1144), .A4(new_n1145), .ZN(new_n1146));
  OAI211_X1 g721(.A(new_n1141), .B(new_n633), .C1(new_n1118), .C2(new_n1117), .ZN(new_n1147));
  AND2_X1   g722(.A1(new_n1147), .A2(new_n1139), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1093), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1058), .A2(KEYINPUT62), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT62), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1055), .A2(new_n1151), .A3(new_n1057), .ZN(new_n1152));
  AND4_X1   g727(.A1(new_n1045), .A2(new_n1083), .A3(new_n1089), .A4(new_n1091), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1150), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1094), .A2(G8), .ZN(new_n1155));
  OAI21_X1  g730(.A(KEYINPUT52), .B1(new_n1155), .B2(new_n1066), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1082), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1064), .A2(new_n1074), .A3(new_n1076), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1156), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  NOR2_X1   g734(.A1(G288), .A2(G1976), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1072), .B1(new_n1158), .B2(new_n1160), .ZN(new_n1161));
  OAI22_X1  g736(.A1(new_n1159), .A2(new_n1091), .B1(new_n1161), .B2(new_n1155), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(KEYINPUT120), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT120), .ZN(new_n1164));
  OAI221_X1 g739(.A(new_n1164), .B1(new_n1161), .B2(new_n1155), .C1(new_n1159), .C2(new_n1091), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1166));
  AND2_X1   g741(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1167));
  AOI211_X1 g742(.A(new_n1063), .B(G286), .C1(new_n1053), .C2(new_n1047), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n1167), .A2(KEYINPUT63), .A3(new_n1083), .A4(new_n1168), .ZN(new_n1169));
  NAND4_X1  g744(.A1(new_n1083), .A2(new_n1168), .A3(new_n1089), .A4(new_n1091), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT63), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1169), .A2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1154), .A2(new_n1166), .A3(new_n1173), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1015), .B1(new_n1149), .B2(new_n1174), .ZN(new_n1175));
  NOR2_X1   g750(.A1(G290), .A2(G1986), .ZN(new_n1176));
  AOI21_X1  g751(.A(KEYINPUT48), .B1(new_n1001), .B2(new_n1176), .ZN(new_n1177));
  AND3_X1   g752(.A1(new_n1001), .A2(KEYINPUT48), .A3(new_n1176), .ZN(new_n1178));
  AOI211_X1 g753(.A(new_n1177), .B(new_n1178), .C1(new_n1001), .C2(new_n1013), .ZN(new_n1179));
  AOI21_X1  g754(.A(KEYINPUT46), .B1(new_n1001), .B2(new_n1007), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1000), .B1(new_n822), .B2(new_n1005), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT46), .ZN(new_n1182));
  NOR3_X1   g757(.A1(new_n1000), .A2(new_n1182), .A3(G1996), .ZN(new_n1183));
  NOR3_X1   g758(.A1(new_n1180), .A2(new_n1181), .A3(new_n1183), .ZN(new_n1184));
  XNOR2_X1  g759(.A(new_n1184), .B(KEYINPUT47), .ZN(new_n1185));
  XOR2_X1   g760(.A(new_n1011), .B(KEYINPUT127), .Z(new_n1186));
  OAI21_X1  g761(.A(new_n1003), .B1(new_n1009), .B2(new_n1186), .ZN(new_n1187));
  AOI211_X1 g762(.A(new_n1179), .B(new_n1185), .C1(new_n1001), .C2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1175), .A2(new_n1188), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g764(.A(G319), .B1(new_n670), .B2(new_n671), .ZN(new_n1191));
  NOR3_X1   g765(.A1(G229), .A2(G227), .A3(new_n1191), .ZN(new_n1192));
  NAND2_X1  g766(.A1(new_n911), .A2(new_n1192), .ZN(new_n1193));
  NOR2_X1   g767(.A1(new_n991), .A2(new_n1193), .ZN(G308));
  NAND2_X1  g768(.A1(new_n984), .A2(new_n986), .ZN(new_n1195));
  NAND2_X1  g769(.A1(new_n988), .A2(new_n990), .ZN(new_n1196));
  NAND2_X1  g770(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  NAND3_X1  g771(.A1(new_n1197), .A2(new_n911), .A3(new_n1192), .ZN(G225));
endmodule


