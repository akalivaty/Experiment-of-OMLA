//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 1 1 0 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 0 0 0 0 0 1 1 0 1 0 1 1 0 1 0 1 1 1 0 0 0 1 1 1 0 0 0 0 0 0 1 0 0 1 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n773, new_n774, new_n775, new_n777, new_n778,
    new_n779, new_n781, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n792, new_n793, new_n794, new_n796,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n857, new_n858, new_n859, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n907, new_n908, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n924, new_n925, new_n926, new_n927,
    new_n929, new_n930, new_n931, new_n932, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n947, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n961, new_n962, new_n963;
  INV_X1    g000(.A(KEYINPUT95), .ZN(new_n202));
  XNOR2_X1  g001(.A(G78gat), .B(G106gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT31), .B(G50gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  INV_X1    g004(.A(KEYINPUT29), .ZN(new_n206));
  XNOR2_X1  g005(.A(G211gat), .B(G218gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(G197gat), .B(G204gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT22), .ZN(new_n209));
  INV_X1    g008(.A(G211gat), .ZN(new_n210));
  INV_X1    g009(.A(G218gat), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n207), .A2(new_n208), .A3(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n207), .B1(new_n212), .B2(new_n208), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n206), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT3), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(G141gat), .A2(G148gat), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  NOR2_X1   g019(.A1(G141gat), .A2(G148gat), .ZN(new_n221));
  OAI21_X1  g020(.A(KEYINPUT79), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(G141gat), .ZN(new_n223));
  INV_X1    g022(.A(G148gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT79), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n225), .A2(new_n226), .A3(new_n219), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT2), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n222), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  XOR2_X1   g028(.A(G155gat), .B(G162gat), .Z(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n225), .A2(new_n219), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT80), .ZN(new_n233));
  INV_X1    g032(.A(G155gat), .ZN(new_n234));
  INV_X1    g033(.A(G162gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n228), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(G155gat), .A2(G162gat), .ZN(new_n237));
  AOI22_X1  g036(.A1(new_n232), .A2(new_n233), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n225), .A2(KEYINPUT80), .A3(new_n219), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n231), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n218), .A2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(G228gat), .ZN(new_n243));
  INV_X1    g042(.A(G233gat), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  OR2_X1    g044(.A1(new_n214), .A2(new_n215), .ZN(new_n246));
  AOI22_X1  g045(.A1(new_n229), .A2(new_n230), .B1(new_n238), .B2(new_n239), .ZN(new_n247));
  AOI21_X1  g046(.A(KEYINPUT29), .B1(new_n247), .B2(new_n217), .ZN(new_n248));
  OAI211_X1 g047(.A(new_n242), .B(new_n245), .C1(new_n246), .C2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n245), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n231), .A2(new_n240), .A3(new_n217), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n246), .B1(new_n251), .B2(new_n206), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n247), .B1(new_n217), .B2(new_n216), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n250), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n249), .A2(new_n254), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n205), .B1(new_n255), .B2(G22gat), .ZN(new_n256));
  INV_X1    g055(.A(G22gat), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n249), .A2(new_n254), .A3(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT82), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n249), .A2(new_n254), .A3(KEYINPUT82), .A4(new_n257), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n256), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(KEYINPUT83), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT83), .ZN(new_n264));
  NAND4_X1  g063(.A1(new_n256), .A2(new_n260), .A3(new_n264), .A4(new_n261), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n255), .A2(G22gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(new_n258), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(new_n205), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(G1gat), .B(G29gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n271), .B(KEYINPUT0), .ZN(new_n272));
  XNOR2_X1  g071(.A(G57gat), .B(G85gat), .ZN(new_n273));
  XOR2_X1   g072(.A(new_n272), .B(new_n273), .Z(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(G225gat), .A2(G233gat), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n277));
  XNOR2_X1  g076(.A(G113gat), .B(G120gat), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT73), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT1), .ZN(new_n281));
  INV_X1    g080(.A(G113gat), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n282), .A2(KEYINPUT73), .A3(G120gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(G127gat), .B(G134gat), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n280), .A2(new_n281), .A3(new_n283), .A4(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT72), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n282), .A2(G120gat), .ZN(new_n287));
  INV_X1    g086(.A(G120gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(G113gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(new_n281), .ZN(new_n291));
  XOR2_X1   g090(.A(G127gat), .B(G134gat), .Z(new_n292));
  AOI21_X1  g091(.A(new_n286), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(KEYINPUT1), .B1(new_n287), .B2(new_n289), .ZN(new_n294));
  NOR3_X1   g093(.A1(new_n294), .A2(KEYINPUT72), .A3(new_n284), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n285), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n277), .B1(new_n296), .B2(new_n241), .ZN(new_n297));
  OAI211_X1 g096(.A(new_n292), .B(new_n286), .C1(KEYINPUT1), .C2(new_n278), .ZN(new_n298));
  OAI21_X1  g097(.A(KEYINPUT72), .B1(new_n294), .B2(new_n284), .ZN(new_n299));
  AND3_X1   g098(.A1(new_n284), .A2(new_n281), .A3(new_n283), .ZN(new_n300));
  AOI22_X1  g099(.A1(new_n298), .A2(new_n299), .B1(new_n300), .B2(new_n280), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n301), .A2(new_n247), .A3(KEYINPUT4), .ZN(new_n302));
  AND2_X1   g101(.A1(new_n297), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n301), .B1(KEYINPUT3), .B2(new_n241), .ZN(new_n304));
  AOI21_X1  g103(.A(KEYINPUT81), .B1(new_n304), .B2(new_n251), .ZN(new_n305));
  INV_X1    g104(.A(new_n230), .ZN(new_n306));
  AOI21_X1  g105(.A(KEYINPUT2), .B1(new_n232), .B2(KEYINPUT79), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n306), .B1(new_n307), .B2(new_n227), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n233), .B1(new_n220), .B2(new_n221), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n236), .A2(new_n237), .ZN(new_n310));
  AND3_X1   g109(.A1(new_n309), .A2(new_n310), .A3(new_n239), .ZN(new_n311));
  OAI21_X1  g110(.A(KEYINPUT3), .B1(new_n308), .B2(new_n311), .ZN(new_n312));
  NAND4_X1  g111(.A1(new_n312), .A2(KEYINPUT81), .A3(new_n251), .A4(new_n296), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  OAI211_X1 g113(.A(new_n276), .B(new_n303), .C1(new_n305), .C2(new_n314), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n315), .A2(KEYINPUT5), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n296), .A2(new_n241), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n247), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n276), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(KEYINPUT5), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n297), .A2(new_n302), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n312), .A2(new_n251), .A3(new_n296), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT81), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n323), .B1(new_n326), .B2(new_n313), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n322), .B1(new_n327), .B2(new_n276), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n275), .B1(new_n316), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT6), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT5), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n327), .A2(new_n331), .A3(new_n276), .ZN(new_n332));
  INV_X1    g131(.A(new_n315), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n274), .B(new_n332), .C1(new_n333), .C2(new_n322), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n329), .A2(new_n330), .A3(new_n334), .ZN(new_n335));
  OAI211_X1 g134(.A(KEYINPUT6), .B(new_n275), .C1(new_n316), .C2(new_n328), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  XOR2_X1   g136(.A(G8gat), .B(G36gat), .Z(new_n338));
  XNOR2_X1  g137(.A(new_n338), .B(KEYINPUT78), .ZN(new_n339));
  XNOR2_X1  g138(.A(G64gat), .B(G92gat), .ZN(new_n340));
  XOR2_X1   g139(.A(new_n339), .B(new_n340), .Z(new_n341));
  NAND2_X1  g140(.A1(G226gat), .A2(G233gat), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(G183gat), .A2(G190gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(G169gat), .A2(G176gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(KEYINPUT67), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT67), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n347), .A2(G169gat), .A3(G176gat), .ZN(new_n348));
  AND2_X1   g147(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT26), .ZN(new_n350));
  INV_X1    g149(.A(G169gat), .ZN(new_n351));
  INV_X1    g150(.A(G176gat), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n350), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n344), .B1(new_n349), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT71), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n346), .A2(new_n348), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n359), .A2(new_n354), .A3(new_n353), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n360), .A2(KEYINPUT71), .A3(new_n344), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT70), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT27), .ZN(new_n364));
  INV_X1    g163(.A(G183gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(KEYINPUT68), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT68), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(G183gat), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n364), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  NOR2_X1   g168(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n363), .B1(new_n371), .B2(G190gat), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT28), .ZN(new_n373));
  INV_X1    g172(.A(G190gat), .ZN(new_n374));
  OAI211_X1 g173(.A(KEYINPUT70), .B(new_n374), .C1(new_n369), .C2(new_n370), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n372), .A2(new_n373), .A3(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(KEYINPUT27), .B(G183gat), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n377), .A2(KEYINPUT28), .A3(new_n374), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n362), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT23), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n382), .A2(new_n351), .A3(new_n352), .ZN(new_n383));
  OAI21_X1  g182(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(new_n359), .ZN(new_n386));
  NOR2_X1   g185(.A1(G183gat), .A2(G190gat), .ZN(new_n387));
  AND2_X1   g186(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n387), .B1(new_n388), .B2(G190gat), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT65), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT24), .ZN(new_n391));
  AND3_X1   g190(.A1(new_n344), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n390), .B1(new_n344), .B2(new_n391), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n389), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n386), .B1(new_n394), .B2(KEYINPUT66), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT66), .ZN(new_n396));
  OAI211_X1 g195(.A(new_n389), .B(new_n396), .C1(new_n392), .C2(new_n393), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n381), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT69), .ZN(new_n399));
  AND3_X1   g198(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n400));
  AOI21_X1  g199(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n366), .A2(new_n368), .A3(new_n374), .ZN(new_n403));
  AND2_X1   g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n385), .A2(new_n359), .A3(KEYINPUT25), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n399), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n402), .A2(new_n403), .ZN(new_n407));
  AOI22_X1  g206(.A1(new_n384), .A2(new_n383), .B1(new_n346), .B2(new_n348), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n407), .A2(new_n408), .A3(KEYINPUT69), .A4(KEYINPUT25), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n406), .A2(new_n409), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n398), .A2(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n343), .B1(new_n379), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n413), .B1(G183gat), .B2(G190gat), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n344), .A2(new_n391), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(KEYINPUT65), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n401), .A2(new_n390), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n414), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n408), .B1(new_n418), .B2(new_n396), .ZN(new_n419));
  INV_X1    g218(.A(new_n397), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n380), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n421), .A2(new_n406), .A3(new_n409), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n375), .A2(new_n373), .ZN(new_n423));
  INV_X1    g222(.A(new_n370), .ZN(new_n424));
  XNOR2_X1  g223(.A(KEYINPUT68), .B(G183gat), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n424), .B1(new_n425), .B2(new_n364), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT70), .B1(new_n426), .B2(new_n374), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n378), .B1(new_n423), .B2(new_n427), .ZN(new_n428));
  AND3_X1   g227(.A1(new_n360), .A2(KEYINPUT71), .A3(new_n344), .ZN(new_n429));
  AOI21_X1  g228(.A(KEYINPUT71), .B1(new_n360), .B2(new_n344), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n428), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(KEYINPUT29), .B1(new_n422), .B2(new_n432), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n412), .B(new_n246), .C1(new_n433), .C2(new_n343), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  AND2_X1   g234(.A1(new_n406), .A2(new_n409), .ZN(new_n436));
  AOI22_X1  g235(.A1(new_n421), .A2(new_n436), .B1(new_n428), .B2(new_n431), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n342), .B1(new_n437), .B2(KEYINPUT29), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n246), .B1(new_n438), .B2(new_n412), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n341), .B1(new_n435), .B2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n246), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n422), .A2(new_n432), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n343), .B1(new_n442), .B2(new_n206), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n437), .A2(new_n342), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n441), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n341), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n445), .A2(new_n446), .A3(new_n434), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n440), .A2(KEYINPUT30), .A3(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT30), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n445), .A2(new_n449), .A3(new_n446), .A4(new_n434), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n270), .B1(new_n337), .B2(new_n451), .ZN(new_n452));
  AND2_X1   g251(.A1(new_n266), .A2(new_n269), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n317), .A2(new_n318), .A3(new_n276), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n454), .A2(KEYINPUT85), .A3(KEYINPUT39), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(KEYINPUT39), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT85), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  OAI211_X1 g257(.A(new_n455), .B(new_n458), .C1(new_n327), .C2(new_n276), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n303), .B1(new_n305), .B2(new_n314), .ZN(new_n460));
  XNOR2_X1  g259(.A(KEYINPUT84), .B(KEYINPUT39), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n460), .A2(new_n320), .A3(new_n461), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n459), .A2(new_n462), .A3(KEYINPUT40), .A4(new_n274), .ZN(new_n463));
  AND2_X1   g262(.A1(new_n329), .A2(new_n463), .ZN(new_n464));
  AND3_X1   g263(.A1(new_n464), .A2(new_n450), .A3(new_n448), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n459), .A2(new_n462), .A3(new_n274), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT86), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n459), .A2(new_n462), .A3(KEYINPUT86), .A4(new_n274), .ZN(new_n469));
  XNOR2_X1  g268(.A(KEYINPUT87), .B(KEYINPUT40), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n453), .B1(new_n465), .B2(new_n471), .ZN(new_n472));
  AND3_X1   g271(.A1(new_n335), .A2(new_n336), .A3(new_n447), .ZN(new_n473));
  OAI21_X1  g272(.A(KEYINPUT37), .B1(new_n435), .B2(new_n439), .ZN(new_n474));
  XNOR2_X1  g273(.A(KEYINPUT88), .B(KEYINPUT37), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n445), .A2(new_n434), .A3(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n474), .A2(new_n341), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(KEYINPUT38), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT38), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n474), .A2(new_n479), .A3(new_n476), .A4(new_n341), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(KEYINPUT89), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n445), .A2(new_n434), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n446), .B1(new_n482), .B2(KEYINPUT37), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT89), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n483), .A2(new_n484), .A3(new_n479), .A4(new_n476), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n473), .A2(new_n478), .A3(new_n481), .A4(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n452), .B1(new_n472), .B2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(G227gat), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n488), .A2(new_n244), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  NOR3_X1   g289(.A1(new_n379), .A2(new_n411), .A3(new_n301), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n296), .B1(new_n422), .B2(new_n432), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  XNOR2_X1  g292(.A(KEYINPUT75), .B(KEYINPUT34), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  OAI211_X1 g295(.A(new_n490), .B(new_n494), .C1(new_n491), .C2(new_n492), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n301), .B1(new_n379), .B2(new_n411), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n422), .A2(new_n432), .A3(new_n296), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n499), .A2(new_n489), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(KEYINPUT32), .ZN(new_n502));
  XOR2_X1   g301(.A(G71gat), .B(G99gat), .Z(new_n503));
  XNOR2_X1  g302(.A(G15gat), .B(G43gat), .ZN(new_n504));
  XNOR2_X1  g303(.A(new_n503), .B(new_n504), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n499), .A2(new_n489), .A3(new_n500), .A4(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(KEYINPUT33), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT74), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n502), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n507), .A2(new_n509), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n501), .A2(KEYINPUT32), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n498), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n509), .B1(new_n506), .B2(new_n507), .ZN(new_n514));
  AND2_X1   g313(.A1(new_n501), .A2(KEYINPUT32), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n512), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  AND2_X1   g315(.A1(new_n496), .A2(new_n497), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n513), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g318(.A(KEYINPUT77), .B1(new_n519), .B2(KEYINPUT36), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n516), .A2(new_n517), .ZN(new_n521));
  OAI211_X1 g320(.A(new_n498), .B(new_n512), .C1(new_n515), .C2(new_n514), .ZN(new_n522));
  AOI21_X1  g321(.A(KEYINPUT36), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT77), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT76), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n526), .B1(new_n516), .B2(new_n517), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT36), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n528), .B1(new_n516), .B2(new_n517), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n510), .A2(KEYINPUT76), .A3(new_n498), .A4(new_n512), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n527), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n520), .A2(new_n525), .A3(new_n531), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n270), .A2(new_n521), .A3(new_n527), .A4(new_n530), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n337), .A2(new_n451), .ZN(new_n534));
  OAI21_X1  g333(.A(KEYINPUT35), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  AND2_X1   g334(.A1(new_n337), .A2(new_n451), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT35), .ZN(new_n537));
  AOI22_X1  g336(.A1(new_n266), .A2(new_n269), .B1(new_n517), .B2(new_n516), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n536), .A2(new_n537), .A3(new_n522), .A4(new_n538), .ZN(new_n539));
  AOI22_X1  g338(.A1(new_n487), .A2(new_n532), .B1(new_n535), .B2(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(G113gat), .B(G141gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n541), .B(G197gat), .ZN(new_n542));
  XOR2_X1   g341(.A(KEYINPUT11), .B(G169gat), .Z(new_n543));
  XNOR2_X1  g342(.A(new_n542), .B(new_n543), .ZN(new_n544));
  XOR2_X1   g343(.A(new_n544), .B(KEYINPUT12), .Z(new_n545));
  XNOR2_X1  g344(.A(G43gat), .B(G50gat), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n546), .A2(KEYINPUT15), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(KEYINPUT91), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n546), .A2(KEYINPUT15), .ZN(new_n549));
  NOR2_X1   g348(.A1(G29gat), .A2(G36gat), .ZN(new_n550));
  OR2_X1    g349(.A1(new_n550), .A2(KEYINPUT14), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(KEYINPUT14), .ZN(new_n552));
  XNOR2_X1  g351(.A(KEYINPUT90), .B(G29gat), .ZN(new_n553));
  INV_X1    g352(.A(G36gat), .ZN(new_n554));
  OAI211_X1 g353(.A(new_n551), .B(new_n552), .C1(new_n553), .C2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n548), .A2(new_n549), .A3(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT92), .ZN(new_n558));
  INV_X1    g357(.A(new_n549), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n558), .B1(new_n555), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g360(.A1(new_n548), .A2(new_n558), .A3(new_n549), .A4(new_n556), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(KEYINPUT17), .ZN(new_n564));
  XNOR2_X1  g363(.A(G15gat), .B(G22gat), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT16), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n565), .B1(new_n566), .B2(G1gat), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n567), .B1(G1gat), .B2(new_n565), .ZN(new_n568));
  INV_X1    g367(.A(G8gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT17), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n561), .A2(new_n571), .A3(new_n562), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n564), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT93), .ZN(new_n574));
  AND2_X1   g373(.A1(new_n561), .A2(new_n562), .ZN(new_n575));
  INV_X1    g374(.A(new_n570), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n574), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n573), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n564), .A2(new_n574), .A3(new_n570), .A4(new_n572), .ZN(new_n579));
  AOI22_X1  g378(.A1(new_n578), .A2(new_n579), .B1(G229gat), .B2(G233gat), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(KEYINPUT18), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n563), .B(new_n576), .ZN(new_n583));
  NAND2_X1  g382(.A1(G229gat), .A2(G233gat), .ZN(new_n584));
  XOR2_X1   g383(.A(new_n584), .B(KEYINPUT13), .Z(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  OR2_X1    g385(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n587), .B1(new_n580), .B2(KEYINPUT18), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n545), .B1(new_n582), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n578), .A2(new_n579), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(new_n584), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT18), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n545), .ZN(new_n594));
  NAND4_X1  g393(.A1(new_n593), .A2(new_n594), .A3(new_n581), .A4(new_n587), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT94), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n589), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  OAI211_X1 g396(.A(KEYINPUT94), .B(new_n545), .C1(new_n582), .C2(new_n588), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n202), .B1(new_n540), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n535), .A2(new_n539), .ZN(new_n601));
  INV_X1    g400(.A(new_n452), .ZN(new_n602));
  NAND4_X1  g401(.A1(new_n478), .A2(new_n336), .A3(new_n335), .A4(new_n447), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n481), .A2(new_n485), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND4_X1  g404(.A1(new_n471), .A2(new_n450), .A3(new_n464), .A4(new_n448), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(new_n270), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n602), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n531), .B1(new_n523), .B2(new_n524), .ZN(new_n609));
  AND2_X1   g408(.A1(new_n523), .A2(new_n524), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n601), .B1(new_n608), .B2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n599), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n612), .A2(KEYINPUT95), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n600), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT99), .ZN(new_n616));
  INV_X1    g415(.A(G85gat), .ZN(new_n617));
  INV_X1    g416(.A(G92gat), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(KEYINPUT99), .A2(G85gat), .A3(G92gat), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n619), .A2(KEYINPUT7), .A3(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT7), .ZN(new_n622));
  OAI211_X1 g421(.A(new_n616), .B(new_n622), .C1(new_n617), .C2(new_n618), .ZN(new_n623));
  NAND2_X1  g422(.A1(G99gat), .A2(G106gat), .ZN(new_n624));
  AOI22_X1  g423(.A1(KEYINPUT8), .A2(new_n624), .B1(new_n617), .B2(new_n618), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n621), .A2(new_n623), .A3(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(G99gat), .B(G106gat), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n626), .B(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(G64gat), .ZN(new_n631));
  AND2_X1   g430(.A1(new_n631), .A2(G57gat), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n631), .A2(G57gat), .ZN(new_n633));
  AND2_X1   g432(.A1(G71gat), .A2(G78gat), .ZN(new_n634));
  OAI22_X1  g433(.A1(new_n632), .A2(new_n633), .B1(KEYINPUT9), .B2(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(G71gat), .B(G78gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n630), .A2(KEYINPUT10), .A3(new_n637), .ZN(new_n638));
  OR2_X1    g437(.A1(new_n626), .A2(new_n628), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(KEYINPUT101), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(new_n637), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(new_n630), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n640), .A2(new_n629), .A3(new_n637), .ZN(new_n643));
  AOI21_X1  g442(.A(KEYINPUT10), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT102), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AOI211_X1 g445(.A(KEYINPUT102), .B(KEYINPUT10), .C1(new_n642), .C2(new_n643), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n638), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(G230gat), .A2(G233gat), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(G120gat), .B(G148gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(G176gat), .B(G204gat), .ZN(new_n652));
  XOR2_X1   g451(.A(new_n651), .B(new_n652), .Z(new_n653));
  INV_X1    g452(.A(new_n649), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n642), .A2(new_n654), .A3(new_n643), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  OR2_X1    g455(.A1(new_n656), .A2(KEYINPUT103), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(KEYINPUT103), .ZN(new_n658));
  NAND4_X1  g457(.A1(new_n650), .A2(new_n653), .A3(new_n657), .A4(new_n658), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n656), .B1(new_n648), .B2(new_n649), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n659), .B1(new_n660), .B2(new_n653), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(G190gat), .B(G218gat), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n564), .A2(new_n572), .A3(new_n629), .ZN(new_n665));
  AND2_X1   g464(.A1(G232gat), .A2(G233gat), .ZN(new_n666));
  AOI22_X1  g465(.A1(new_n575), .A2(new_n630), .B1(KEYINPUT41), .B2(new_n666), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n664), .B1(new_n665), .B2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n665), .A2(new_n667), .A3(new_n664), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n666), .A2(KEYINPUT41), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(G134gat), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(new_n235), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n674), .B1(new_n668), .B2(KEYINPUT100), .ZN(new_n675));
  OR2_X1    g474(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n671), .A2(new_n675), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n637), .A2(KEYINPUT21), .ZN(new_n680));
  XOR2_X1   g479(.A(G127gat), .B(G155gat), .Z(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(KEYINPUT98), .ZN(new_n682));
  XOR2_X1   g481(.A(new_n680), .B(new_n682), .Z(new_n683));
  AOI21_X1  g482(.A(new_n576), .B1(KEYINPUT21), .B2(new_n637), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(KEYINPUT97), .B(KEYINPUT19), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(KEYINPUT20), .ZN(new_n687));
  NAND2_X1  g486(.A1(G231gat), .A2(G233gat), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(KEYINPUT96), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n687), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g489(.A(G183gat), .B(G211gat), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n685), .B(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n679), .A2(new_n694), .ZN(new_n695));
  AND3_X1   g494(.A1(new_n615), .A2(new_n662), .A3(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n337), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(G1gat), .ZN(G1324gat));
  INV_X1    g498(.A(new_n451), .ZN(new_n700));
  AND2_X1   g499(.A1(new_n696), .A2(new_n700), .ZN(new_n701));
  XOR2_X1   g500(.A(KEYINPUT16), .B(G8gat), .Z(new_n702));
  AND2_X1   g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n701), .A2(new_n569), .ZN(new_n704));
  OAI21_X1  g503(.A(KEYINPUT42), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n705), .B1(KEYINPUT42), .B2(new_n703), .ZN(G1325gat));
  INV_X1    g505(.A(G15gat), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n696), .A2(new_n707), .A3(new_n519), .ZN(new_n708));
  AND2_X1   g507(.A1(new_n696), .A2(new_n611), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n708), .B1(new_n709), .B2(new_n707), .ZN(G1326gat));
  NAND2_X1  g509(.A1(new_n696), .A2(new_n453), .ZN(new_n711));
  XNOR2_X1  g510(.A(KEYINPUT43), .B(G22gat), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n711), .B(new_n712), .ZN(G1327gat));
  NAND2_X1  g512(.A1(new_n662), .A2(new_n694), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n714), .A2(new_n678), .ZN(new_n715));
  AND2_X1   g514(.A1(new_n615), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n716), .A2(new_n697), .A3(new_n553), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT45), .ZN(new_n718));
  OR2_X1    g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n717), .A2(new_n718), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT104), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n721), .A2(KEYINPUT44), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n722), .B1(new_n540), .B2(new_n678), .ZN(new_n723));
  XNOR2_X1  g522(.A(KEYINPUT104), .B(KEYINPUT44), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n612), .A2(new_n679), .A3(new_n724), .ZN(new_n725));
  AND2_X1   g524(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n599), .A2(new_n714), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n728), .A2(new_n337), .ZN(new_n729));
  OAI211_X1 g528(.A(new_n719), .B(new_n720), .C1(new_n553), .C2(new_n729), .ZN(G1328gat));
  NAND3_X1  g529(.A1(new_n716), .A2(new_n554), .A3(new_n700), .ZN(new_n731));
  OR2_X1    g530(.A1(new_n731), .A2(KEYINPUT46), .ZN(new_n732));
  OAI21_X1  g531(.A(G36gat), .B1(new_n728), .B2(new_n451), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n731), .A2(KEYINPUT46), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n732), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT105), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n735), .B(new_n736), .ZN(G1329gat));
  INV_X1    g536(.A(new_n519), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n738), .A2(G43gat), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n716), .A2(new_n739), .ZN(new_n740));
  OR2_X1    g539(.A1(new_n740), .A2(KEYINPUT107), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n726), .A2(new_n611), .A3(new_n727), .ZN(new_n742));
  AOI22_X1  g541(.A1(new_n740), .A2(KEYINPUT107), .B1(G43gat), .B2(new_n742), .ZN(new_n743));
  AOI21_X1  g542(.A(KEYINPUT106), .B1(new_n741), .B2(new_n743), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n744), .A2(KEYINPUT47), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT47), .ZN(new_n746));
  AOI211_X1 g545(.A(KEYINPUT106), .B(new_n746), .C1(new_n741), .C2(new_n743), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n745), .A2(new_n747), .ZN(G1330gat));
  NAND4_X1  g547(.A1(new_n723), .A2(new_n453), .A3(new_n725), .A4(new_n727), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(G50gat), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n270), .A2(G50gat), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n540), .A2(new_n202), .A3(new_n599), .ZN(new_n752));
  AOI21_X1  g551(.A(KEYINPUT95), .B1(new_n612), .B2(new_n613), .ZN(new_n753));
  OAI211_X1 g552(.A(new_n715), .B(new_n751), .C1(new_n752), .C2(new_n753), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n750), .A2(KEYINPUT48), .A3(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT108), .ZN(new_n756));
  AOI22_X1  g555(.A1(new_n754), .A2(new_n756), .B1(new_n749), .B2(G50gat), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n615), .A2(KEYINPUT108), .A3(new_n715), .A4(new_n751), .ZN(new_n758));
  AOI211_X1 g557(.A(KEYINPUT109), .B(KEYINPUT48), .C1(new_n757), .C2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT109), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n754), .A2(new_n756), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n761), .A2(new_n758), .A3(new_n750), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT48), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n760), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n755), .B1(new_n759), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(KEYINPUT110), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT110), .ZN(new_n767));
  OAI211_X1 g566(.A(new_n767), .B(new_n755), .C1(new_n759), .C2(new_n764), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n766), .A2(new_n768), .ZN(G1331gat));
  AND4_X1   g568(.A1(new_n612), .A2(new_n599), .A3(new_n661), .A4(new_n695), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(new_n697), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g571(.A1(new_n770), .A2(new_n700), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n773), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n774));
  XOR2_X1   g573(.A(KEYINPUT49), .B(G64gat), .Z(new_n775));
  OAI21_X1  g574(.A(new_n774), .B1(new_n773), .B2(new_n775), .ZN(G1333gat));
  NAND2_X1  g575(.A1(new_n770), .A2(new_n611), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n738), .A2(G71gat), .ZN(new_n778));
  AOI22_X1  g577(.A1(new_n777), .A2(G71gat), .B1(new_n770), .B2(new_n778), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g579(.A1(new_n770), .A2(new_n453), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g581(.A1(new_n613), .A2(new_n693), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(new_n661), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(KEYINPUT111), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(new_n726), .ZN(new_n786));
  OAI21_X1  g585(.A(G85gat), .B1(new_n786), .B2(new_n337), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n612), .A2(new_n783), .A3(new_n679), .ZN(new_n788));
  XOR2_X1   g587(.A(new_n788), .B(KEYINPUT51), .Z(new_n789));
  NAND4_X1  g588(.A1(new_n789), .A2(new_n617), .A3(new_n697), .A4(new_n661), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n787), .A2(new_n790), .ZN(G1336gat));
  OAI21_X1  g590(.A(G92gat), .B1(new_n786), .B2(new_n451), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n789), .A2(new_n618), .A3(new_n700), .A4(new_n661), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n794), .B(KEYINPUT52), .ZN(G1337gat));
  XNOR2_X1  g594(.A(KEYINPUT112), .B(G99gat), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n789), .A2(new_n519), .A3(new_n661), .A4(new_n796), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n786), .A2(new_n532), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n797), .B1(new_n798), .B2(new_n796), .ZN(G1338gat));
  INV_X1    g598(.A(KEYINPUT53), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n662), .A2(G106gat), .A3(new_n270), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n789), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n785), .A2(new_n726), .A3(new_n453), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(KEYINPUT114), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(G106gat), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n803), .A2(KEYINPUT114), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n800), .B(new_n802), .C1(new_n805), .C2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n803), .A2(G106gat), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n802), .ZN(new_n809));
  AND3_X1   g608(.A1(new_n809), .A2(KEYINPUT113), .A3(KEYINPUT53), .ZN(new_n810));
  AOI21_X1  g609(.A(KEYINPUT113), .B1(new_n809), .B2(KEYINPUT53), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n807), .B1(new_n810), .B2(new_n811), .ZN(G1339gat));
  INV_X1    g611(.A(new_n659), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n654), .B(new_n638), .C1(new_n646), .C2(new_n647), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n650), .A2(KEYINPUT54), .A3(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(new_n653), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT54), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n648), .A2(new_n817), .A3(new_n649), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n815), .A2(new_n816), .A3(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT55), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n813), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n815), .A2(KEYINPUT55), .A3(new_n816), .A4(new_n818), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n597), .A2(new_n821), .A3(new_n598), .A4(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n583), .A2(new_n586), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n824), .B1(new_n590), .B2(new_n584), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(new_n544), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n661), .A2(new_n595), .A3(new_n826), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n679), .B1(new_n823), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n821), .A2(new_n822), .ZN(new_n829));
  AND3_X1   g628(.A1(new_n595), .A2(KEYINPUT116), .A3(new_n826), .ZN(new_n830));
  AOI21_X1  g629(.A(KEYINPUT116), .B1(new_n595), .B2(new_n826), .ZN(new_n831));
  NOR4_X1   g630(.A1(new_n829), .A2(new_n830), .A3(new_n831), .A4(new_n678), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n694), .B1(new_n828), .B2(new_n832), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n599), .A2(new_n695), .A3(new_n662), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT115), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n599), .A2(new_n695), .A3(KEYINPUT115), .A4(new_n662), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n337), .B1(new_n833), .B2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(new_n533), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT117), .ZN(new_n842));
  XNOR2_X1  g641(.A(new_n841), .B(new_n842), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n843), .A2(new_n451), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n613), .A2(new_n282), .ZN(new_n845));
  XNOR2_X1  g644(.A(new_n845), .B(KEYINPUT118), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n833), .A2(new_n838), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n538), .A2(new_n522), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n700), .A2(new_n337), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n848), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(G113gat), .B1(new_n851), .B2(new_n599), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n847), .A2(new_n852), .ZN(G1340gat));
  NOR3_X1   g652(.A1(new_n851), .A2(new_n288), .A3(new_n662), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n844), .A2(new_n661), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n854), .B1(new_n855), .B2(new_n288), .ZN(G1341gat));
  INV_X1    g655(.A(G127gat), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n844), .A2(new_n857), .A3(new_n693), .ZN(new_n858));
  OAI21_X1  g657(.A(G127gat), .B1(new_n851), .B2(new_n694), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(G1342gat));
  INV_X1    g659(.A(G134gat), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n678), .A2(new_n700), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n843), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  OR2_X1    g662(.A1(new_n863), .A2(KEYINPUT56), .ZN(new_n864));
  OAI21_X1  g663(.A(G134gat), .B1(new_n851), .B2(new_n678), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n863), .A2(KEYINPUT56), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(G1343gat));
  OR2_X1    g666(.A1(new_n839), .A2(KEYINPUT119), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n611), .A2(new_n270), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n870), .B1(new_n839), .B2(KEYINPUT119), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n868), .A2(new_n451), .A3(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n223), .B1(new_n872), .B2(new_n599), .ZN(new_n873));
  AND2_X1   g672(.A1(new_n532), .A2(new_n850), .ZN(new_n874));
  AOI21_X1  g673(.A(KEYINPUT57), .B1(new_n848), .B2(new_n453), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT57), .ZN(new_n876));
  AOI211_X1 g675(.A(new_n876), .B(new_n270), .C1(new_n833), .C2(new_n838), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n874), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n613), .A2(G141gat), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n873), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT58), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  OAI211_X1 g681(.A(new_n873), .B(KEYINPUT58), .C1(new_n878), .C2(new_n879), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(G1344gat));
  INV_X1    g683(.A(KEYINPUT121), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n833), .A2(new_n834), .ZN(new_n886));
  AOI21_X1  g685(.A(KEYINPUT57), .B1(new_n886), .B2(new_n453), .ZN(new_n887));
  OAI211_X1 g686(.A(new_n661), .B(new_n874), .C1(new_n887), .C2(new_n877), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(G148gat), .ZN(new_n889));
  XOR2_X1   g688(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  OAI211_X1 g690(.A(new_n661), .B(new_n874), .C1(new_n875), .C2(new_n877), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n224), .A2(KEYINPUT59), .ZN(new_n893));
  AOI22_X1  g692(.A1(new_n889), .A2(new_n891), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n872), .A2(G148gat), .A3(new_n662), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n885), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n868), .A2(new_n871), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n897), .A2(new_n700), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n898), .A2(new_n224), .A3(new_n661), .ZN(new_n899));
  AND2_X1   g698(.A1(new_n892), .A2(new_n893), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n890), .B1(new_n888), .B2(G148gat), .ZN(new_n901));
  OAI211_X1 g700(.A(new_n899), .B(KEYINPUT121), .C1(new_n900), .C2(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n896), .A2(new_n902), .ZN(G1345gat));
  OAI21_X1  g702(.A(G155gat), .B1(new_n878), .B2(new_n694), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n693), .A2(new_n234), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n904), .B1(new_n872), .B2(new_n905), .ZN(G1346gat));
  OAI21_X1  g705(.A(G162gat), .B1(new_n878), .B2(new_n678), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n862), .A2(new_n235), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n907), .B1(new_n897), .B2(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT122), .ZN(new_n910));
  XNOR2_X1  g709(.A(new_n909), .B(new_n910), .ZN(G1347gat));
  AOI21_X1  g710(.A(new_n697), .B1(new_n833), .B2(new_n838), .ZN(new_n912));
  AND3_X1   g711(.A1(new_n912), .A2(new_n700), .A3(new_n840), .ZN(new_n913));
  AOI21_X1  g712(.A(G169gat), .B1(new_n913), .B2(new_n613), .ZN(new_n914));
  AND4_X1   g713(.A1(new_n337), .A2(new_n848), .A3(new_n700), .A4(new_n849), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n599), .A2(new_n351), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n914), .B1(new_n915), .B2(new_n916), .ZN(G1348gat));
  AOI21_X1  g716(.A(G176gat), .B1(new_n913), .B2(new_n661), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT123), .ZN(new_n919));
  OR2_X1    g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n918), .A2(new_n919), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n662), .A2(new_n352), .ZN(new_n922));
  AOI22_X1  g721(.A1(new_n920), .A2(new_n921), .B1(new_n915), .B2(new_n922), .ZN(G1349gat));
  AOI21_X1  g722(.A(new_n425), .B1(new_n915), .B2(new_n693), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n693), .A2(new_n377), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n924), .B1(new_n913), .B2(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT60), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n926), .B(new_n927), .ZN(G1350gat));
  AOI21_X1  g727(.A(new_n374), .B1(new_n915), .B2(new_n679), .ZN(new_n929));
  XOR2_X1   g728(.A(new_n929), .B(KEYINPUT61), .Z(new_n930));
  NAND3_X1  g729(.A1(new_n913), .A2(new_n374), .A3(new_n679), .ZN(new_n931));
  XOR2_X1   g730(.A(new_n931), .B(KEYINPUT124), .Z(new_n932));
  NAND2_X1  g731(.A1(new_n930), .A2(new_n932), .ZN(G1351gat));
  NAND2_X1  g732(.A1(new_n869), .A2(new_n700), .ZN(new_n934));
  INV_X1    g733(.A(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n912), .A2(new_n935), .ZN(new_n936));
  INV_X1    g735(.A(new_n936), .ZN(new_n937));
  AOI21_X1  g736(.A(G197gat), .B1(new_n937), .B2(new_n613), .ZN(new_n938));
  OR2_X1    g737(.A1(new_n887), .A2(new_n877), .ZN(new_n939));
  NOR3_X1   g738(.A1(new_n611), .A2(new_n697), .A3(new_n451), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n613), .A2(G197gat), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n938), .B1(new_n941), .B2(new_n942), .ZN(G1352gat));
  NAND2_X1  g742(.A1(new_n941), .A2(new_n661), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(G204gat), .ZN(new_n945));
  NOR3_X1   g744(.A1(new_n936), .A2(G204gat), .A3(new_n662), .ZN(new_n946));
  XNOR2_X1  g745(.A(new_n946), .B(KEYINPUT62), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n945), .A2(new_n947), .ZN(G1353gat));
  OAI211_X1 g747(.A(new_n693), .B(new_n940), .C1(new_n887), .C2(new_n877), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT126), .ZN(new_n950));
  OAI21_X1  g749(.A(G211gat), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  INV_X1    g750(.A(new_n951), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT63), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n949), .A2(new_n950), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  INV_X1    g754(.A(new_n954), .ZN(new_n956));
  OAI21_X1  g755(.A(KEYINPUT63), .B1(new_n956), .B2(new_n951), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n937), .A2(new_n210), .A3(new_n693), .ZN(new_n958));
  XNOR2_X1  g757(.A(new_n958), .B(KEYINPUT125), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n955), .A2(new_n957), .A3(new_n959), .ZN(G1354gat));
  AOI21_X1  g759(.A(G218gat), .B1(new_n937), .B2(new_n679), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n678), .A2(new_n211), .ZN(new_n962));
  XNOR2_X1  g761(.A(new_n962), .B(KEYINPUT127), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n961), .B1(new_n941), .B2(new_n963), .ZN(G1355gat));
endmodule


