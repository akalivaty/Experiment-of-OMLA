//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 0 1 0 0 1 0 0 1 0 1 1 1 0 1 1 0 0 0 1 0 1 1 0 1 0 1 0 0 0 1 0 0 0 1 1 0 1 0 0 0 0 0 1 1 1 1 0 0 0 0 0 1 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:41 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n575, new_n576, new_n578, new_n579, new_n580,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n592, new_n593, new_n594, new_n596, new_n597,
    new_n598, new_n599, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n626, new_n627, new_n629, new_n630, new_n631, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n832, new_n833, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1174, new_n1175, new_n1176;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT64), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G567), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT66), .ZN(new_n458));
  INV_X1    g033(.A(G2106), .ZN(new_n459));
  OAI21_X1  g034(.A(new_n458), .B1(new_n452), .B2(new_n459), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT67), .Z(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NAND2_X1  g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  OAI211_X1 g040(.A(G137), .B(new_n462), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G101), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT69), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n466), .A2(KEYINPUT69), .A3(new_n469), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT68), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n475), .B1(new_n464), .B2(new_n465), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT3), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(new_n467), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n478), .A2(KEYINPUT68), .A3(new_n463), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n476), .A2(new_n479), .A3(G125), .ZN(new_n480));
  NAND2_X1  g055(.A1(G113), .A2(G2104), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n462), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n474), .A2(new_n482), .ZN(G160));
  OAI21_X1  g058(.A(KEYINPUT70), .B1(G100), .B2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  NOR3_X1   g060(.A1(KEYINPUT70), .A2(G100), .A3(G2105), .ZN(new_n486));
  OAI221_X1 g061(.A(G2104), .B1(G112), .B2(new_n462), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  AOI21_X1  g062(.A(G2105), .B1(new_n478), .B2(new_n463), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G136), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n462), .B1(new_n478), .B2(new_n463), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G124), .ZN(new_n491));
  AND3_X1   g066(.A1(new_n487), .A2(new_n489), .A3(new_n491), .ZN(G162));
  NAND2_X1  g067(.A1(new_n490), .A2(G126), .ZN(new_n493));
  MUX2_X1   g068(.A(G102), .B(G114), .S(G2105), .Z(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G2104), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT71), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n488), .A2(new_n497), .A3(G138), .ZN(new_n498));
  OAI211_X1 g073(.A(G138), .B(new_n462), .C1(new_n464), .C2(new_n465), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT71), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n498), .A2(new_n500), .A3(KEYINPUT4), .ZN(new_n501));
  INV_X1    g076(.A(G138), .ZN(new_n502));
  NOR3_X1   g077(.A1(new_n502), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n476), .A2(new_n479), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n496), .B1(new_n501), .B2(new_n504), .ZN(G164));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n506), .A2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  OAI21_X1  g083(.A(KEYINPUT73), .B1(new_n508), .B2(KEYINPUT5), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT73), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n510), .A2(new_n506), .A3(G543), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n507), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n512), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT6), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n516), .A2(G651), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT72), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n518), .B1(new_n514), .B2(KEYINPUT6), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n516), .A2(KEYINPUT72), .A3(G651), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n517), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  AND3_X1   g096(.A1(new_n512), .A2(new_n521), .A3(KEYINPUT74), .ZN(new_n522));
  AOI21_X1  g097(.A(KEYINPUT74), .B1(new_n512), .B2(new_n521), .ZN(new_n523));
  INV_X1    g098(.A(G88), .ZN(new_n524));
  NOR3_X1   g099(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  AOI211_X1 g100(.A(new_n508), .B(new_n517), .C1(new_n519), .C2(new_n520), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G50), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(new_n528));
  OAI21_X1  g103(.A(KEYINPUT75), .B1(new_n525), .B2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT74), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n509), .A2(new_n511), .ZN(new_n531));
  INV_X1    g106(.A(new_n507), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(new_n517), .ZN(new_n534));
  AND3_X1   g109(.A1(new_n516), .A2(KEYINPUT72), .A3(G651), .ZN(new_n535));
  AOI21_X1  g110(.A(KEYINPUT72), .B1(new_n516), .B2(G651), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n530), .B1(new_n533), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n512), .A2(new_n521), .A3(KEYINPUT74), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n538), .A2(G88), .A3(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT75), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n540), .A2(new_n541), .A3(new_n527), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n515), .B1(new_n529), .B2(new_n542), .ZN(G166));
  NAND3_X1  g118(.A1(new_n512), .A2(G63), .A3(G651), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n521), .A2(G543), .ZN(new_n545));
  INV_X1    g120(.A(G51), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  OR2_X1    g122(.A1(new_n547), .A2(KEYINPUT76), .ZN(new_n548));
  NAND3_X1  g123(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n549));
  XOR2_X1   g124(.A(new_n549), .B(KEYINPUT7), .Z(new_n550));
  AOI21_X1  g125(.A(new_n550), .B1(new_n547), .B2(KEYINPUT76), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n522), .A2(new_n523), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G89), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n548), .A2(new_n551), .A3(new_n553), .ZN(G286));
  INV_X1    g129(.A(G286), .ZN(G168));
  NAND2_X1  g130(.A1(G77), .A2(G543), .ZN(new_n556));
  INV_X1    g131(.A(G64), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n533), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G651), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT77), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n559), .B(new_n560), .ZN(new_n561));
  XNOR2_X1  g136(.A(KEYINPUT79), .B(G90), .ZN(new_n562));
  XNOR2_X1  g137(.A(KEYINPUT78), .B(G52), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n552), .A2(new_n562), .B1(new_n526), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n561), .A2(new_n564), .ZN(G301));
  INV_X1    g140(.A(G301), .ZN(G171));
  NAND2_X1  g141(.A1(new_n552), .A2(G81), .ZN(new_n567));
  NAND2_X1  g142(.A1(G68), .A2(G543), .ZN(new_n568));
  INV_X1    g143(.A(G56), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n533), .B2(new_n569), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n570), .A2(G651), .B1(G43), .B2(new_n526), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(G860), .ZN(G153));
  AND3_X1   g149(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(G36), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n576), .B(KEYINPUT80), .ZN(G176));
  NAND2_X1  g152(.A1(G1), .A2(G3), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n578), .B(KEYINPUT8), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n575), .A2(new_n579), .ZN(new_n580));
  XOR2_X1   g155(.A(new_n580), .B(KEYINPUT81), .Z(G188));
  NAND2_X1  g156(.A1(new_n519), .A2(new_n520), .ZN(new_n582));
  NAND4_X1  g157(.A1(new_n582), .A2(G53), .A3(G543), .A4(new_n534), .ZN(new_n583));
  AND2_X1   g158(.A1(KEYINPUT82), .A2(KEYINPUT9), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n583), .B(new_n584), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n512), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n586));
  OR2_X1    g161(.A1(new_n586), .A2(new_n514), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  AND3_X1   g163(.A1(new_n538), .A2(G91), .A3(new_n539), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(G299));
  INV_X1    g166(.A(new_n515), .ZN(new_n592));
  AND3_X1   g167(.A1(new_n540), .A2(new_n541), .A3(new_n527), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n541), .B1(new_n540), .B2(new_n527), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n592), .B1(new_n593), .B2(new_n594), .ZN(G303));
  OR2_X1    g170(.A1(new_n512), .A2(G74), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n596), .A2(G651), .B1(G49), .B2(new_n526), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n538), .A2(new_n539), .ZN(new_n598));
  INV_X1    g173(.A(G87), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n597), .B1(new_n598), .B2(new_n599), .ZN(G288));
  NAND2_X1  g175(.A1(G73), .A2(G543), .ZN(new_n601));
  INV_X1    g176(.A(G61), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n533), .B2(new_n602), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n603), .A2(G651), .B1(G48), .B2(new_n526), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n538), .A2(G86), .A3(new_n539), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(G305));
  AOI22_X1  g181(.A1(new_n552), .A2(G85), .B1(G47), .B2(new_n526), .ZN(new_n607));
  AND2_X1   g182(.A1(new_n607), .A2(KEYINPUT83), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n607), .A2(KEYINPUT83), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n610));
  OAI22_X1  g185(.A1(new_n608), .A2(new_n609), .B1(new_n514), .B2(new_n610), .ZN(G290));
  INV_X1    g186(.A(KEYINPUT10), .ZN(new_n612));
  INV_X1    g187(.A(G92), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n598), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n552), .A2(KEYINPUT10), .A3(G92), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(G79), .A2(G543), .ZN(new_n617));
  INV_X1    g192(.A(G66), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n533), .B2(new_n618), .ZN(new_n619));
  AOI22_X1  g194(.A1(new_n619), .A2(G651), .B1(G54), .B2(new_n526), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n616), .A2(new_n620), .ZN(new_n621));
  MUX2_X1   g196(.A(new_n621), .B(G301), .S(G868), .Z(G284));
  XOR2_X1   g197(.A(G284), .B(KEYINPUT84), .Z(G321));
  MUX2_X1   g198(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g199(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g200(.A(new_n621), .ZN(new_n626));
  INV_X1    g201(.A(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n627), .B2(G860), .ZN(G148));
  NOR2_X1   g203(.A1(new_n621), .A2(G559), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT85), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(G868), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n631), .B1(G868), .B2(new_n573), .ZN(G323));
  XNOR2_X1  g207(.A(G323), .B(KEYINPUT11), .ZN(G282));
  MUX2_X1   g208(.A(G99), .B(G111), .S(G2105), .Z(new_n634));
  AOI22_X1  g209(.A1(G123), .A2(new_n490), .B1(new_n634), .B2(G2104), .ZN(new_n635));
  INV_X1    g210(.A(G135), .ZN(new_n636));
  INV_X1    g211(.A(new_n488), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n635), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(KEYINPUT87), .Z(new_n639));
  INV_X1    g214(.A(G2096), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n476), .A2(new_n479), .ZN(new_n642));
  INV_X1    g217(.A(new_n468), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(KEYINPUT12), .Z(new_n645));
  XOR2_X1   g220(.A(KEYINPUT86), .B(KEYINPUT13), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2100), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n645), .B(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n639), .A2(new_n640), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n641), .A2(new_n648), .A3(new_n649), .ZN(G156));
  XNOR2_X1  g225(.A(G2451), .B(G2454), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT16), .ZN(new_n652));
  XOR2_X1   g227(.A(G2443), .B(G2446), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G1341), .B(G1348), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(KEYINPUT14), .ZN(new_n657));
  XOR2_X1   g232(.A(KEYINPUT15), .B(G2435), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(G2438), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2427), .B(G2430), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT88), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n657), .B1(new_n659), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n662), .B1(new_n659), .B2(new_n661), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n656), .A2(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(G14), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n665), .B1(new_n656), .B2(new_n663), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n667), .B(KEYINPUT89), .Z(G401));
  XOR2_X1   g243(.A(G2067), .B(G2678), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT90), .ZN(new_n670));
  XOR2_X1   g245(.A(G2072), .B(G2078), .Z(new_n671));
  XOR2_X1   g246(.A(G2084), .B(G2090), .Z(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  NOR3_X1   g248(.A1(new_n670), .A2(new_n671), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT18), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n670), .A2(new_n671), .ZN(new_n676));
  XOR2_X1   g251(.A(KEYINPUT91), .B(KEYINPUT17), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n671), .B(new_n677), .ZN(new_n678));
  OAI211_X1 g253(.A(new_n676), .B(new_n673), .C1(new_n670), .C2(new_n678), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n678), .A2(new_n670), .A3(new_n672), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n675), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(new_n640), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(G2100), .ZN(G227));
  XOR2_X1   g258(.A(G1971), .B(G1976), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT19), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1956), .B(G2474), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1961), .B(G1966), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  AND2_X1   g263(.A1(new_n686), .A2(new_n687), .ZN(new_n689));
  NOR3_X1   g264(.A1(new_n685), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n685), .A2(new_n688), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n691), .B(KEYINPUT20), .Z(new_n692));
  AOI211_X1 g267(.A(new_n690), .B(new_n692), .C1(new_n685), .C2(new_n689), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT92), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n693), .B(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1991), .B(G1996), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1981), .B(G1986), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n696), .B(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(G229));
  MUX2_X1   g276(.A(G6), .B(G305), .S(G16), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT94), .ZN(new_n703));
  XOR2_X1   g278(.A(KEYINPUT32), .B(G1981), .Z(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  NOR2_X1   g280(.A1(G16), .A2(G23), .ZN(new_n706));
  INV_X1    g281(.A(G288), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n706), .B1(new_n707), .B2(G16), .ZN(new_n708));
  XOR2_X1   g283(.A(KEYINPUT33), .B(G1976), .Z(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(KEYINPUT95), .Z(new_n710));
  XNOR2_X1  g285(.A(new_n708), .B(new_n710), .ZN(new_n711));
  NOR2_X1   g286(.A1(G16), .A2(G22), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(G166), .B2(G16), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n711), .B1(G1971), .B2(new_n713), .ZN(new_n714));
  OAI211_X1 g289(.A(new_n705), .B(new_n714), .C1(G1971), .C2(new_n713), .ZN(new_n715));
  OR2_X1    g290(.A1(new_n715), .A2(KEYINPUT34), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n715), .A2(KEYINPUT34), .ZN(new_n717));
  MUX2_X1   g292(.A(G95), .B(G107), .S(G2105), .Z(new_n718));
  AOI22_X1  g293(.A1(G119), .A2(new_n490), .B1(new_n718), .B2(G2104), .ZN(new_n719));
  INV_X1    g294(.A(G131), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n719), .B1(new_n720), .B2(new_n637), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT93), .Z(new_n722));
  MUX2_X1   g297(.A(G25), .B(new_n722), .S(G29), .Z(new_n723));
  XOR2_X1   g298(.A(KEYINPUT35), .B(G1991), .Z(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(G290), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(G16), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(G16), .B2(G24), .ZN(new_n728));
  INV_X1    g303(.A(G1986), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n725), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(new_n729), .B2(new_n728), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n716), .A2(new_n717), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(KEYINPUT36), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT36), .ZN(new_n734));
  NAND4_X1  g309(.A1(new_n716), .A2(new_n734), .A3(new_n717), .A4(new_n731), .ZN(new_n735));
  NOR2_X1   g310(.A1(G16), .A2(G21), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(G168), .B2(G16), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT102), .ZN(new_n738));
  AND2_X1   g313(.A1(new_n738), .A2(G1966), .ZN(new_n739));
  INV_X1    g314(.A(G16), .ZN(new_n740));
  NOR2_X1   g315(.A1(G171), .A2(new_n740), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(G5), .B2(new_n740), .ZN(new_n742));
  INV_X1    g317(.A(G1961), .ZN(new_n743));
  AND2_X1   g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n639), .A2(G29), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT103), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n488), .A2(G139), .ZN(new_n747));
  OR2_X1    g322(.A1(new_n747), .A2(KEYINPUT98), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n747), .A2(KEYINPUT98), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT25), .ZN(new_n750));
  INV_X1    g325(.A(G103), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n750), .B1(new_n643), .B2(new_n751), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n468), .A2(KEYINPUT25), .A3(G103), .ZN(new_n753));
  AOI22_X1  g328(.A1(new_n748), .A2(new_n749), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  AND2_X1   g329(.A1(new_n476), .A2(new_n479), .ZN(new_n755));
  AOI22_X1  g330(.A1(new_n755), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n754), .B1(new_n462), .B2(new_n756), .ZN(new_n757));
  MUX2_X1   g332(.A(G33), .B(new_n757), .S(G29), .Z(new_n758));
  NOR2_X1   g333(.A1(G29), .A2(G35), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(G162), .B2(G29), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT29), .Z(new_n761));
  INV_X1    g336(.A(G2090), .ZN(new_n762));
  AOI22_X1  g337(.A1(G2072), .A2(new_n758), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  OAI211_X1 g338(.A(new_n746), .B(new_n763), .C1(G2072), .C2(new_n758), .ZN(new_n764));
  NAND2_X1  g339(.A1(G160), .A2(G29), .ZN(new_n765));
  INV_X1    g340(.A(G29), .ZN(new_n766));
  AND2_X1   g341(.A1(KEYINPUT24), .A2(G34), .ZN(new_n767));
  NOR2_X1   g342(.A1(KEYINPUT24), .A2(G34), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n766), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n765), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT99), .ZN(new_n771));
  OAI22_X1  g346(.A1(new_n742), .A2(new_n743), .B1(G2084), .B2(new_n771), .ZN(new_n772));
  NOR4_X1   g347(.A1(new_n739), .A2(new_n744), .A3(new_n764), .A4(new_n772), .ZN(new_n773));
  NOR2_X1   g348(.A1(G16), .A2(G19), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(new_n573), .B2(G16), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT96), .Z(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(G1341), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n771), .A2(G2084), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT100), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n738), .A2(G1966), .ZN(new_n780));
  NOR3_X1   g355(.A1(new_n777), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT31), .B(G11), .ZN(new_n782));
  XOR2_X1   g357(.A(KEYINPUT30), .B(G28), .Z(new_n783));
  OAI21_X1  g358(.A(new_n782), .B1(new_n783), .B2(G29), .ZN(new_n784));
  AOI22_X1  g359(.A1(G129), .A2(new_n490), .B1(new_n488), .B2(G141), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n468), .A2(G105), .ZN(new_n786));
  NAND3_X1  g361(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT26), .Z(new_n788));
  NAND3_X1  g363(.A1(new_n785), .A2(new_n786), .A3(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n790), .A2(new_n766), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(new_n766), .B2(G32), .ZN(new_n792));
  XOR2_X1   g367(.A(KEYINPUT27), .B(G1996), .Z(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT101), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n784), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(new_n794), .B2(new_n792), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n761), .A2(new_n762), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g373(.A1(G4), .A2(G16), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(new_n626), .B2(G16), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n800), .A2(G1348), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n766), .A2(G26), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT28), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n488), .A2(G140), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n490), .A2(G128), .ZN(new_n805));
  AND2_X1   g380(.A1(G116), .A2(G2105), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(G104), .B2(new_n462), .ZN(new_n807));
  OAI211_X1 g382(.A(new_n804), .B(new_n805), .C1(new_n467), .C2(new_n807), .ZN(new_n808));
  AND3_X1   g383(.A1(new_n808), .A2(KEYINPUT97), .A3(G29), .ZN(new_n809));
  AOI21_X1  g384(.A(KEYINPUT97), .B1(new_n808), .B2(G29), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n803), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(G2067), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NOR2_X1   g388(.A1(G27), .A2(G29), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(G164), .B2(G29), .ZN(new_n815));
  INV_X1    g390(.A(G2078), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  NAND4_X1  g392(.A1(new_n798), .A2(new_n801), .A3(new_n813), .A4(new_n817), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n800), .A2(G1348), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n740), .A2(G20), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT105), .ZN(new_n821));
  XNOR2_X1  g396(.A(KEYINPUT104), .B(KEYINPUT23), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n823), .B1(G299), .B2(G16), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(G1956), .Z(new_n825));
  NOR3_X1   g400(.A1(new_n818), .A2(new_n819), .A3(new_n825), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n773), .A2(new_n781), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n827), .A2(KEYINPUT106), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT106), .ZN(new_n829));
  NAND4_X1  g404(.A1(new_n773), .A2(new_n781), .A3(new_n829), .A4(new_n826), .ZN(new_n830));
  AOI22_X1  g405(.A1(new_n733), .A2(new_n735), .B1(new_n828), .B2(new_n830), .ZN(G311));
  NAND2_X1  g406(.A1(new_n733), .A2(new_n735), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n828), .A2(new_n830), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(G150));
  NAND2_X1  g409(.A1(new_n626), .A2(G559), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT38), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n572), .A2(KEYINPUT107), .ZN(new_n837));
  INV_X1    g412(.A(G93), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n598), .A2(new_n838), .ZN(new_n839));
  AOI22_X1  g414(.A1(new_n512), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n840));
  INV_X1    g415(.A(G55), .ZN(new_n841));
  OAI22_X1  g416(.A1(new_n840), .A2(new_n514), .B1(new_n841), .B2(new_n545), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT108), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n837), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT107), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n846), .B1(new_n567), .B2(new_n571), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n839), .A2(new_n842), .ZN(new_n848));
  OAI21_X1  g423(.A(KEYINPUT108), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n572), .A2(KEYINPUT107), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n845), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n850), .B1(new_n845), .B2(new_n849), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n836), .B(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT39), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT109), .ZN(new_n859));
  AOI21_X1  g434(.A(G860), .B1(new_n856), .B2(new_n857), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n843), .A2(G860), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT110), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT37), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n861), .A2(new_n864), .ZN(G145));
  XNOR2_X1  g440(.A(new_n645), .B(new_n721), .ZN(new_n866));
  MUX2_X1   g441(.A(G106), .B(G118), .S(G2105), .Z(new_n867));
  AOI22_X1  g442(.A1(G130), .A2(new_n490), .B1(new_n867), .B2(G2104), .ZN(new_n868));
  INV_X1    g443(.A(G142), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n868), .B1(new_n869), .B2(new_n637), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n866), .B(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(G164), .B(new_n808), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n871), .B(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n757), .B(new_n790), .ZN(new_n874));
  OR2_X1    g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n873), .A2(new_n874), .ZN(new_n876));
  XOR2_X1   g451(.A(G160), .B(G162), .Z(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(new_n639), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n875), .A2(new_n876), .A3(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(G37), .ZN(new_n881));
  AND2_X1   g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n879), .B1(new_n875), .B2(new_n876), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n882), .A2(KEYINPUT40), .A3(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT40), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n880), .A2(new_n881), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n886), .B1(new_n887), .B2(new_n883), .ZN(new_n888));
  AND2_X1   g463(.A1(new_n885), .A2(new_n888), .ZN(G395));
  NOR2_X1   g464(.A1(new_n843), .A2(G868), .ZN(new_n890));
  XNOR2_X1  g465(.A(G166), .B(G305), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(G290), .A2(G288), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  NOR2_X1   g469(.A1(G290), .A2(G288), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n892), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n895), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n897), .A2(new_n893), .A3(new_n891), .ZN(new_n898));
  AND2_X1   g473(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(KEYINPUT111), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT41), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n621), .A2(G299), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n621), .A2(G299), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n901), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n626), .A2(new_n590), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n906), .A2(KEYINPUT41), .A3(new_n902), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n854), .A2(new_n630), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n854), .A2(new_n630), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n908), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n911), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n903), .A2(new_n904), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n913), .A2(new_n915), .A3(new_n909), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n912), .A2(new_n916), .A3(KEYINPUT42), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(KEYINPUT42), .B1(new_n912), .B2(new_n916), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n900), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n912), .A2(new_n916), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT42), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n923), .A2(KEYINPUT111), .A3(new_n899), .A4(new_n917), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n920), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n890), .B1(new_n925), .B2(G868), .ZN(G295));
  AOI21_X1  g501(.A(new_n890), .B1(new_n925), .B2(G868), .ZN(G331));
  XNOR2_X1  g502(.A(G301), .B(G286), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n928), .B1(new_n852), .B2(new_n853), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n845), .A2(new_n849), .ZN(new_n930));
  INV_X1    g505(.A(new_n850), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  XNOR2_X1  g507(.A(G301), .B(G168), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n932), .A2(new_n933), .A3(new_n851), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n929), .A2(new_n934), .A3(new_n914), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n908), .B1(new_n929), .B2(new_n934), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n896), .A2(new_n898), .ZN(new_n938));
  NOR3_X1   g513(.A1(new_n936), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n929), .A2(new_n934), .ZN(new_n940));
  AND2_X1   g515(.A1(new_n905), .A2(new_n907), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n899), .B1(new_n942), .B2(new_n935), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n881), .B1(new_n939), .B2(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n944), .A2(KEYINPUT114), .A3(KEYINPUT43), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT114), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n938), .B1(new_n936), .B2(new_n937), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n942), .A2(new_n899), .A3(new_n935), .ZN(new_n948));
  AOI21_X1  g523(.A(G37), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT43), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n946), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  OAI211_X1 g526(.A(KEYINPUT113), .B(new_n899), .C1(new_n936), .C2(new_n937), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT113), .ZN(new_n953));
  OAI211_X1 g528(.A(new_n942), .B(new_n935), .C1(new_n953), .C2(new_n938), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n952), .A2(new_n954), .A3(new_n950), .A4(new_n881), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n945), .A2(new_n951), .A3(KEYINPUT44), .A4(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n952), .A2(new_n954), .A3(new_n881), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(KEYINPUT43), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n949), .A2(new_n950), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  XOR2_X1   g535(.A(KEYINPUT112), .B(KEYINPUT44), .Z(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n956), .A2(new_n962), .ZN(G397));
  OAI21_X1  g538(.A(KEYINPUT4), .B1(new_n499), .B2(KEYINPUT71), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n497), .B1(new_n488), .B2(G138), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n504), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(new_n496), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  XNOR2_X1  g543(.A(KEYINPUT115), .B(G1384), .ZN(new_n969));
  AOI21_X1  g544(.A(KEYINPUT45), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(G40), .ZN(new_n971));
  NOR3_X1   g546(.A1(new_n474), .A2(new_n482), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(G1996), .ZN(new_n974));
  NOR3_X1   g549(.A1(new_n973), .A2(new_n974), .A3(new_n790), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n975), .B(KEYINPUT116), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n973), .A2(G1996), .ZN(new_n977));
  INV_X1    g552(.A(new_n973), .ZN(new_n978));
  XNOR2_X1  g553(.A(new_n808), .B(G2067), .ZN(new_n979));
  AOI22_X1  g554(.A1(new_n977), .A2(new_n790), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n721), .B(new_n724), .ZN(new_n981));
  OAI211_X1 g556(.A(new_n976), .B(new_n980), .C1(new_n973), .C2(new_n981), .ZN(new_n982));
  XNOR2_X1  g557(.A(G290), .B(G1986), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n982), .B1(new_n978), .B2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(G8), .ZN(new_n985));
  AOI21_X1  g560(.A(G1384), .B1(new_n966), .B2(new_n967), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n985), .B1(new_n972), .B2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT49), .ZN(new_n988));
  INV_X1    g563(.A(G1981), .ZN(new_n989));
  AND3_X1   g564(.A1(new_n604), .A2(new_n989), .A3(new_n605), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n989), .B1(new_n604), .B2(new_n605), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n988), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(G305), .A2(G1981), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n604), .A2(new_n989), .A3(new_n605), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n993), .A2(KEYINPUT49), .A3(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n992), .A2(new_n995), .A3(new_n987), .ZN(new_n996));
  INV_X1    g571(.A(G1976), .ZN(new_n997));
  AND3_X1   g572(.A1(new_n996), .A2(new_n997), .A3(new_n707), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n987), .B1(new_n998), .B2(new_n990), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n987), .B1(new_n997), .B2(G288), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(KEYINPUT52), .ZN(new_n1001));
  AOI21_X1  g576(.A(KEYINPUT52), .B1(G288), .B2(new_n997), .ZN(new_n1002));
  OAI211_X1 g577(.A(new_n1002), .B(new_n987), .C1(new_n997), .C2(G288), .ZN(new_n1003));
  AND3_X1   g578(.A1(new_n1001), .A2(new_n996), .A3(new_n1003), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n972), .B1(new_n986), .B2(KEYINPUT45), .ZN(new_n1005));
  AND3_X1   g580(.A1(new_n968), .A2(KEYINPUT45), .A3(new_n969), .ZN(new_n1006));
  OAI21_X1  g581(.A(KEYINPUT117), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(G1971), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT45), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1009), .B1(G164), .B2(G1384), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n968), .A2(KEYINPUT45), .A3(new_n969), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT117), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1010), .A2(new_n1011), .A3(new_n1012), .A4(new_n972), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1007), .A2(new_n1008), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n480), .A2(new_n481), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(G2105), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1016), .A2(G40), .A3(new_n472), .A4(new_n473), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n986), .A2(KEYINPUT50), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT50), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1019), .B1(G164), .B2(G1384), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1017), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(new_n762), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n985), .B1(new_n1014), .B2(new_n1022), .ZN(new_n1023));
  XOR2_X1   g598(.A(KEYINPUT118), .B(KEYINPUT55), .Z(new_n1024));
  NOR3_X1   g599(.A1(G166), .A2(new_n985), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1024), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1026), .B1(G303), .B2(G8), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1004), .A2(new_n1023), .A3(new_n1028), .ZN(new_n1029));
  AND2_X1   g604(.A1(new_n999), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1014), .A2(new_n1022), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(G8), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1028), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1023), .A2(new_n1028), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n986), .A2(KEYINPUT45), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1036), .A2(new_n1010), .A3(new_n972), .ZN(new_n1037));
  INV_X1    g612(.A(G1966), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1040));
  INV_X1    g615(.A(G2084), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1040), .A2(new_n1041), .A3(new_n972), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1039), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(G8), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1044), .A2(G286), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1034), .A2(new_n1035), .A3(new_n1004), .A4(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1030), .B1(new_n1046), .B2(KEYINPUT63), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT63), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1004), .B1(new_n1023), .B2(new_n1028), .ZN(new_n1049));
  AND3_X1   g624(.A1(new_n1031), .A2(new_n1028), .A3(G8), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1048), .B1(new_n1051), .B2(new_n1045), .ZN(new_n1052));
  OAI21_X1  g627(.A(KEYINPUT119), .B1(new_n1047), .B2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1051), .A2(new_n1048), .A3(new_n1045), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1046), .A2(KEYINPUT63), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT119), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1054), .A2(new_n1055), .A3(new_n1056), .A4(new_n1030), .ZN(new_n1057));
  AND2_X1   g632(.A1(new_n1053), .A2(new_n1057), .ZN(new_n1058));
  XOR2_X1   g633(.A(KEYINPUT56), .B(G2072), .Z(new_n1059));
  INV_X1    g634(.A(new_n1059), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1010), .A2(new_n1011), .A3(new_n972), .A4(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1061), .B1(new_n1021), .B2(G1956), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT57), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1063), .B1(new_n588), .B2(new_n589), .ZN(new_n1064));
  INV_X1    g639(.A(new_n589), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1065), .A2(KEYINPUT57), .A3(new_n585), .A4(new_n587), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1062), .A2(new_n1064), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT121), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n972), .A2(new_n986), .ZN(new_n1069));
  OAI22_X1  g644(.A1(new_n1021), .A2(G1348), .B1(G2067), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(new_n626), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT60), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n1068), .B(KEYINPUT61), .C1(new_n1071), .C2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1066), .A2(new_n1064), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n1074), .B(new_n1061), .C1(new_n1021), .C2(G1956), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1073), .A2(new_n1076), .ZN(new_n1077));
  AND3_X1   g652(.A1(new_n1075), .A2(new_n1068), .A3(KEYINPUT61), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n621), .A2(KEYINPUT60), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n626), .A2(new_n1072), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1070), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1071), .B1(new_n1078), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1077), .A2(new_n1082), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1076), .A2(new_n1071), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT120), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1010), .A2(new_n1011), .A3(new_n974), .A4(new_n972), .ZN(new_n1086));
  XOR2_X1   g661(.A(KEYINPUT58), .B(G1341), .Z(new_n1087));
  NAND2_X1  g662(.A1(new_n1069), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1085), .B1(new_n1089), .B2(new_n573), .ZN(new_n1090));
  AOI211_X1 g665(.A(KEYINPUT120), .B(new_n572), .C1(new_n1086), .C2(new_n1088), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(KEYINPUT59), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT59), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1094), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1084), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1067), .B1(new_n1083), .B2(new_n1096), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1021), .A2(G1961), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n816), .A2(KEYINPUT53), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1037), .A2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(G2078), .B1(new_n1007), .B2(new_n1013), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1101), .B1(KEYINPUT53), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(G171), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1017), .A2(new_n1099), .ZN(new_n1105));
  AND2_X1   g680(.A1(new_n1105), .A2(new_n1011), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT123), .ZN(new_n1107));
  INV_X1    g682(.A(new_n970), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1106), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1105), .A2(new_n1011), .ZN(new_n1110));
  OAI21_X1  g685(.A(KEYINPUT123), .B1(new_n1110), .B2(new_n970), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1098), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1112), .B1(KEYINPUT53), .B2(new_n1102), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1104), .B1(G171), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT54), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n985), .B1(new_n1039), .B2(new_n1042), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT51), .ZN(new_n1117));
  NOR2_X1   g692(.A1(G168), .A2(new_n985), .ZN(new_n1118));
  NOR4_X1   g693(.A1(new_n1116), .A2(KEYINPUT122), .A3(new_n1117), .A4(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1116), .A2(G286), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1120), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT122), .ZN(new_n1123));
  OAI21_X1  g698(.A(KEYINPUT51), .B1(new_n1116), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1118), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1044), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  AOI22_X1  g702(.A1(new_n1114), .A2(new_n1115), .B1(new_n1122), .B2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1107), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1129));
  NOR3_X1   g704(.A1(new_n1110), .A2(KEYINPUT123), .A3(new_n970), .ZN(new_n1130));
  OAI22_X1  g705(.A1(new_n1129), .A2(new_n1130), .B1(G1961), .B2(new_n1021), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1007), .A2(new_n1013), .ZN(new_n1132));
  AOI21_X1  g707(.A(KEYINPUT53), .B1(new_n1132), .B2(new_n816), .ZN(new_n1133));
  OAI21_X1  g708(.A(G171), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1134));
  OAI211_X1 g709(.A(new_n1101), .B(G301), .C1(KEYINPUT53), .C2(new_n1102), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1134), .A2(KEYINPUT54), .A3(new_n1135), .ZN(new_n1136));
  AND2_X1   g711(.A1(new_n1136), .A2(new_n1051), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1097), .A2(new_n1128), .A3(new_n1137), .ZN(new_n1138));
  NOR3_X1   g713(.A1(new_n1104), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT124), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT62), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1044), .A2(new_n1123), .A3(KEYINPUT51), .A4(new_n1125), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1127), .A2(new_n1141), .A3(new_n1142), .A4(new_n1120), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1139), .A2(new_n1140), .A3(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1122), .A2(new_n1127), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(KEYINPUT62), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1140), .B1(new_n1139), .B2(new_n1143), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1138), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n984), .B1(new_n1058), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n724), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n722), .A2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n976), .A2(new_n980), .A3(new_n1152), .ZN(new_n1153));
  OR2_X1    g728(.A1(new_n808), .A2(G2067), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n973), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT125), .ZN(new_n1156));
  OR2_X1    g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1158));
  NOR3_X1   g733(.A1(G290), .A2(G1986), .A3(new_n973), .ZN(new_n1159));
  XNOR2_X1  g734(.A(new_n1159), .B(KEYINPUT48), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n982), .A2(new_n1160), .ZN(new_n1161));
  OR2_X1    g736(.A1(new_n977), .A2(KEYINPUT46), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n977), .A2(KEYINPUT46), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n978), .B1(new_n789), .B2(new_n979), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1162), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  XOR2_X1   g740(.A(KEYINPUT126), .B(KEYINPUT47), .Z(new_n1166));
  XNOR2_X1  g741(.A(new_n1165), .B(new_n1166), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1161), .A2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1157), .A2(new_n1158), .A3(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT127), .ZN(new_n1170));
  XNOR2_X1  g745(.A(new_n1169), .B(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1150), .A2(new_n1171), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g747(.A1(new_n882), .A2(new_n884), .ZN(new_n1174));
  INV_X1    g748(.A(new_n667), .ZN(new_n1175));
  NOR4_X1   g749(.A1(G229), .A2(new_n460), .A3(new_n1175), .A4(G227), .ZN(new_n1176));
  AND3_X1   g750(.A1(new_n1174), .A2(new_n960), .A3(new_n1176), .ZN(G308));
  NAND3_X1  g751(.A1(new_n1174), .A2(new_n960), .A3(new_n1176), .ZN(G225));
endmodule


