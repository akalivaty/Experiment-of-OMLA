

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584;

  XNOR2_X1 U322 ( .A(n378), .B(n377), .ZN(n380) );
  XNOR2_X1 U323 ( .A(n394), .B(KEYINPUT68), .ZN(n303) );
  XNOR2_X1 U324 ( .A(n368), .B(n367), .ZN(n369) );
  INV_X1 U325 ( .A(KEYINPUT47), .ZN(n424) );
  XNOR2_X1 U326 ( .A(n370), .B(n369), .ZN(n372) );
  XNOR2_X1 U327 ( .A(n376), .B(n375), .ZN(n377) );
  NOR2_X1 U328 ( .A1(n538), .A2(n447), .ZN(n457) );
  INV_X1 U329 ( .A(KEYINPUT69), .ZN(n301) );
  XNOR2_X1 U330 ( .A(n302), .B(n301), .ZN(n394) );
  XNOR2_X1 U331 ( .A(n449), .B(n448), .ZN(n578) );
  XNOR2_X1 U332 ( .A(n308), .B(n307), .ZN(n567) );
  XOR2_X1 U333 ( .A(n361), .B(n360), .Z(n538) );
  XNOR2_X1 U334 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U335 ( .A(n455), .B(n454), .ZN(G1352GAT) );
  NAND2_X1 U336 ( .A1(G229GAT), .A2(G233GAT), .ZN(n295) );
  XOR2_X1 U337 ( .A(G141GAT), .B(G197GAT), .Z(n291) );
  XNOR2_X1 U338 ( .A(G169GAT), .B(G113GAT), .ZN(n290) );
  XNOR2_X1 U339 ( .A(n291), .B(n290), .ZN(n293) );
  XOR2_X1 U340 ( .A(G36GAT), .B(G50GAT), .Z(n292) );
  XNOR2_X1 U341 ( .A(n293), .B(n292), .ZN(n294) );
  XNOR2_X1 U342 ( .A(n295), .B(n294), .ZN(n308) );
  XOR2_X1 U343 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n297) );
  XNOR2_X1 U344 ( .A(G22GAT), .B(G8GAT), .ZN(n296) );
  XNOR2_X1 U345 ( .A(n297), .B(n296), .ZN(n306) );
  XNOR2_X1 U346 ( .A(G15GAT), .B(G1GAT), .ZN(n298) );
  XNOR2_X1 U347 ( .A(n298), .B(KEYINPUT70), .ZN(n402) );
  XOR2_X1 U348 ( .A(n402), .B(KEYINPUT67), .Z(n304) );
  XOR2_X1 U349 ( .A(KEYINPUT8), .B(KEYINPUT7), .Z(n300) );
  XNOR2_X1 U350 ( .A(G43GAT), .B(G29GAT), .ZN(n299) );
  XNOR2_X1 U351 ( .A(n300), .B(n299), .ZN(n302) );
  XNOR2_X1 U352 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U353 ( .A(n306), .B(n305), .Z(n307) );
  XOR2_X1 U354 ( .A(G22GAT), .B(G155GAT), .Z(n403) );
  XOR2_X1 U355 ( .A(KEYINPUT3), .B(KEYINPUT92), .Z(n310) );
  XNOR2_X1 U356 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n309) );
  XNOR2_X1 U357 ( .A(n310), .B(n309), .ZN(n357) );
  XOR2_X1 U358 ( .A(n403), .B(n357), .Z(n312) );
  NAND2_X1 U359 ( .A1(G228GAT), .A2(G233GAT), .ZN(n311) );
  XNOR2_X1 U360 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U361 ( .A(n313), .B(KEYINPUT22), .Z(n317) );
  XOR2_X1 U362 ( .A(G162GAT), .B(KEYINPUT79), .Z(n315) );
  XNOR2_X1 U363 ( .A(G50GAT), .B(G218GAT), .ZN(n314) );
  XNOR2_X1 U364 ( .A(n315), .B(n314), .ZN(n388) );
  XNOR2_X1 U365 ( .A(n388), .B(KEYINPUT93), .ZN(n316) );
  XNOR2_X1 U366 ( .A(n317), .B(n316), .ZN(n321) );
  XOR2_X1 U367 ( .A(KEYINPUT24), .B(KEYINPUT90), .Z(n319) );
  XNOR2_X1 U368 ( .A(G106GAT), .B(KEYINPUT23), .ZN(n318) );
  XNOR2_X1 U369 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U370 ( .A(n321), .B(n320), .Z(n327) );
  XOR2_X1 U371 ( .A(G211GAT), .B(KEYINPUT91), .Z(n323) );
  XNOR2_X1 U372 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n322) );
  XNOR2_X1 U373 ( .A(n323), .B(n322), .ZN(n434) );
  XOR2_X1 U374 ( .A(G78GAT), .B(G148GAT), .Z(n325) );
  XNOR2_X1 U375 ( .A(KEYINPUT75), .B(G204GAT), .ZN(n324) );
  XNOR2_X1 U376 ( .A(n325), .B(n324), .ZN(n375) );
  XNOR2_X1 U377 ( .A(n434), .B(n375), .ZN(n326) );
  XNOR2_X1 U378 ( .A(n327), .B(n326), .ZN(n476) );
  XOR2_X1 U379 ( .A(G176GAT), .B(G183GAT), .Z(n329) );
  XNOR2_X1 U380 ( .A(G43GAT), .B(KEYINPUT20), .ZN(n328) );
  XNOR2_X1 U381 ( .A(n329), .B(n328), .ZN(n343) );
  XOR2_X1 U382 ( .A(KEYINPUT64), .B(KEYINPUT89), .Z(n331) );
  NAND2_X1 U383 ( .A1(G227GAT), .A2(G233GAT), .ZN(n330) );
  XNOR2_X1 U384 ( .A(n331), .B(n330), .ZN(n334) );
  XOR2_X1 U385 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n333) );
  XNOR2_X1 U386 ( .A(G169GAT), .B(KEYINPUT19), .ZN(n332) );
  XNOR2_X1 U387 ( .A(n333), .B(n332), .ZN(n439) );
  XOR2_X1 U388 ( .A(n334), .B(n439), .Z(n338) );
  XOR2_X1 U389 ( .A(G127GAT), .B(KEYINPUT0), .Z(n336) );
  XNOR2_X1 U390 ( .A(G113GAT), .B(G134GAT), .ZN(n335) );
  XNOR2_X1 U391 ( .A(n336), .B(n335), .ZN(n345) );
  XNOR2_X1 U392 ( .A(G15GAT), .B(n345), .ZN(n337) );
  XNOR2_X1 U393 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U394 ( .A(G120GAT), .B(G71GAT), .Z(n362) );
  XOR2_X1 U395 ( .A(n339), .B(n362), .Z(n341) );
  XNOR2_X1 U396 ( .A(G99GAT), .B(G190GAT), .ZN(n340) );
  XNOR2_X1 U397 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U398 ( .A(n343), .B(n342), .ZN(n459) );
  INV_X1 U399 ( .A(n459), .ZN(n540) );
  NOR2_X1 U400 ( .A1(n476), .A2(n540), .ZN(n344) );
  XNOR2_X1 U401 ( .A(n344), .B(KEYINPUT26), .ZN(n471) );
  XOR2_X1 U402 ( .A(n345), .B(G1GAT), .Z(n347) );
  NAND2_X1 U403 ( .A1(G225GAT), .A2(G233GAT), .ZN(n346) );
  XNOR2_X1 U404 ( .A(n347), .B(n346), .ZN(n361) );
  XOR2_X1 U405 ( .A(G85GAT), .B(G162GAT), .Z(n349) );
  XNOR2_X1 U406 ( .A(G29GAT), .B(G120GAT), .ZN(n348) );
  XNOR2_X1 U407 ( .A(n349), .B(n348), .ZN(n353) );
  XOR2_X1 U408 ( .A(KEYINPUT94), .B(G57GAT), .Z(n351) );
  XNOR2_X1 U409 ( .A(KEYINPUT1), .B(KEYINPUT5), .ZN(n350) );
  XNOR2_X1 U410 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U411 ( .A(n353), .B(n352), .Z(n359) );
  XOR2_X1 U412 ( .A(KEYINPUT6), .B(KEYINPUT4), .Z(n355) );
  XNOR2_X1 U413 ( .A(G148GAT), .B(G155GAT), .ZN(n354) );
  XNOR2_X1 U414 ( .A(n355), .B(n354), .ZN(n356) );
  XNOR2_X1 U415 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U416 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U417 ( .A(KEYINPUT32), .B(KEYINPUT77), .Z(n364) );
  XOR2_X1 U418 ( .A(G176GAT), .B(G64GAT), .Z(n433) );
  XNOR2_X1 U419 ( .A(n362), .B(n433), .ZN(n363) );
  XNOR2_X1 U420 ( .A(n364), .B(n363), .ZN(n370) );
  XOR2_X1 U421 ( .A(KEYINPUT33), .B(KEYINPUT76), .Z(n366) );
  XNOR2_X1 U422 ( .A(KEYINPUT72), .B(KEYINPUT31), .ZN(n365) );
  XOR2_X1 U423 ( .A(n366), .B(n365), .Z(n368) );
  NAND2_X1 U424 ( .A1(G230GAT), .A2(G233GAT), .ZN(n367) );
  INV_X1 U425 ( .A(KEYINPUT73), .ZN(n371) );
  XNOR2_X1 U426 ( .A(n372), .B(n371), .ZN(n378) );
  XOR2_X1 U427 ( .A(G92GAT), .B(G85GAT), .Z(n374) );
  XNOR2_X1 U428 ( .A(G99GAT), .B(G106GAT), .ZN(n373) );
  XNOR2_X1 U429 ( .A(n374), .B(n373), .ZN(n383) );
  XNOR2_X1 U430 ( .A(n383), .B(KEYINPUT74), .ZN(n376) );
  XNOR2_X1 U431 ( .A(G57GAT), .B(KEYINPUT71), .ZN(n379) );
  XOR2_X1 U432 ( .A(n379), .B(KEYINPUT13), .Z(n399) );
  XNOR2_X1 U433 ( .A(n380), .B(n399), .ZN(n486) );
  XOR2_X1 U434 ( .A(KEYINPUT45), .B(KEYINPUT114), .Z(n416) );
  XOR2_X1 U435 ( .A(KEYINPUT65), .B(KEYINPUT9), .Z(n382) );
  XNOR2_X1 U436 ( .A(KEYINPUT10), .B(KEYINPUT80), .ZN(n381) );
  XNOR2_X1 U437 ( .A(n382), .B(n381), .ZN(n387) );
  XOR2_X1 U438 ( .A(n383), .B(G134GAT), .Z(n385) );
  NAND2_X1 U439 ( .A1(G232GAT), .A2(G233GAT), .ZN(n384) );
  XNOR2_X1 U440 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U441 ( .A(n387), .B(n386), .ZN(n392) );
  XOR2_X1 U442 ( .A(KEYINPUT11), .B(KEYINPUT81), .Z(n390) );
  XOR2_X1 U443 ( .A(G36GAT), .B(G190GAT), .Z(n435) );
  XNOR2_X1 U444 ( .A(n388), .B(n435), .ZN(n389) );
  XNOR2_X1 U445 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U446 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U447 ( .A(n394), .B(n393), .ZN(n564) );
  XNOR2_X1 U448 ( .A(KEYINPUT82), .B(n564), .ZN(n572) );
  XNOR2_X1 U449 ( .A(KEYINPUT36), .B(KEYINPUT103), .ZN(n395) );
  XNOR2_X1 U450 ( .A(n572), .B(n395), .ZN(n580) );
  XOR2_X1 U451 ( .A(KEYINPUT85), .B(KEYINPUT84), .Z(n401) );
  XOR2_X1 U452 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n397) );
  XNOR2_X1 U453 ( .A(KEYINPUT86), .B(KEYINPUT15), .ZN(n396) );
  XNOR2_X1 U454 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U455 ( .A(n399), .B(n398), .Z(n400) );
  XNOR2_X1 U456 ( .A(n401), .B(n400), .ZN(n414) );
  XOR2_X1 U457 ( .A(n403), .B(n402), .Z(n405) );
  NAND2_X1 U458 ( .A1(G231GAT), .A2(G233GAT), .ZN(n404) );
  XNOR2_X1 U459 ( .A(n405), .B(n404), .ZN(n412) );
  XOR2_X1 U460 ( .A(KEYINPUT83), .B(G64GAT), .Z(n407) );
  XNOR2_X1 U461 ( .A(G211GAT), .B(G78GAT), .ZN(n406) );
  XNOR2_X1 U462 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U463 ( .A(G8GAT), .B(G183GAT), .Z(n432) );
  XOR2_X1 U464 ( .A(n408), .B(n432), .Z(n410) );
  XNOR2_X1 U465 ( .A(G127GAT), .B(G71GAT), .ZN(n409) );
  XNOR2_X1 U466 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U467 ( .A(n412), .B(n411), .Z(n413) );
  XNOR2_X1 U468 ( .A(n414), .B(n413), .ZN(n577) );
  INV_X1 U469 ( .A(n577), .ZN(n500) );
  NOR2_X1 U470 ( .A1(n580), .A2(n500), .ZN(n415) );
  XOR2_X1 U471 ( .A(n416), .B(n415), .Z(n417) );
  NAND2_X1 U472 ( .A1(n486), .A2(n417), .ZN(n418) );
  NOR2_X1 U473 ( .A1(n567), .A2(n418), .ZN(n427) );
  XNOR2_X1 U474 ( .A(n486), .B(KEYINPUT41), .ZN(n456) );
  NAND2_X1 U475 ( .A1(n456), .A2(n567), .ZN(n420) );
  XNOR2_X1 U476 ( .A(KEYINPUT46), .B(KEYINPUT112), .ZN(n419) );
  XNOR2_X1 U477 ( .A(n420), .B(n419), .ZN(n421) );
  AND2_X1 U478 ( .A1(n421), .A2(n500), .ZN(n422) );
  XNOR2_X1 U479 ( .A(n422), .B(KEYINPUT113), .ZN(n423) );
  NOR2_X1 U480 ( .A1(n423), .A2(n564), .ZN(n425) );
  XNOR2_X1 U481 ( .A(n425), .B(n424), .ZN(n426) );
  NOR2_X1 U482 ( .A1(n427), .A2(n426), .ZN(n429) );
  INV_X1 U483 ( .A(KEYINPUT48), .ZN(n428) );
  XNOR2_X1 U484 ( .A(n429), .B(n428), .ZN(n537) );
  XOR2_X1 U485 ( .A(KEYINPUT95), .B(G92GAT), .Z(n431) );
  XNOR2_X1 U486 ( .A(G204GAT), .B(G218GAT), .ZN(n430) );
  XNOR2_X1 U487 ( .A(n431), .B(n430), .ZN(n445) );
  XNOR2_X1 U488 ( .A(n433), .B(n432), .ZN(n443) );
  XOR2_X1 U489 ( .A(n435), .B(n434), .Z(n437) );
  NAND2_X1 U490 ( .A1(G226GAT), .A2(G233GAT), .ZN(n436) );
  XNOR2_X1 U491 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U492 ( .A(n438), .B(KEYINPUT96), .Z(n441) );
  XNOR2_X1 U493 ( .A(n439), .B(KEYINPUT97), .ZN(n440) );
  XNOR2_X1 U494 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U495 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U496 ( .A(n445), .B(n444), .Z(n529) );
  AND2_X1 U497 ( .A1(n537), .A2(n529), .ZN(n446) );
  XOR2_X1 U498 ( .A(n446), .B(KEYINPUT54), .Z(n447) );
  NAND2_X1 U499 ( .A1(n471), .A2(n457), .ZN(n449) );
  INV_X1 U500 ( .A(KEYINPUT124), .ZN(n448) );
  NAND2_X1 U501 ( .A1(n567), .A2(n578), .ZN(n451) );
  XOR2_X1 U502 ( .A(KEYINPUT126), .B(KEYINPUT60), .Z(n450) );
  XNOR2_X1 U503 ( .A(n451), .B(n450), .ZN(n455) );
  XNOR2_X1 U504 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n453) );
  INV_X1 U505 ( .A(KEYINPUT125), .ZN(n452) );
  XOR2_X1 U506 ( .A(n456), .B(KEYINPUT107), .Z(n543) );
  AND2_X1 U507 ( .A1(n476), .A2(n457), .ZN(n458) );
  XNOR2_X1 U508 ( .A(KEYINPUT55), .B(n458), .ZN(n460) );
  NOR2_X2 U509 ( .A1(n460), .A2(n459), .ZN(n573) );
  NAND2_X1 U510 ( .A1(n543), .A2(n573), .ZN(n463) );
  XOR2_X1 U511 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n461) );
  XNOR2_X1 U512 ( .A(n461), .B(G176GAT), .ZN(n462) );
  XNOR2_X1 U513 ( .A(n463), .B(n462), .ZN(G1349GAT) );
  INV_X1 U514 ( .A(G204GAT), .ZN(n467) );
  XOR2_X1 U515 ( .A(KEYINPUT127), .B(KEYINPUT61), .Z(n465) );
  INV_X1 U516 ( .A(n578), .ZN(n581) );
  OR2_X1 U517 ( .A1(n581), .A2(n486), .ZN(n464) );
  XNOR2_X1 U518 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U519 ( .A(n467), .B(n466), .ZN(G1353GAT) );
  NAND2_X1 U520 ( .A1(n540), .A2(n529), .ZN(n468) );
  NAND2_X1 U521 ( .A1(n476), .A2(n468), .ZN(n469) );
  XOR2_X1 U522 ( .A(KEYINPUT25), .B(n469), .Z(n473) );
  XOR2_X1 U523 ( .A(KEYINPUT27), .B(KEYINPUT98), .Z(n470) );
  XNOR2_X1 U524 ( .A(n529), .B(n470), .ZN(n478) );
  INV_X1 U525 ( .A(n478), .ZN(n472) );
  NAND2_X1 U526 ( .A1(n472), .A2(n471), .ZN(n554) );
  NAND2_X1 U527 ( .A1(n473), .A2(n554), .ZN(n474) );
  XNOR2_X1 U528 ( .A(KEYINPUT99), .B(n474), .ZN(n475) );
  NOR2_X1 U529 ( .A1(n538), .A2(n475), .ZN(n481) );
  XNOR2_X1 U530 ( .A(n476), .B(KEYINPUT66), .ZN(n477) );
  XOR2_X1 U531 ( .A(n477), .B(KEYINPUT28), .Z(n534) );
  NOR2_X1 U532 ( .A1(n478), .A2(n534), .ZN(n539) );
  NAND2_X1 U533 ( .A1(n538), .A2(n539), .ZN(n479) );
  NOR2_X1 U534 ( .A1(n540), .A2(n479), .ZN(n480) );
  NOR2_X1 U535 ( .A1(n481), .A2(n480), .ZN(n498) );
  XNOR2_X1 U536 ( .A(KEYINPUT88), .B(KEYINPUT87), .ZN(n483) );
  NOR2_X1 U537 ( .A1(n572), .A2(n500), .ZN(n482) );
  XNOR2_X1 U538 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U539 ( .A(n484), .B(KEYINPUT16), .ZN(n485) );
  NOR2_X1 U540 ( .A1(n498), .A2(n485), .ZN(n515) );
  NAND2_X1 U541 ( .A1(n486), .A2(n567), .ZN(n487) );
  XOR2_X1 U542 ( .A(KEYINPUT78), .B(n487), .Z(n502) );
  AND2_X1 U543 ( .A1(n515), .A2(n502), .ZN(n495) );
  NAND2_X1 U544 ( .A1(n495), .A2(n538), .ZN(n491) );
  XOR2_X1 U545 ( .A(KEYINPUT101), .B(KEYINPUT100), .Z(n489) );
  XNOR2_X1 U546 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n488) );
  XNOR2_X1 U547 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U548 ( .A(n491), .B(n490), .ZN(G1324GAT) );
  NAND2_X1 U549 ( .A1(n495), .A2(n529), .ZN(n492) );
  XNOR2_X1 U550 ( .A(n492), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U551 ( .A(G15GAT), .B(KEYINPUT35), .Z(n494) );
  NAND2_X1 U552 ( .A1(n495), .A2(n540), .ZN(n493) );
  XNOR2_X1 U553 ( .A(n494), .B(n493), .ZN(G1326GAT) );
  NAND2_X1 U554 ( .A1(n534), .A2(n495), .ZN(n496) );
  XNOR2_X1 U555 ( .A(n496), .B(KEYINPUT102), .ZN(n497) );
  XNOR2_X1 U556 ( .A(G22GAT), .B(n497), .ZN(G1327GAT) );
  XOR2_X1 U557 ( .A(G29GAT), .B(KEYINPUT39), .Z(n505) );
  NOR2_X1 U558 ( .A1(n580), .A2(n498), .ZN(n499) );
  NAND2_X1 U559 ( .A1(n500), .A2(n499), .ZN(n501) );
  XNOR2_X1 U560 ( .A(KEYINPUT37), .B(n501), .ZN(n527) );
  NAND2_X1 U561 ( .A1(n527), .A2(n502), .ZN(n503) );
  XOR2_X1 U562 ( .A(KEYINPUT38), .B(n503), .Z(n511) );
  NAND2_X1 U563 ( .A1(n538), .A2(n511), .ZN(n504) );
  XNOR2_X1 U564 ( .A(n505), .B(n504), .ZN(G1328GAT) );
  XOR2_X1 U565 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n507) );
  NAND2_X1 U566 ( .A1(n529), .A2(n511), .ZN(n506) );
  XNOR2_X1 U567 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U568 ( .A(G36GAT), .B(n508), .ZN(G1329GAT) );
  NAND2_X1 U569 ( .A1(n511), .A2(n540), .ZN(n509) );
  XNOR2_X1 U570 ( .A(n509), .B(KEYINPUT40), .ZN(n510) );
  XNOR2_X1 U571 ( .A(G43GAT), .B(n510), .ZN(G1330GAT) );
  NAND2_X1 U572 ( .A1(n511), .A2(n534), .ZN(n512) );
  XNOR2_X1 U573 ( .A(n512), .B(KEYINPUT106), .ZN(n513) );
  XNOR2_X1 U574 ( .A(G50GAT), .B(n513), .ZN(G1331GAT) );
  XOR2_X1 U575 ( .A(KEYINPUT42), .B(KEYINPUT109), .Z(n518) );
  INV_X1 U576 ( .A(n543), .ZN(n514) );
  NOR2_X1 U577 ( .A1(n567), .A2(n514), .ZN(n526) );
  NAND2_X1 U578 ( .A1(n515), .A2(n526), .ZN(n516) );
  XOR2_X1 U579 ( .A(KEYINPUT108), .B(n516), .Z(n522) );
  NAND2_X1 U580 ( .A1(n538), .A2(n522), .ZN(n517) );
  XNOR2_X1 U581 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U582 ( .A(G57GAT), .B(n519), .ZN(G1332GAT) );
  NAND2_X1 U583 ( .A1(n522), .A2(n529), .ZN(n520) );
  XNOR2_X1 U584 ( .A(n520), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U585 ( .A1(n522), .A2(n540), .ZN(n521) );
  XNOR2_X1 U586 ( .A(n521), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U587 ( .A(KEYINPUT110), .B(KEYINPUT43), .Z(n524) );
  NAND2_X1 U588 ( .A1(n522), .A2(n534), .ZN(n523) );
  XNOR2_X1 U589 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U590 ( .A(G78GAT), .B(n525), .ZN(G1335GAT) );
  AND2_X1 U591 ( .A1(n527), .A2(n526), .ZN(n533) );
  NAND2_X1 U592 ( .A1(n538), .A2(n533), .ZN(n528) );
  XNOR2_X1 U593 ( .A(G85GAT), .B(n528), .ZN(G1336GAT) );
  XOR2_X1 U594 ( .A(G92GAT), .B(KEYINPUT111), .Z(n531) );
  NAND2_X1 U595 ( .A1(n533), .A2(n529), .ZN(n530) );
  XNOR2_X1 U596 ( .A(n531), .B(n530), .ZN(G1337GAT) );
  NAND2_X1 U597 ( .A1(n533), .A2(n540), .ZN(n532) );
  XNOR2_X1 U598 ( .A(n532), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U599 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U600 ( .A(n535), .B(KEYINPUT44), .ZN(n536) );
  XNOR2_X1 U601 ( .A(G106GAT), .B(n536), .ZN(G1339GAT) );
  NAND2_X1 U602 ( .A1(n538), .A2(n537), .ZN(n555) );
  NAND2_X1 U603 ( .A1(n540), .A2(n539), .ZN(n541) );
  NOR2_X1 U604 ( .A1(n555), .A2(n541), .ZN(n550) );
  NAND2_X1 U605 ( .A1(n567), .A2(n550), .ZN(n542) );
  XNOR2_X1 U606 ( .A(G113GAT), .B(n542), .ZN(G1340GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT49), .B(KEYINPUT116), .Z(n545) );
  NAND2_X1 U608 ( .A1(n550), .A2(n543), .ZN(n544) );
  XNOR2_X1 U609 ( .A(n545), .B(n544), .ZN(n547) );
  XOR2_X1 U610 ( .A(G120GAT), .B(KEYINPUT115), .Z(n546) );
  XNOR2_X1 U611 ( .A(n547), .B(n546), .ZN(G1341GAT) );
  NAND2_X1 U612 ( .A1(n577), .A2(n550), .ZN(n548) );
  XNOR2_X1 U613 ( .A(n548), .B(KEYINPUT50), .ZN(n549) );
  XNOR2_X1 U614 ( .A(G127GAT), .B(n549), .ZN(G1342GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n552) );
  NAND2_X1 U616 ( .A1(n550), .A2(n572), .ZN(n551) );
  XNOR2_X1 U617 ( .A(n552), .B(n551), .ZN(n553) );
  XOR2_X1 U618 ( .A(G134GAT), .B(n553), .Z(G1343GAT) );
  XOR2_X1 U619 ( .A(G141GAT), .B(KEYINPUT119), .Z(n558) );
  NOR2_X1 U620 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U621 ( .A(n556), .B(KEYINPUT118), .ZN(n565) );
  NAND2_X1 U622 ( .A1(n567), .A2(n565), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n558), .B(n557), .ZN(G1344GAT) );
  XOR2_X1 U624 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n560) );
  NAND2_X1 U625 ( .A1(n456), .A2(n565), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U627 ( .A(G148GAT), .B(n561), .ZN(G1345GAT) );
  NAND2_X1 U628 ( .A1(n565), .A2(n577), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n562), .B(KEYINPUT120), .ZN(n563) );
  XNOR2_X1 U630 ( .A(G155GAT), .B(n563), .ZN(G1346GAT) );
  NAND2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n566), .B(G162GAT), .ZN(G1347GAT) );
  XOR2_X1 U633 ( .A(G169GAT), .B(KEYINPUT121), .Z(n569) );
  NAND2_X1 U634 ( .A1(n573), .A2(n567), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(G1348GAT) );
  NAND2_X1 U636 ( .A1(n577), .A2(n573), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n570), .B(KEYINPUT122), .ZN(n571) );
  XNOR2_X1 U638 ( .A(G183GAT), .B(n571), .ZN(G1350GAT) );
  XOR2_X1 U639 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n575) );
  NAND2_X1 U640 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U642 ( .A(G190GAT), .B(n576), .ZN(G1351GAT) );
  NAND2_X1 U643 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n579), .B(G211GAT), .ZN(G1354GAT) );
  INV_X1 U645 ( .A(KEYINPUT62), .ZN(n583) );
  NOR2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(n584), .ZN(G1355GAT) );
endmodule

