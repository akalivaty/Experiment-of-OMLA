//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 0 0 0 0 0 1 0 0 0 1 0 1 0 0 1 1 0 0 1 1 1 0 0 1 1 1 1 0 0 0 0 0 0 0 0 1 0 1 1 0 0 1 0 0 0 1 0 0 0 0 0 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:56 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n444, new_n448, new_n449, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n565, new_n567, new_n568, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n623, new_n624, new_n626,
    new_n627, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1163, new_n1164, new_n1165;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  XOR2_X1   g016(.A(KEYINPUT65), .B(G108), .Z(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT66), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT67), .Z(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NOR4_X1   g029(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(new_n455), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(G567), .ZN(new_n459));
  OR2_X1    g034(.A1(new_n459), .A2(KEYINPUT68), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(KEYINPUT68), .ZN(new_n461));
  INV_X1    g036(.A(G2106), .ZN(new_n462));
  OAI211_X1 g037(.A(new_n460), .B(new_n461), .C1(new_n462), .C2(new_n454), .ZN(new_n463));
  XOR2_X1   g038(.A(new_n463), .B(KEYINPUT69), .Z(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(G319));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G125), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n466), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(G101), .A2(G2104), .ZN(new_n475));
  INV_X1    g050(.A(G137), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n475), .B1(new_n471), .B2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n474), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G160));
  NOR2_X1   g056(.A1(new_n471), .A2(G2105), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  NOR2_X1   g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(new_n478), .B2(G112), .ZN(new_n485));
  INV_X1    g060(.A(new_n471), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n486), .A2(KEYINPUT70), .A3(G2105), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT70), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n488), .B1(new_n471), .B2(new_n478), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(G124), .ZN(new_n491));
  OAI221_X1 g066(.A(new_n483), .B1(new_n484), .B2(new_n485), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  NAND4_X1  g068(.A1(new_n468), .A2(new_n470), .A3(G138), .A4(new_n478), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  OR2_X1    g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n494), .A2(new_n495), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OAI21_X1  g073(.A(KEYINPUT71), .B1(new_n478), .B2(G114), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT71), .ZN(new_n500));
  INV_X1    g075(.A(G114), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n500), .A2(new_n501), .A3(G2105), .ZN(new_n502));
  OR2_X1    g077(.A1(G102), .A2(G2105), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n499), .A2(new_n502), .A3(G2104), .A4(new_n503), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n468), .A2(new_n470), .A3(G126), .A4(G2105), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n498), .A2(new_n506), .ZN(G164));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(KEYINPUT5), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT5), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n513), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AND2_X1   g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  NOR2_X1   g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  OR2_X1    g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G543), .ZN(new_n520));
  INV_X1    g095(.A(G50), .ZN(new_n521));
  INV_X1    g096(.A(G88), .ZN(new_n522));
  OAI211_X1 g097(.A(new_n509), .B(new_n511), .C1(new_n517), .C2(new_n518), .ZN(new_n523));
  OAI22_X1  g098(.A1(new_n520), .A2(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n516), .A2(new_n524), .ZN(G166));
  NOR2_X1   g100(.A1(new_n510), .A2(G543), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n508), .A2(KEYINPUT5), .ZN(new_n527));
  OAI21_X1  g102(.A(KEYINPUT72), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT72), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n509), .A2(new_n511), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n531), .A2(G63), .A3(G651), .ZN(new_n532));
  INV_X1    g107(.A(new_n532), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n513), .A2(new_n519), .A3(G89), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n519), .A2(G51), .A3(G543), .ZN(new_n535));
  NAND3_X1  g110(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT7), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n534), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n533), .A2(new_n538), .ZN(G168));
  AOI22_X1  g114(.A1(new_n531), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n540), .A2(new_n515), .ZN(new_n541));
  INV_X1    g116(.A(G52), .ZN(new_n542));
  XNOR2_X1  g117(.A(KEYINPUT73), .B(G90), .ZN(new_n543));
  OAI22_X1  g118(.A1(new_n520), .A2(new_n542), .B1(new_n523), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n541), .A2(new_n544), .ZN(G171));
  AND3_X1   g120(.A1(new_n509), .A2(new_n511), .A3(new_n529), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n529), .B1(new_n509), .B2(new_n511), .ZN(new_n547));
  OAI21_X1  g122(.A(G56), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(G68), .A2(G543), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n515), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  OAI211_X1 g125(.A(G43), .B(G543), .C1(new_n517), .C2(new_n518), .ZN(new_n551));
  INV_X1    g126(.A(G81), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n551), .B1(new_n523), .B2(new_n552), .ZN(new_n553));
  NOR3_X1   g128(.A1(new_n550), .A2(KEYINPUT74), .A3(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT74), .ZN(new_n555));
  INV_X1    g130(.A(G56), .ZN(new_n556));
  AOI21_X1  g131(.A(new_n556), .B1(new_n528), .B2(new_n530), .ZN(new_n557));
  INV_X1    g132(.A(new_n549), .ZN(new_n558));
  OAI21_X1  g133(.A(G651), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n553), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n555), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n554), .A2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(G153));
  AND3_X1   g139(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G36), .ZN(G176));
  NAND2_X1  g141(.A1(G1), .A2(G3), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT8), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n565), .A2(new_n568), .ZN(G188));
  INV_X1    g144(.A(new_n520), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n570), .A2(KEYINPUT9), .A3(G53), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT9), .ZN(new_n572));
  INV_X1    g147(.A(G53), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n520), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(G78), .A2(G543), .ZN(new_n576));
  XOR2_X1   g151(.A(KEYINPUT75), .B(G65), .Z(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n577), .B2(new_n512), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(G651), .ZN(new_n579));
  INV_X1    g154(.A(G91), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n580), .B2(new_n523), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n575), .A2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(G299));
  INV_X1    g158(.A(G171), .ZN(G301));
  INV_X1    g159(.A(G168), .ZN(G286));
  INV_X1    g160(.A(G166), .ZN(G303));
  INV_X1    g161(.A(G49), .ZN(new_n587));
  INV_X1    g162(.A(G87), .ZN(new_n588));
  OAI22_X1  g163(.A1(new_n520), .A2(new_n587), .B1(new_n588), .B2(new_n523), .ZN(new_n589));
  OR2_X1    g164(.A1(new_n531), .A2(G74), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n589), .B1(new_n590), .B2(G651), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(G288));
  INV_X1    g167(.A(G48), .ZN(new_n593));
  INV_X1    g168(.A(G86), .ZN(new_n594));
  OAI22_X1  g169(.A1(new_n520), .A2(new_n593), .B1(new_n594), .B2(new_n523), .ZN(new_n595));
  NAND2_X1  g170(.A1(G73), .A2(G543), .ZN(new_n596));
  INV_X1    g171(.A(G61), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n512), .B2(new_n597), .ZN(new_n598));
  AND2_X1   g173(.A1(new_n598), .A2(G651), .ZN(new_n599));
  OR2_X1    g174(.A1(new_n595), .A2(new_n599), .ZN(G305));
  AOI22_X1  g175(.A1(new_n531), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n601), .A2(new_n515), .ZN(new_n602));
  XNOR2_X1  g177(.A(KEYINPUT76), .B(G47), .ZN(new_n603));
  INV_X1    g178(.A(G85), .ZN(new_n604));
  OAI22_X1  g179(.A1(new_n520), .A2(new_n603), .B1(new_n604), .B2(new_n523), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(G290));
  NAND2_X1  g182(.A1(G79), .A2(G543), .ZN(new_n608));
  INV_X1    g183(.A(G66), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n512), .B2(new_n609), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n570), .A2(G54), .B1(new_n610), .B2(G651), .ZN(new_n611));
  INV_X1    g186(.A(G92), .ZN(new_n612));
  OAI21_X1  g187(.A(KEYINPUT10), .B1(new_n523), .B2(new_n612), .ZN(new_n613));
  OR3_X1    g188(.A1(new_n523), .A2(KEYINPUT10), .A3(new_n612), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n611), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(G868), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(G171), .B2(new_n616), .ZN(G284));
  OAI21_X1  g193(.A(new_n617), .B1(G171), .B2(new_n616), .ZN(G321));
  NAND2_X1  g194(.A1(G286), .A2(G868), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(G868), .B2(new_n582), .ZN(G297));
  XOR2_X1   g196(.A(G297), .B(KEYINPUT77), .Z(G280));
  INV_X1    g197(.A(new_n615), .ZN(new_n623));
  INV_X1    g198(.A(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n623), .B1(new_n624), .B2(G860), .ZN(G148));
  NAND2_X1  g200(.A1(new_n562), .A2(new_n616), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n615), .A2(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n616), .B2(new_n627), .ZN(G323));
  XNOR2_X1  g203(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g204(.A(G2100), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n630), .A2(KEYINPUT79), .ZN(new_n631));
  INV_X1    g206(.A(new_n490), .ZN(new_n632));
  AOI22_X1  g207(.A1(new_n632), .A2(G123), .B1(G135), .B2(new_n482), .ZN(new_n633));
  OR2_X1    g208(.A1(G99), .A2(G2105), .ZN(new_n634));
  OAI211_X1 g209(.A(new_n634), .B(G2104), .C1(G111), .C2(new_n478), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n631), .B1(new_n636), .B2(G2096), .ZN(new_n637));
  XOR2_X1   g212(.A(KEYINPUT78), .B(KEYINPUT12), .Z(new_n638));
  NOR3_X1   g213(.A1(new_n469), .A2(new_n467), .A3(G2105), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n630), .A2(KEYINPUT79), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(KEYINPUT13), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n640), .B(new_n642), .ZN(new_n643));
  OAI211_X1 g218(.A(new_n637), .B(new_n643), .C1(G2096), .C2(new_n636), .ZN(G156));
  XNOR2_X1  g219(.A(KEYINPUT15), .B(G2430), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2435), .ZN(new_n646));
  XOR2_X1   g221(.A(G2427), .B(G2438), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n648), .A2(KEYINPUT14), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2451), .B(G2454), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT80), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT16), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n649), .B(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G1341), .B(G1348), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2443), .B(G2446), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n655), .A2(new_n656), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n657), .A2(G14), .A3(new_n658), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(G401));
  XNOR2_X1  g235(.A(G2072), .B(G2078), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2067), .B(G2678), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G2084), .B(G2090), .Z(new_n664));
  NOR2_X1   g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n661), .B(KEYINPUT17), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(new_n662), .ZN(new_n668));
  OAI21_X1  g243(.A(new_n665), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT81), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n664), .A2(new_n661), .A3(new_n662), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(KEYINPUT18), .Z(new_n672));
  NAND3_X1  g247(.A1(new_n667), .A2(new_n664), .A3(new_n668), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n670), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n674), .B(G2096), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(new_n630), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(G227));
  XNOR2_X1  g252(.A(G1971), .B(G1976), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT19), .ZN(new_n679));
  XOR2_X1   g254(.A(G1956), .B(G2474), .Z(new_n680));
  XOR2_X1   g255(.A(G1961), .B(G1966), .Z(new_n681));
  NAND2_X1  g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT82), .B(KEYINPUT20), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n680), .A2(new_n681), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n687), .A2(new_n679), .A3(new_n682), .ZN(new_n688));
  OAI211_X1 g263(.A(new_n685), .B(new_n688), .C1(new_n679), .C2(new_n687), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT83), .B(G1981), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n689), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1991), .B(G1996), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(G1986), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n693), .B(new_n695), .ZN(G229));
  INV_X1    g271(.A(G16), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(G23), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n698), .B1(new_n591), .B2(new_n697), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT33), .B(G1976), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT87), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n699), .B(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n697), .A2(G22), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(G166), .B2(new_n697), .ZN(new_n704));
  XOR2_X1   g279(.A(KEYINPUT88), .B(G1971), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n697), .A2(G6), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n595), .A2(new_n599), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n707), .B1(new_n708), .B2(new_n697), .ZN(new_n709));
  XOR2_X1   g284(.A(KEYINPUT32), .B(G1981), .Z(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n702), .A2(new_n706), .A3(new_n711), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(KEYINPUT34), .Z(new_n713));
  NOR2_X1   g288(.A1(G16), .A2(G24), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n606), .B(KEYINPUT86), .Z(new_n715));
  AOI21_X1  g290(.A(new_n714), .B1(new_n715), .B2(G16), .ZN(new_n716));
  INV_X1    g291(.A(G1986), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT84), .B(G29), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n719), .A2(G25), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n632), .A2(G119), .ZN(new_n721));
  NOR2_X1   g296(.A1(G95), .A2(G2105), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(KEYINPUT85), .Z(new_n723));
  INV_X1    g298(.A(G107), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n467), .B1(new_n724), .B2(G2105), .ZN(new_n725));
  AOI22_X1  g300(.A1(new_n723), .A2(new_n725), .B1(new_n482), .B2(G131), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n721), .A2(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(new_n727), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n720), .B1(new_n728), .B2(new_n719), .ZN(new_n729));
  XOR2_X1   g304(.A(KEYINPUT35), .B(G1991), .Z(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n713), .A2(new_n718), .A3(new_n731), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT36), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n563), .A2(new_n697), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(new_n697), .B2(G19), .ZN(new_n735));
  XNOR2_X1  g310(.A(KEYINPUT91), .B(G1341), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n632), .A2(G129), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n478), .A2(G105), .A3(G2104), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n482), .A2(G141), .ZN(new_n740));
  NAND3_X1  g315(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT26), .Z(new_n742));
  NAND4_X1  g317(.A1(new_n738), .A2(new_n739), .A3(new_n740), .A4(new_n742), .ZN(new_n743));
  MUX2_X1   g318(.A(G32), .B(new_n743), .S(G29), .Z(new_n744));
  XOR2_X1   g319(.A(KEYINPUT27), .B(G1996), .Z(new_n745));
  NOR2_X1   g320(.A1(G5), .A2(G16), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(G171), .B2(G16), .ZN(new_n747));
  OAI22_X1  g322(.A1(new_n744), .A2(new_n745), .B1(G1961), .B2(new_n747), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n737), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n697), .A2(G4), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(new_n623), .B2(new_n697), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT90), .ZN(new_n752));
  XNOR2_X1  g327(.A(KEYINPUT89), .B(G1348), .ZN(new_n753));
  AOI22_X1  g328(.A1(new_n752), .A2(new_n753), .B1(G1961), .B2(new_n747), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n735), .A2(new_n736), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n749), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(new_n719), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n757), .A2(G35), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G162), .B2(new_n757), .ZN(new_n759));
  XOR2_X1   g334(.A(KEYINPUT29), .B(G2090), .Z(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n482), .A2(G139), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n478), .A2(G103), .A3(G2104), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT25), .Z(new_n764));
  AOI22_X1  g339(.A1(new_n486), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n765));
  OAI211_X1 g340(.A(new_n762), .B(new_n764), .C1(new_n765), .C2(new_n478), .ZN(new_n766));
  MUX2_X1   g341(.A(G33), .B(new_n766), .S(G29), .Z(new_n767));
  NOR2_X1   g342(.A1(new_n767), .A2(G2072), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n719), .A2(G27), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(G164), .B2(new_n719), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n768), .B1(G2078), .B2(new_n770), .ZN(new_n771));
  OAI211_X1 g346(.A(new_n761), .B(new_n771), .C1(G2078), .C2(new_n770), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n697), .A2(KEYINPUT23), .A3(G20), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT23), .ZN(new_n774));
  INV_X1    g349(.A(G20), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n774), .B1(new_n775), .B2(G16), .ZN(new_n776));
  OAI211_X1 g351(.A(new_n773), .B(new_n776), .C1(new_n582), .C2(new_n697), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(G1956), .ZN(new_n778));
  INV_X1    g353(.A(G29), .ZN(new_n779));
  XNOR2_X1  g354(.A(KEYINPUT30), .B(G28), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n778), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT24), .B(G34), .ZN(new_n782));
  AOI22_X1  g357(.A1(G160), .A2(G29), .B1(new_n757), .B2(new_n782), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(G2084), .Z(new_n784));
  NAND3_X1  g359(.A1(new_n633), .A2(new_n635), .A3(new_n719), .ZN(new_n785));
  AOI22_X1  g360(.A1(new_n744), .A2(new_n745), .B1(G2072), .B2(new_n767), .ZN(new_n786));
  NAND4_X1  g361(.A1(new_n781), .A2(new_n784), .A3(new_n785), .A4(new_n786), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n752), .A2(new_n753), .ZN(new_n788));
  NOR4_X1   g363(.A1(new_n756), .A2(new_n772), .A3(new_n787), .A4(new_n788), .ZN(new_n789));
  AND2_X1   g364(.A1(new_n733), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n482), .A2(G140), .ZN(new_n791));
  NOR2_X1   g366(.A1(G104), .A2(G2105), .ZN(new_n792));
  OAI21_X1  g367(.A(G2104), .B1(new_n478), .B2(G116), .ZN(new_n793));
  INV_X1    g368(.A(G128), .ZN(new_n794));
  OAI221_X1 g369(.A(new_n791), .B1(new_n792), .B2(new_n793), .C1(new_n490), .C2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n795), .A2(G29), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT92), .Z(new_n797));
  NAND2_X1  g372(.A1(new_n757), .A2(G26), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT28), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  XNOR2_X1  g375(.A(KEYINPUT93), .B(G2067), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n697), .A2(G21), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(G168), .B2(new_n697), .ZN(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT94), .B(G1966), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  XNOR2_X1  g383(.A(KEYINPUT31), .B(G11), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n790), .A2(new_n803), .A3(new_n808), .A4(new_n809), .ZN(G150));
  INV_X1    g385(.A(G150), .ZN(G311));
  OAI211_X1 g386(.A(G55), .B(G543), .C1(new_n517), .C2(new_n518), .ZN(new_n812));
  INV_X1    g387(.A(G93), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n812), .B1(new_n523), .B2(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  AOI22_X1  g390(.A1(new_n531), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n815), .B1(new_n816), .B2(new_n515), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n817), .A2(G860), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT37), .Z(new_n819));
  NAND2_X1  g394(.A1(new_n548), .A2(new_n549), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n553), .B1(new_n820), .B2(G651), .ZN(new_n821));
  OAI21_X1  g396(.A(KEYINPUT95), .B1(new_n817), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n559), .A2(new_n560), .ZN(new_n823));
  OAI21_X1  g398(.A(G67), .B1(new_n546), .B2(new_n547), .ZN(new_n824));
  NAND2_X1  g399(.A1(G80), .A2(G543), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n814), .B1(new_n826), .B2(G651), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT95), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n823), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n822), .A2(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT96), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n817), .B1(new_n554), .B2(new_n561), .ZN(new_n832));
  AND3_X1   g407(.A1(new_n830), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n831), .B1(new_n830), .B2(new_n832), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n615), .A2(new_n624), .ZN(new_n836));
  XOR2_X1   g411(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n837));
  XOR2_X1   g412(.A(new_n836), .B(new_n837), .Z(new_n838));
  XNOR2_X1  g413(.A(new_n835), .B(new_n838), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n819), .B1(new_n839), .B2(G860), .ZN(G145));
  NAND2_X1  g415(.A1(new_n506), .A2(KEYINPUT97), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT97), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n504), .A2(new_n842), .A3(new_n505), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  AND2_X1   g419(.A1(new_n496), .A2(new_n497), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n795), .B(new_n846), .ZN(new_n847));
  AOI22_X1  g422(.A1(new_n632), .A2(G130), .B1(G142), .B2(new_n482), .ZN(new_n848));
  NOR2_X1   g423(.A1(G106), .A2(G2105), .ZN(new_n849));
  OAI21_X1  g424(.A(G2104), .B1(new_n478), .B2(G118), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n848), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n847), .B(new_n851), .Z(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n743), .B(new_n727), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n766), .B(new_n640), .Z(new_n855));
  OR2_X1    g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n854), .A2(new_n855), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n853), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n852), .A2(new_n856), .A3(new_n857), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT98), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n636), .B(G160), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(G162), .ZN(new_n864));
  AND3_X1   g439(.A1(new_n861), .A2(new_n862), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n862), .B1(new_n861), .B2(new_n864), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n861), .A2(new_n864), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n868), .A2(G37), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g446(.A1(new_n817), .A2(new_n616), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n835), .B(new_n627), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n582), .B(new_n615), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  OR3_X1    g450(.A1(new_n873), .A2(KEYINPUT99), .A3(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n874), .B(KEYINPUT41), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n873), .A2(new_n878), .ZN(new_n879));
  OAI21_X1  g454(.A(KEYINPUT99), .B1(new_n873), .B2(new_n875), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n876), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n606), .B(new_n591), .ZN(new_n882));
  XNOR2_X1  g457(.A(G166), .B(new_n708), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n882), .B(new_n883), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n884), .A2(KEYINPUT100), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(KEYINPUT42), .ZN(new_n886));
  XOR2_X1   g461(.A(new_n881), .B(new_n886), .Z(new_n887));
  OAI21_X1  g462(.A(new_n872), .B1(new_n887), .B2(new_n616), .ZN(G295));
  OAI21_X1  g463(.A(new_n872), .B1(new_n887), .B2(new_n616), .ZN(G331));
  INV_X1    g464(.A(KEYINPUT101), .ZN(new_n890));
  NAND2_X1  g465(.A1(G168), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g466(.A(KEYINPUT101), .B1(new_n533), .B2(new_n538), .ZN(new_n892));
  AOI21_X1  g467(.A(G171), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n891), .A2(G171), .A3(new_n892), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n896), .B1(new_n833), .B2(new_n834), .ZN(new_n897));
  NOR3_X1   g472(.A1(new_n817), .A2(new_n821), .A3(KEYINPUT95), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n828), .B1(new_n823), .B2(new_n827), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n832), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(KEYINPUT96), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n830), .A2(new_n831), .A3(new_n832), .ZN(new_n902));
  AND3_X1   g477(.A1(new_n891), .A2(G171), .A3(new_n892), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n903), .A2(new_n893), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n901), .A2(new_n902), .A3(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT102), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n897), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  OAI211_X1 g482(.A(KEYINPUT102), .B(new_n896), .C1(new_n833), .C2(new_n834), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n907), .A2(new_n908), .A3(new_n878), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n897), .A2(new_n905), .A3(new_n874), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n909), .A2(new_n884), .A3(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(G37), .ZN(new_n912));
  AND2_X1   g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT104), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT43), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n884), .B(KEYINPUT103), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n875), .B1(new_n907), .B2(new_n908), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n877), .B1(new_n897), .B2(new_n905), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n916), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n913), .A2(new_n914), .A3(new_n915), .A4(new_n919), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n919), .A2(new_n915), .A3(new_n912), .A4(new_n911), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(KEYINPUT104), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n911), .A2(new_n912), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT103), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n884), .B(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n925), .B1(new_n909), .B2(new_n910), .ZN(new_n926));
  OAI21_X1  g501(.A(KEYINPUT43), .B1(new_n923), .B2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n920), .A2(new_n922), .A3(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT44), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n923), .A2(new_n926), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n929), .B1(new_n931), .B2(new_n915), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT105), .ZN(new_n933));
  INV_X1    g508(.A(new_n919), .ZN(new_n934));
  OAI21_X1  g509(.A(KEYINPUT43), .B1(new_n934), .B2(new_n923), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n932), .A2(new_n933), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n933), .B1(new_n932), .B2(new_n935), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n930), .B1(new_n936), .B2(new_n937), .ZN(G397));
  INV_X1    g513(.A(KEYINPUT106), .ZN(new_n939));
  AOI21_X1  g514(.A(G1384), .B1(new_n844), .B2(new_n845), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT45), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  AND3_X1   g518(.A1(new_n474), .A2(new_n479), .A3(G40), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n939), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n941), .A2(KEYINPUT106), .A3(new_n942), .A4(new_n944), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n727), .B(new_n730), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n950), .B(KEYINPUT107), .ZN(new_n951));
  INV_X1    g526(.A(G2067), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n795), .B(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(G1996), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n743), .B(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n951), .A2(new_n953), .A3(new_n955), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n606), .B(new_n717), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n949), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT124), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n940), .A2(KEYINPUT45), .ZN(new_n960));
  INV_X1    g535(.A(G1384), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n961), .B1(new_n498), .B2(new_n506), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(new_n942), .ZN(new_n963));
  INV_X1    g538(.A(G2078), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n960), .A2(new_n963), .A3(new_n964), .A4(new_n944), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT53), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT50), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n846), .A2(new_n967), .A3(new_n961), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n962), .A2(KEYINPUT50), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n968), .A2(new_n969), .A3(new_n944), .ZN(new_n970));
  INV_X1    g545(.A(G1961), .ZN(new_n971));
  AOI22_X1  g546(.A1(new_n965), .A2(new_n966), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n966), .A2(G2078), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n943), .A2(new_n944), .A3(new_n960), .A4(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n972), .A2(G301), .A3(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT54), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  OAI211_X1 g552(.A(KEYINPUT45), .B(new_n961), .C1(new_n498), .C2(new_n506), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n943), .A2(new_n944), .A3(new_n978), .A4(new_n973), .ZN(new_n979));
  AOI21_X1  g554(.A(G301), .B1(new_n972), .B2(new_n979), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n977), .A2(new_n980), .ZN(new_n981));
  AND2_X1   g556(.A1(new_n972), .A2(G301), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n979), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n965), .A2(new_n966), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n970), .A2(new_n971), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n984), .A2(new_n985), .A3(new_n974), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT123), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n972), .A2(KEYINPUT123), .A3(new_n974), .ZN(new_n989));
  AND2_X1   g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n983), .B1(new_n990), .B2(G301), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n981), .B1(new_n991), .B2(KEYINPUT54), .ZN(new_n992));
  INV_X1    g567(.A(G8), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n944), .B1(new_n940), .B2(new_n967), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT112), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(G2090), .ZN(new_n997));
  OR2_X1    g572(.A1(new_n962), .A2(KEYINPUT50), .ZN(new_n998));
  OAI211_X1 g573(.A(KEYINPUT112), .B(new_n944), .C1(new_n940), .C2(new_n967), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n996), .A2(new_n997), .A3(new_n998), .A4(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n960), .A2(new_n963), .A3(new_n944), .ZN(new_n1001));
  INV_X1    g576(.A(G1971), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n993), .B1(new_n1000), .B2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g579(.A1(G166), .A2(new_n993), .ZN(new_n1005));
  XNOR2_X1  g580(.A(new_n1005), .B(KEYINPUT55), .ZN(new_n1006));
  OR2_X1    g581(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT108), .ZN(new_n1008));
  OR3_X1    g583(.A1(new_n970), .A2(new_n1008), .A3(G2090), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1008), .B1(new_n970), .B2(G2090), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1009), .A2(new_n1003), .A3(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1011), .A2(G8), .A3(new_n1006), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT110), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1013), .B1(G305), .B2(G1981), .ZN(new_n1014));
  INV_X1    g589(.A(G1981), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n708), .A2(KEYINPUT110), .A3(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n595), .B(KEYINPUT111), .ZN(new_n1018));
  OAI21_X1  g593(.A(G1981), .B1(new_n1018), .B2(new_n599), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT49), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n993), .B1(new_n940), .B2(new_n944), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1017), .A2(new_n1019), .A3(KEYINPUT49), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n591), .A2(G1976), .ZN(new_n1026));
  AOI21_X1  g601(.A(KEYINPUT52), .B1(new_n1023), .B2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(KEYINPUT109), .B1(new_n591), .B2(G1976), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1023), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n1023), .B(new_n1028), .C1(KEYINPUT52), .C2(new_n1026), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  AND2_X1   g607(.A1(new_n1025), .A2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1007), .A2(new_n1012), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  NOR2_X1   g610(.A1(G168), .A2(new_n993), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1036), .ZN(new_n1037));
  OAI211_X1 g612(.A(new_n944), .B(new_n978), .C1(new_n940), .C2(KEYINPUT45), .ZN(new_n1038));
  INV_X1    g613(.A(G1966), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(KEYINPUT113), .ZN(new_n1041));
  OR2_X1    g616(.A1(new_n970), .A2(G2084), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT113), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1038), .A2(new_n1043), .A3(new_n1039), .ZN(new_n1044));
  AND3_X1   g619(.A1(new_n1041), .A2(new_n1042), .A3(new_n1044), .ZN(new_n1045));
  OAI211_X1 g620(.A(KEYINPUT51), .B(new_n1037), .C1(new_n1045), .C2(new_n993), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT51), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1041), .A2(new_n1042), .A3(new_n1044), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n1047), .B(G8), .C1(new_n1048), .C2(G286), .ZN(new_n1049));
  AND3_X1   g624(.A1(new_n1048), .A2(KEYINPUT122), .A3(new_n1036), .ZN(new_n1050));
  AOI21_X1  g625(.A(KEYINPUT122), .B1(new_n1048), .B2(new_n1036), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1046), .B(new_n1049), .C1(new_n1050), .C2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1035), .A2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n959), .B1(new_n992), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(new_n753), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n970), .A2(new_n1055), .ZN(new_n1056));
  AND3_X1   g631(.A1(new_n940), .A2(new_n952), .A3(new_n944), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT117), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n940), .A2(new_n944), .ZN(new_n1060));
  OAI21_X1  g635(.A(KEYINPUT117), .B1(new_n1060), .B2(G2067), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1056), .A2(new_n1059), .A3(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(KEYINPUT118), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT118), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1056), .A2(new_n1059), .A3(new_n1064), .A4(new_n1061), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n615), .A2(KEYINPUT121), .ZN(new_n1067));
  OR2_X1    g642(.A1(new_n615), .A2(KEYINPUT121), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1066), .A2(KEYINPUT60), .A3(new_n1067), .A4(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT60), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1063), .A2(new_n1065), .A3(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1070), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n1069), .B(new_n1071), .C1(new_n1067), .C2(new_n1072), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n960), .A2(new_n963), .A3(new_n954), .A4(new_n944), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT120), .ZN(new_n1075));
  XOR2_X1   g650(.A(KEYINPUT58), .B(G1341), .Z(new_n1076));
  NAND2_X1  g651(.A1(new_n1060), .A2(new_n1076), .ZN(new_n1077));
  AND3_X1   g652(.A1(new_n1074), .A2(new_n1075), .A3(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1075), .B1(new_n1074), .B2(new_n1077), .ZN(new_n1079));
  NOR3_X1   g654(.A1(new_n1078), .A2(new_n1079), .A3(new_n562), .ZN(new_n1080));
  XOR2_X1   g655(.A(new_n1080), .B(KEYINPUT59), .Z(new_n1081));
  INV_X1    g656(.A(KEYINPUT61), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n996), .A2(new_n998), .A3(new_n999), .ZN(new_n1083));
  XNOR2_X1  g658(.A(KEYINPUT114), .B(G1956), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  XOR2_X1   g660(.A(KEYINPUT56), .B(G2072), .Z(new_n1086));
  OR2_X1    g661(.A1(new_n1001), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1088), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n575), .A2(KEYINPUT115), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT115), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1091), .B1(new_n571), .B2(new_n574), .ZN(new_n1092));
  OR3_X1    g667(.A1(new_n1090), .A2(new_n581), .A3(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT57), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(KEYINPUT116), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT116), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1093), .A2(new_n1097), .A3(new_n1094), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1096), .B(new_n1098), .C1(new_n1094), .C2(G299), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1082), .B1(new_n1089), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1089), .A2(new_n1099), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1089), .A2(new_n1082), .A3(new_n1099), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1073), .A2(new_n1081), .A3(new_n1102), .A4(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1099), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT119), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1105), .A2(new_n1106), .A3(new_n1088), .ZN(new_n1107));
  OAI21_X1  g682(.A(KEYINPUT119), .B1(new_n1089), .B2(new_n1099), .ZN(new_n1108));
  OAI211_X1 g683(.A(new_n1107), .B(new_n1108), .C1(new_n615), .C2(new_n1066), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(new_n1101), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1104), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(new_n983), .ZN(new_n1112));
  AOI21_X1  g687(.A(G301), .B1(new_n988), .B2(new_n989), .ZN(new_n1113));
  OAI21_X1  g688(.A(KEYINPUT54), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1114), .B1(new_n980), .B2(new_n977), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1115), .A2(KEYINPUT124), .A3(new_n1035), .A4(new_n1052), .ZN(new_n1116));
  AND3_X1   g691(.A1(new_n1054), .A2(new_n1111), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1033), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1118), .A2(new_n1012), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1023), .ZN(new_n1120));
  INV_X1    g695(.A(G1976), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1025), .A2(new_n1121), .A3(new_n591), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1120), .B1(new_n1122), .B2(new_n1017), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT63), .ZN(new_n1124));
  NOR3_X1   g699(.A1(new_n1045), .A2(new_n993), .A3(G286), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1125), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1124), .B1(new_n1034), .B2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1006), .B1(new_n1011), .B2(G8), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1128), .A2(new_n1124), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1129), .A2(new_n1012), .A3(new_n1033), .A4(new_n1125), .ZN(new_n1130));
  AOI211_X1 g705(.A(new_n1119), .B(new_n1123), .C1(new_n1127), .C2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1052), .A2(KEYINPUT62), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1132), .A2(KEYINPUT125), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT125), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1052), .A2(new_n1134), .A3(KEYINPUT62), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1136));
  OAI211_X1 g711(.A(new_n1035), .B(new_n980), .C1(new_n1052), .C2(KEYINPUT62), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1131), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n958), .B1(new_n1117), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(new_n953), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n949), .B1(new_n743), .B2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n949), .A2(KEYINPUT46), .A3(new_n954), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT46), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1143), .B1(new_n948), .B2(G1996), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1141), .A2(new_n1142), .A3(new_n1144), .ZN(new_n1145));
  XOR2_X1   g720(.A(new_n1145), .B(KEYINPUT47), .Z(new_n1146));
  NAND4_X1  g721(.A1(new_n955), .A2(new_n730), .A3(new_n728), .A4(new_n953), .ZN(new_n1147));
  OR2_X1    g722(.A1(new_n795), .A2(G2067), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n948), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NOR3_X1   g724(.A1(new_n948), .A2(G1986), .A3(G290), .ZN(new_n1150));
  XNOR2_X1  g725(.A(new_n1150), .B(KEYINPUT48), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1151), .B1(new_n949), .B2(new_n956), .ZN(new_n1152));
  NOR3_X1   g727(.A1(new_n1146), .A2(new_n1149), .A3(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1139), .A2(new_n1153), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g729(.A1(G229), .A2(new_n464), .ZN(new_n1156));
  NAND3_X1  g730(.A1(new_n1156), .A2(new_n676), .A3(new_n659), .ZN(new_n1157));
  INV_X1    g731(.A(KEYINPUT126), .ZN(new_n1158));
  NAND2_X1  g732(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NAND4_X1  g733(.A1(new_n1156), .A2(new_n676), .A3(new_n659), .A4(KEYINPUT126), .ZN(new_n1160));
  AOI22_X1  g734(.A1(new_n867), .A2(new_n869), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g735(.A1(new_n928), .A2(new_n1161), .ZN(G225));
  NAND2_X1  g736(.A1(G225), .A2(KEYINPUT127), .ZN(new_n1163));
  INV_X1    g737(.A(KEYINPUT127), .ZN(new_n1164));
  NAND3_X1  g738(.A1(new_n928), .A2(new_n1161), .A3(new_n1164), .ZN(new_n1165));
  NAND2_X1  g739(.A1(new_n1163), .A2(new_n1165), .ZN(G308));
endmodule


