//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 0 1 0 1 0 0 0 0 1 0 0 1 0 1 1 0 1 0 0 0 1 0 0 1 0 0 0 0 1 1 1 0 1 1 1 1 1 1 0 1 1 1 1 0 0 1 0 0 0 0 0 0 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:08 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1067, new_n1068, new_n1069, new_n1070, new_n1071, new_n1072,
    new_n1073, new_n1074, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1129, new_n1130, new_n1131, new_n1132, new_n1133,
    new_n1134, new_n1135, new_n1136, new_n1137, new_n1138, new_n1139,
    new_n1140, new_n1141, new_n1142, new_n1143, new_n1144, new_n1145,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1160, new_n1161, new_n1162, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  XOR2_X1   g0003(.A(KEYINPUT65), .B(G244), .Z(new_n204));
  INV_X1    g0004(.A(G77), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G58), .A2(G232), .B1(G87), .B2(G250), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G50), .A2(G226), .B1(G107), .B2(G264), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G68), .A2(G238), .B1(G97), .B2(G257), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G116), .A2(G270), .ZN(new_n210));
  NAND4_X1  g0010(.A1(new_n207), .A2(new_n208), .A3(new_n209), .A4(new_n210), .ZN(new_n211));
  OAI21_X1  g0011(.A(new_n203), .B1(new_n206), .B2(new_n211), .ZN(new_n212));
  OR2_X1    g0012(.A1(new_n212), .A2(KEYINPUT1), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n212), .A2(KEYINPUT1), .ZN(new_n214));
  OAI21_X1  g0014(.A(G50), .B1(G58), .B2(G68), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  NAND3_X1  g0018(.A1(new_n216), .A2(G20), .A3(new_n218), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n203), .A2(G13), .ZN(new_n220));
  OAI211_X1 g0020(.A(new_n220), .B(G250), .C1(G257), .C2(G264), .ZN(new_n221));
  XOR2_X1   g0021(.A(KEYINPUT64), .B(KEYINPUT0), .Z(new_n222));
  XNOR2_X1  g0022(.A(new_n221), .B(new_n222), .ZN(new_n223));
  AND4_X1   g0023(.A1(new_n213), .A2(new_n214), .A3(new_n219), .A4(new_n223), .ZN(G361));
  XNOR2_X1  g0024(.A(G250), .B(G257), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT66), .ZN(new_n226));
  XOR2_X1   g0026(.A(G264), .B(G270), .Z(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  INV_X1    g0029(.A(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n228), .B(new_n233), .Z(G358));
  XOR2_X1   g0034(.A(G68), .B(G77), .Z(new_n235));
  XNOR2_X1  g0035(.A(G50), .B(G58), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G351));
  XNOR2_X1  g0041(.A(KEYINPUT15), .B(G87), .ZN(new_n242));
  INV_X1    g0042(.A(new_n242), .ZN(new_n243));
  INV_X1    g0043(.A(G33), .ZN(new_n244));
  NOR2_X1   g0044(.A1(new_n244), .A2(G20), .ZN(new_n245));
  AOI22_X1  g0045(.A1(new_n243), .A2(new_n245), .B1(G20), .B2(G77), .ZN(new_n246));
  NOR2_X1   g0046(.A1(G20), .A2(G33), .ZN(new_n247));
  INV_X1    g0047(.A(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(KEYINPUT8), .B(G58), .ZN(new_n249));
  OAI21_X1  g0049(.A(new_n246), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  OAI21_X1  g0050(.A(new_n217), .B1(new_n203), .B2(new_n244), .ZN(new_n251));
  INV_X1    g0051(.A(G1), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n252), .A2(G13), .A3(G20), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(KEYINPUT70), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT70), .ZN(new_n255));
  NAND4_X1  g0055(.A1(new_n255), .A2(new_n252), .A3(G13), .A4(G20), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  AOI22_X1  g0058(.A1(new_n250), .A2(new_n251), .B1(new_n205), .B2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n251), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n252), .A2(G20), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n262), .A2(G77), .A3(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n259), .A2(new_n264), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n217), .B1(G33), .B2(G41), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT3), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(new_n244), .ZN(new_n269));
  NAND2_X1  g0069(.A1(KEYINPUT3), .A2(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n230), .A2(G1698), .ZN(new_n272));
  INV_X1    g0072(.A(G238), .ZN(new_n273));
  INV_X1    g0073(.A(G1698), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n271), .B1(new_n272), .B2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G107), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n276), .B1(new_n277), .B2(new_n271), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT72), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n267), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n280), .B1(new_n279), .B2(new_n278), .ZN(new_n281));
  INV_X1    g0081(.A(G274), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n252), .B1(G41), .B2(G45), .ZN(new_n283));
  OR3_X1    g0083(.A1(new_n266), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(new_n204), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n267), .A2(new_n283), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n285), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n281), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n265), .B1(new_n291), .B2(G190), .ZN(new_n292));
  INV_X1    g0092(.A(G200), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n292), .B1(new_n293), .B2(new_n291), .ZN(new_n294));
  INV_X1    g0094(.A(G179), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n291), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G169), .ZN(new_n297));
  AOI22_X1  g0097(.A1(new_n290), .A2(new_n297), .B1(new_n264), .B2(new_n259), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  AND2_X1   g0099(.A1(new_n294), .A2(new_n299), .ZN(new_n300));
  OR2_X1    g0100(.A1(new_n300), .A2(KEYINPUT73), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(KEYINPUT73), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n271), .A2(G222), .A3(new_n274), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT67), .ZN(new_n304));
  XNOR2_X1  g0104(.A(new_n303), .B(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n271), .A2(G1698), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  AND2_X1   g0107(.A1(KEYINPUT3), .A2(G33), .ZN(new_n308));
  NOR2_X1   g0108(.A1(KEYINPUT3), .A2(G33), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  AOI22_X1  g0110(.A1(new_n307), .A2(G223), .B1(G77), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n305), .A2(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n267), .B1(new_n312), .B2(KEYINPUT68), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n313), .B1(KEYINPUT68), .B2(new_n312), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n285), .B1(G226), .B2(new_n288), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(new_n297), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT69), .ZN(new_n318));
  XNOR2_X1  g0118(.A(new_n249), .B(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n245), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(G150), .ZN(new_n322));
  NOR3_X1   g0122(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n323));
  INV_X1    g0123(.A(G20), .ZN(new_n324));
  OAI22_X1  g0124(.A1(new_n322), .A2(new_n248), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n251), .B1(new_n321), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n263), .A2(G50), .ZN(new_n327));
  XNOR2_X1  g0127(.A(new_n327), .B(KEYINPUT71), .ZN(new_n328));
  INV_X1    g0128(.A(G50), .ZN(new_n329));
  AOI22_X1  g0129(.A1(new_n262), .A2(new_n328), .B1(new_n329), .B2(new_n258), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n326), .A2(new_n330), .ZN(new_n331));
  OAI211_X1 g0131(.A(new_n317), .B(new_n331), .C1(G179), .C2(new_n316), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n301), .A2(new_n302), .A3(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT74), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n273), .B1(new_n287), .B2(new_n334), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n335), .B1(new_n334), .B2(new_n287), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n230), .A2(G1698), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n271), .B(new_n337), .C1(G226), .C2(G1698), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(G97), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n244), .A2(new_n340), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n266), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n336), .A2(new_n284), .A3(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT13), .ZN(new_n344));
  XNOR2_X1  g0144(.A(new_n343), .B(new_n344), .ZN(new_n345));
  OR3_X1    g0145(.A1(new_n345), .A2(KEYINPUT14), .A3(new_n297), .ZN(new_n346));
  OAI21_X1  g0146(.A(KEYINPUT14), .B1(new_n345), .B2(new_n297), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n345), .A2(G179), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  OAI22_X1  g0149(.A1(new_n320), .A2(new_n205), .B1(new_n324), .B2(G68), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT76), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n350), .A2(new_n351), .B1(G50), .B2(new_n247), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n352), .B1(new_n351), .B2(new_n350), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(new_n251), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  OR2_X1    g0155(.A1(new_n355), .A2(KEYINPUT11), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(KEYINPUT11), .ZN(new_n357));
  INV_X1    g0157(.A(G68), .ZN(new_n358));
  INV_X1    g0158(.A(new_n263), .ZN(new_n359));
  NOR3_X1   g0159(.A1(new_n261), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  OAI21_X1  g0160(.A(KEYINPUT12), .B1(new_n257), .B2(G68), .ZN(new_n361));
  OR3_X1    g0161(.A1(new_n257), .A2(KEYINPUT12), .A3(G68), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n360), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n356), .A2(new_n357), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n349), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n345), .A2(G190), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT75), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n345), .A2(KEYINPUT75), .A3(G190), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n345), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n364), .B1(new_n371), .B2(G200), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n365), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(KEYINPUT77), .B1(new_n308), .B2(new_n309), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT77), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n269), .A2(new_n376), .A3(new_n270), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n375), .A2(new_n377), .A3(new_n324), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT7), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n271), .A2(G20), .ZN(new_n381));
  XOR2_X1   g0181(.A(KEYINPUT78), .B(KEYINPUT7), .Z(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n380), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(G68), .ZN(new_n385));
  INV_X1    g0185(.A(G58), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n386), .A2(new_n358), .ZN(new_n387));
  NOR2_X1   g0187(.A1(G58), .A2(G68), .ZN(new_n388));
  OAI21_X1  g0188(.A(G20), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n247), .A2(G159), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT16), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n260), .B1(new_n385), .B2(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n310), .A2(KEYINPUT7), .A3(new_n324), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n395), .B1(new_n381), .B2(new_n382), .ZN(new_n396));
  AND2_X1   g0196(.A1(new_n396), .A2(G68), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n392), .B1(new_n397), .B2(new_n391), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n394), .A2(new_n398), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n319), .A2(new_n359), .ZN(new_n400));
  AOI22_X1  g0200(.A1(new_n400), .A2(new_n262), .B1(new_n258), .B2(new_n319), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n284), .B1(new_n230), .B2(new_n287), .ZN(new_n403));
  OR2_X1    g0203(.A1(new_n274), .A2(G226), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n271), .B(new_n404), .C1(G223), .C2(G1698), .ZN(new_n405));
  NAND2_X1  g0205(.A1(G33), .A2(G87), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n267), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n403), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(G179), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n409), .B1(new_n297), .B2(new_n408), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n402), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT18), .ZN(new_n412));
  XNOR2_X1  g0212(.A(new_n411), .B(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n408), .A2(G190), .ZN(new_n414));
  OAI21_X1  g0214(.A(G200), .B1(new_n403), .B2(new_n407), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n399), .A2(new_n401), .A3(new_n414), .A4(new_n415), .ZN(new_n416));
  XNOR2_X1  g0216(.A(new_n416), .B(KEYINPUT17), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n413), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n314), .A2(G190), .A3(new_n315), .ZN(new_n419));
  XNOR2_X1  g0219(.A(new_n331), .B(KEYINPUT9), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n293), .B1(new_n314), .B2(new_n315), .ZN(new_n422));
  OAI21_X1  g0222(.A(KEYINPUT10), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n316), .A2(G200), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT10), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n424), .A2(new_n425), .A3(new_n419), .A4(new_n420), .ZN(new_n426));
  AND2_X1   g0226(.A1(new_n423), .A2(new_n426), .ZN(new_n427));
  NOR4_X1   g0227(.A1(new_n333), .A2(new_n374), .A3(new_n418), .A4(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n277), .A2(KEYINPUT6), .A3(G97), .ZN(new_n429));
  OR2_X1    g0229(.A1(new_n429), .A2(KEYINPUT79), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(KEYINPUT79), .ZN(new_n431));
  XOR2_X1   g0231(.A(G97), .B(G107), .Z(new_n432));
  OAI211_X1 g0232(.A(new_n430), .B(new_n431), .C1(new_n432), .C2(KEYINPUT6), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(G20), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n434), .B1(new_n205), .B2(new_n248), .ZN(new_n435));
  AND2_X1   g0235(.A1(new_n396), .A2(G107), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n251), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n257), .A2(G97), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n261), .B1(new_n252), .B2(G33), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n438), .B1(new_n439), .B2(G97), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n437), .A2(new_n440), .ZN(new_n441));
  XNOR2_X1  g0241(.A(new_n441), .B(KEYINPUT80), .ZN(new_n442));
  XNOR2_X1  g0242(.A(KEYINPUT5), .B(G41), .ZN(new_n443));
  INV_X1    g0243(.A(G45), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n444), .A2(G1), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  NOR3_X1   g0246(.A1(new_n446), .A2(new_n282), .A3(new_n266), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n266), .B1(new_n445), .B2(new_n443), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(G257), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n448), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n271), .A2(G244), .A3(new_n274), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT81), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  XNOR2_X1  g0255(.A(new_n455), .B(KEYINPUT4), .ZN(new_n456));
  NAND2_X1  g0256(.A1(G33), .A2(G283), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n271), .A2(G250), .A3(G1698), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  OR3_X1    g0260(.A1(new_n456), .A2(new_n458), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n452), .B1(new_n461), .B2(new_n266), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n442), .B1(G190), .B2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT82), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n461), .A2(new_n464), .A3(new_n266), .ZN(new_n465));
  NOR3_X1   g0265(.A1(new_n456), .A2(new_n458), .A3(new_n460), .ZN(new_n466));
  OAI21_X1  g0266(.A(KEYINPUT82), .B1(new_n466), .B2(new_n267), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n452), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  OR2_X1    g0268(.A1(new_n468), .A2(new_n293), .ZN(new_n469));
  INV_X1    g0269(.A(new_n462), .ZN(new_n470));
  AOI22_X1  g0270(.A1(new_n468), .A2(new_n295), .B1(new_n470), .B2(new_n297), .ZN(new_n471));
  AOI22_X1  g0271(.A1(new_n463), .A2(new_n469), .B1(new_n471), .B2(new_n441), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n271), .A2(new_n324), .A3(G87), .ZN(new_n473));
  XNOR2_X1  g0273(.A(new_n473), .B(KEYINPUT22), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT23), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n475), .B1(new_n324), .B2(G107), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n277), .A2(KEYINPUT23), .A3(G20), .ZN(new_n477));
  AOI22_X1  g0277(.A1(new_n476), .A2(new_n477), .B1(new_n245), .B2(G116), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n474), .A2(new_n478), .ZN(new_n479));
  XNOR2_X1  g0279(.A(new_n479), .B(KEYINPUT24), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(new_n251), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT25), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n482), .B1(new_n257), .B2(G107), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n258), .A2(KEYINPUT25), .A3(new_n277), .ZN(new_n484));
  AOI22_X1  g0284(.A1(new_n439), .A2(G107), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n481), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n271), .A2(G250), .A3(new_n274), .ZN(new_n487));
  INV_X1    g0287(.A(G294), .ZN(new_n488));
  OAI221_X1 g0288(.A(new_n487), .B1(new_n244), .B2(new_n488), .C1(new_n306), .C2(new_n451), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n447), .B1(new_n489), .B2(new_n266), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n449), .A2(G264), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(G169), .ZN(new_n493));
  XNOR2_X1  g0293(.A(new_n491), .B(KEYINPUT83), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(new_n490), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n493), .B1(new_n295), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n486), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(KEYINPUT84), .ZN(new_n498));
  INV_X1    g0298(.A(new_n486), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n495), .A2(new_n293), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n500), .B1(G190), .B2(new_n492), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT84), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n486), .A2(new_n496), .A3(new_n503), .ZN(new_n504));
  AND3_X1   g0304(.A1(new_n498), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(new_n439), .ZN(new_n506));
  INV_X1    g0306(.A(G116), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n457), .B(new_n324), .C1(G33), .C2(new_n340), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n509), .B(new_n251), .C1(new_n324), .C2(G116), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT20), .ZN(new_n511));
  AND2_X1   g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n510), .A2(new_n511), .ZN(new_n513));
  OAI22_X1  g0313(.A1(new_n512), .A2(new_n513), .B1(G116), .B2(new_n257), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n508), .A2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT21), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n271), .A2(G257), .A3(new_n274), .ZN(new_n517));
  INV_X1    g0317(.A(G303), .ZN(new_n518));
  INV_X1    g0318(.A(G264), .ZN(new_n519));
  OAI221_X1 g0319(.A(new_n517), .B1(new_n518), .B2(new_n271), .C1(new_n306), .C2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n266), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n447), .B1(G270), .B2(new_n449), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(G169), .ZN(new_n524));
  OR3_X1    g0324(.A1(new_n515), .A2(new_n516), .A3(new_n524), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n516), .B1(new_n515), .B2(new_n524), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n523), .A2(new_n295), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n527), .B1(new_n508), .B2(new_n514), .ZN(new_n528));
  AND3_X1   g0328(.A1(new_n525), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n523), .A2(G200), .ZN(new_n530));
  INV_X1    g0330(.A(G190), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n515), .B(new_n530), .C1(new_n531), .C2(new_n523), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n271), .A2(new_n324), .A3(G68), .ZN(new_n533));
  AOI21_X1  g0333(.A(G20), .B1(new_n341), .B2(KEYINPUT19), .ZN(new_n534));
  NOR3_X1   g0334(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n320), .A2(new_n340), .ZN(new_n536));
  OAI221_X1 g0336(.A(new_n533), .B1(new_n534), .B2(new_n535), .C1(new_n536), .C2(KEYINPUT19), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n537), .A2(new_n251), .B1(new_n258), .B2(new_n242), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n439), .A2(G87), .ZN(new_n539));
  AND2_X1   g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n445), .A2(new_n282), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n267), .B(new_n541), .C1(G250), .C2(new_n445), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n273), .A2(new_n274), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n271), .B(new_n544), .C1(G244), .C2(new_n274), .ZN(new_n545));
  NAND2_X1  g0345(.A1(G33), .A2(G116), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n267), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n543), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(G190), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n540), .B(new_n549), .C1(new_n293), .C2(new_n548), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n538), .B1(new_n242), .B2(new_n506), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n548), .A2(new_n295), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n551), .B(new_n552), .C1(G169), .C2(new_n548), .ZN(new_n553));
  AND2_X1   g0353(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  AND3_X1   g0354(.A1(new_n529), .A2(new_n532), .A3(new_n554), .ZN(new_n555));
  AND3_X1   g0355(.A1(new_n472), .A2(new_n505), .A3(new_n555), .ZN(new_n556));
  AND2_X1   g0356(.A1(new_n428), .A2(new_n556), .ZN(G372));
  INV_X1    g0357(.A(KEYINPUT85), .ZN(new_n558));
  OR2_X1    g0358(.A1(new_n547), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n547), .A2(new_n558), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n543), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n540), .B(new_n549), .C1(new_n561), .C2(new_n293), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n551), .B(new_n552), .C1(new_n561), .C2(G169), .ZN(new_n563));
  AND2_X1   g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AND2_X1   g0364(.A1(new_n502), .A2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT86), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n529), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n525), .A2(new_n526), .A3(new_n528), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(KEYINPUT86), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(new_n497), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n472), .B(new_n565), .C1(new_n571), .C2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n468), .A2(new_n295), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n470), .A2(new_n297), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n574), .A2(new_n554), .A3(new_n575), .A4(new_n441), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(KEYINPUT26), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT26), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n471), .A2(new_n564), .A3(new_n578), .A4(new_n442), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n577), .A2(new_n563), .A3(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n573), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n428), .A2(new_n582), .ZN(new_n583));
  XOR2_X1   g0383(.A(new_n583), .B(KEYINPUT87), .Z(new_n584));
  AND3_X1   g0384(.A1(new_n423), .A2(KEYINPUT88), .A3(new_n426), .ZN(new_n585));
  AOI21_X1  g0385(.A(KEYINPUT88), .B1(new_n423), .B2(new_n426), .ZN(new_n586));
  OR2_X1    g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  XOR2_X1   g0387(.A(new_n416), .B(KEYINPUT17), .Z(new_n588));
  INV_X1    g0388(.A(new_n299), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n373), .A2(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n588), .B1(new_n590), .B2(new_n365), .ZN(new_n591));
  XNOR2_X1  g0391(.A(new_n411), .B(KEYINPUT18), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n587), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n332), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT89), .ZN(new_n595));
  XNOR2_X1  g0395(.A(new_n594), .B(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n584), .A2(new_n596), .ZN(new_n597));
  XOR2_X1   g0397(.A(new_n597), .B(KEYINPUT90), .Z(G369));
  NAND3_X1  g0398(.A1(new_n252), .A2(new_n324), .A3(G13), .ZN(new_n599));
  OR2_X1    g0399(.A1(new_n599), .A2(KEYINPUT27), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(KEYINPUT27), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n600), .A2(G213), .A3(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(G343), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n515), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n571), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n529), .A2(new_n532), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n607), .B1(new_n608), .B2(new_n606), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n609), .A2(G330), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n505), .B1(new_n499), .B2(new_n605), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n611), .B1(new_n497), .B2(new_n605), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n529), .A2(new_n604), .ZN(new_n614));
  AOI22_X1  g0414(.A1(new_n505), .A2(new_n614), .B1(new_n572), .B2(new_n605), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n613), .A2(new_n615), .ZN(G399));
  INV_X1    g0416(.A(new_n220), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n617), .A2(G41), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n535), .A2(new_n507), .ZN(new_n619));
  NOR3_X1   g0419(.A1(new_n618), .A2(new_n619), .A3(new_n252), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n620), .B1(new_n216), .B2(new_n618), .ZN(new_n621));
  XOR2_X1   g0421(.A(new_n621), .B(KEYINPUT28), .Z(new_n622));
  INV_X1    g0422(.A(G330), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n489), .A2(new_n266), .ZN(new_n624));
  AND4_X1   g0424(.A1(new_n624), .A2(new_n527), .A3(new_n494), .A4(new_n548), .ZN(new_n625));
  AOI21_X1  g0425(.A(KEYINPUT91), .B1(new_n625), .B2(new_n462), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT30), .ZN(new_n627));
  INV_X1    g0427(.A(new_n561), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n628), .A2(new_n295), .A3(new_n495), .A4(new_n523), .ZN(new_n629));
  OAI22_X1  g0429(.A1(new_n626), .A2(new_n627), .B1(new_n468), .B2(new_n629), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n626), .A2(new_n627), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n604), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT31), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT92), .ZN(new_n635));
  AOI22_X1  g0435(.A1(new_n556), .A2(new_n605), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  OAI211_X1 g0436(.A(KEYINPUT31), .B(new_n604), .C1(new_n630), .C2(new_n631), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n634), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(KEYINPUT92), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n623), .B1(new_n636), .B2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT29), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n576), .A2(new_n578), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(KEYINPUT93), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT93), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n576), .A2(new_n644), .A3(new_n578), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n471), .A2(new_n564), .A3(KEYINPUT26), .A4(new_n442), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n643), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n498), .A2(new_n504), .A3(new_n529), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n472), .A2(new_n565), .A3(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n647), .A2(new_n563), .A3(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n641), .B1(new_n650), .B2(new_n605), .ZN(new_n651));
  AOI211_X1 g0451(.A(KEYINPUT29), .B(new_n604), .C1(new_n573), .C2(new_n581), .ZN(new_n652));
  NOR3_X1   g0452(.A1(new_n640), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n622), .B1(new_n653), .B2(G1), .ZN(G364));
  AND2_X1   g0454(.A1(new_n324), .A2(G13), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n252), .B1(new_n655), .B2(G45), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n657), .A2(new_n618), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(G13), .A2(G33), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n661), .A2(G20), .ZN(new_n662));
  XNOR2_X1  g0462(.A(new_n662), .B(KEYINPUT94), .ZN(new_n663));
  OR2_X1    g0463(.A1(new_n609), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n663), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n217), .B1(G20), .B2(new_n297), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n216), .A2(new_n444), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n375), .A2(new_n377), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n670), .A2(new_n617), .ZN(new_n671));
  OAI211_X1 g0471(.A(new_n669), .B(new_n671), .C1(new_n237), .C2(new_n444), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n617), .A2(new_n310), .ZN(new_n673));
  AOI22_X1  g0473(.A1(new_n673), .A2(G355), .B1(new_n507), .B2(new_n617), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n668), .B1(new_n672), .B2(new_n674), .ZN(new_n675));
  NOR2_X1   g0475(.A1(G179), .A2(G200), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n324), .B1(new_n676), .B2(G190), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(G97), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n324), .A2(new_n295), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(G200), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n681), .A2(new_n531), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n681), .A2(G190), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  OAI221_X1 g0485(.A(new_n679), .B1(new_n683), .B2(new_n329), .C1(new_n358), .C2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT95), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n687), .B1(new_n324), .B2(G190), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n293), .A2(G179), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n531), .A2(KEYINPUT95), .A3(G20), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n688), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n691), .A2(new_n277), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n324), .A2(new_n531), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(new_n689), .ZN(new_n694));
  INV_X1    g0494(.A(G87), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n271), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n693), .A2(G179), .A3(new_n293), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n680), .A2(new_n531), .A3(new_n293), .ZN(new_n698));
  OAI22_X1  g0498(.A1(new_n697), .A2(new_n386), .B1(new_n698), .B2(new_n205), .ZN(new_n699));
  OR4_X1    g0499(.A1(new_n686), .A2(new_n692), .A3(new_n696), .A4(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n688), .A2(new_n676), .A3(new_n690), .ZN(new_n701));
  INV_X1    g0501(.A(G159), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g0503(.A(KEYINPUT96), .B(KEYINPUT32), .ZN(new_n704));
  XNOR2_X1  g0504(.A(new_n703), .B(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(G322), .ZN(new_n706));
  INV_X1    g0506(.A(G311), .ZN(new_n707));
  OAI22_X1  g0507(.A1(new_n697), .A2(new_n706), .B1(new_n698), .B2(new_n707), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n708), .B1(G326), .B2(new_n682), .ZN(new_n709));
  XNOR2_X1  g0509(.A(KEYINPUT33), .B(G317), .ZN(new_n710));
  AOI22_X1  g0510(.A1(new_n684), .A2(new_n710), .B1(G294), .B2(new_n678), .ZN(new_n711));
  INV_X1    g0511(.A(new_n691), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(G283), .ZN(new_n713));
  INV_X1    g0513(.A(new_n701), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(G329), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n709), .A2(new_n711), .A3(new_n713), .A4(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n310), .B1(new_n694), .B2(new_n518), .ZN(new_n717));
  XNOR2_X1  g0517(.A(new_n717), .B(KEYINPUT97), .ZN(new_n718));
  OAI22_X1  g0518(.A1(new_n700), .A2(new_n705), .B1(new_n716), .B2(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n675), .B1(new_n719), .B2(new_n666), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n659), .B1(new_n664), .B2(new_n720), .ZN(new_n721));
  XNOR2_X1  g0521(.A(new_n609), .B(G330), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n721), .B1(new_n659), .B2(new_n722), .ZN(new_n723));
  XNOR2_X1  g0523(.A(new_n723), .B(KEYINPUT98), .ZN(G396));
  NAND2_X1  g0524(.A1(new_n582), .A2(new_n605), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n265), .A2(new_n604), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n589), .B1(new_n294), .B2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n299), .A2(new_n604), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n725), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n463), .A2(new_n469), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n471), .A2(new_n441), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n565), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n572), .B1(new_n567), .B2(new_n569), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  OAI211_X1 g0536(.A(new_n605), .B(new_n729), .C1(new_n736), .C2(new_n580), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n640), .B1(new_n731), .B2(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(new_n658), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n731), .A2(new_n640), .A3(new_n737), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n666), .A2(new_n660), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n659), .B1(new_n205), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n679), .B1(new_n683), .B2(new_n518), .ZN(new_n744));
  OAI22_X1  g0544(.A1(new_n698), .A2(new_n507), .B1(new_n694), .B2(new_n277), .ZN(new_n745));
  INV_X1    g0545(.A(new_n697), .ZN(new_n746));
  AOI211_X1 g0546(.A(new_n271), .B(new_n745), .C1(G294), .C2(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n712), .A2(G87), .ZN(new_n748));
  OAI211_X1 g0548(.A(new_n747), .B(new_n748), .C1(new_n707), .C2(new_n701), .ZN(new_n749));
  AOI211_X1 g0549(.A(new_n744), .B(new_n749), .C1(G283), .C2(new_n684), .ZN(new_n750));
  AOI22_X1  g0550(.A1(G137), .A2(new_n682), .B1(new_n684), .B2(G150), .ZN(new_n751));
  XNOR2_X1  g0551(.A(new_n751), .B(KEYINPUT99), .ZN(new_n752));
  XNOR2_X1  g0552(.A(KEYINPUT100), .B(G143), .ZN(new_n753));
  OAI221_X1 g0553(.A(new_n752), .B1(new_n702), .B2(new_n698), .C1(new_n697), .C2(new_n753), .ZN(new_n754));
  XNOR2_X1  g0554(.A(new_n754), .B(KEYINPUT34), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n691), .A2(new_n358), .ZN(new_n756));
  OAI221_X1 g0556(.A(new_n670), .B1(new_n329), .B2(new_n694), .C1(new_n386), .C2(new_n677), .ZN(new_n757));
  AOI211_X1 g0557(.A(new_n756), .B(new_n757), .C1(G132), .C2(new_n714), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n750), .B1(new_n755), .B2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n666), .ZN(new_n760));
  OAI221_X1 g0560(.A(new_n743), .B1(new_n759), .B2(new_n760), .C1(new_n729), .C2(new_n661), .ZN(new_n761));
  AND2_X1   g0561(.A1(new_n741), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(G384));
  OAI21_X1  g0563(.A(new_n428), .B1(new_n651), .B2(new_n652), .ZN(new_n764));
  AND2_X1   g0564(.A1(new_n596), .A2(new_n764), .ZN(new_n765));
  XOR2_X1   g0565(.A(new_n765), .B(KEYINPUT107), .Z(new_n766));
  INV_X1    g0566(.A(KEYINPUT102), .ZN(new_n767));
  INV_X1    g0567(.A(new_n319), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(new_n263), .ZN(new_n769));
  OAI22_X1  g0569(.A1(new_n769), .A2(new_n261), .B1(new_n257), .B2(new_n768), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n358), .B1(new_n380), .B2(new_n383), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n392), .B1(new_n771), .B2(new_n391), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n770), .B1(new_n394), .B2(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n767), .B1(new_n773), .B2(new_n602), .ZN(new_n774));
  INV_X1    g0574(.A(new_n391), .ZN(new_n775));
  AOI21_X1  g0575(.A(KEYINPUT16), .B1(new_n385), .B2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n393), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n251), .B1(new_n771), .B2(new_n777), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n401), .B1(new_n776), .B2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n602), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n779), .A2(KEYINPUT102), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n779), .A2(new_n410), .ZN(new_n782));
  NAND4_X1  g0582(.A1(new_n774), .A2(new_n781), .A3(new_n416), .A4(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(KEYINPUT37), .ZN(new_n784));
  INV_X1    g0584(.A(KEYINPUT103), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n783), .A2(KEYINPUT103), .A3(KEYINPUT37), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n402), .A2(new_n780), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n411), .A2(new_n788), .A3(new_n416), .ZN(new_n789));
  OR2_X1    g0589(.A1(new_n789), .A2(KEYINPUT37), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n786), .A2(new_n787), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n774), .A2(new_n781), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n792), .B1(new_n588), .B2(new_n592), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n791), .A2(KEYINPUT38), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(KEYINPUT104), .ZN(new_n795));
  AOI21_X1  g0595(.A(KEYINPUT38), .B1(new_n791), .B2(new_n793), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(KEYINPUT104), .ZN(new_n798));
  INV_X1    g0598(.A(KEYINPUT38), .ZN(new_n799));
  AND3_X1   g0599(.A1(new_n783), .A2(KEYINPUT103), .A3(KEYINPUT37), .ZN(new_n800));
  AOI21_X1  g0600(.A(KEYINPUT103), .B1(new_n783), .B2(KEYINPUT37), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n789), .A2(KEYINPUT37), .ZN(new_n802));
  NOR3_X1   g0602(.A1(new_n800), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n413), .A2(new_n417), .B1(new_n774), .B2(new_n781), .ZN(new_n804));
  OAI211_X1 g0604(.A(new_n798), .B(new_n799), .C1(new_n803), .C2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  OAI21_X1  g0606(.A(KEYINPUT39), .B1(new_n797), .B2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(KEYINPUT105), .ZN(new_n808));
  XOR2_X1   g0608(.A(new_n789), .B(KEYINPUT37), .Z(new_n809));
  AOI21_X1  g0609(.A(new_n788), .B1(new_n413), .B2(new_n417), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n799), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  AND2_X1   g0611(.A1(new_n811), .A2(new_n794), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(KEYINPUT39), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n807), .A2(new_n808), .A3(new_n815), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n349), .A2(new_n364), .A3(new_n605), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n799), .B1(new_n803), .B2(new_n804), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n819), .A2(KEYINPUT104), .A3(new_n794), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n814), .B1(new_n820), .B2(new_n805), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n812), .A2(KEYINPUT39), .ZN(new_n822));
  OAI21_X1  g0622(.A(KEYINPUT105), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n816), .A2(new_n818), .A3(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n797), .A2(new_n806), .ZN(new_n825));
  AND2_X1   g0625(.A1(new_n370), .A2(new_n372), .ZN(new_n826));
  OAI211_X1 g0626(.A(new_n364), .B(new_n604), .C1(new_n826), .C2(new_n349), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n364), .A2(new_n604), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n365), .A2(new_n373), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n728), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n831), .B1(new_n737), .B2(new_n832), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n825), .A2(new_n833), .B1(new_n592), .B2(new_n602), .ZN(new_n834));
  AND3_X1   g0634(.A1(new_n824), .A2(KEYINPUT106), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(KEYINPUT106), .B1(new_n824), .B2(new_n834), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n766), .B(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n730), .B1(new_n827), .B2(new_n829), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n472), .A2(new_n505), .A3(new_n555), .A4(new_n605), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n840), .A2(new_n634), .A3(new_n637), .ZN(new_n841));
  AND2_X1   g0641(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT40), .ZN(new_n843));
  NAND4_X1  g0643(.A1(new_n842), .A2(new_n843), .A3(new_n805), .A4(new_n820), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n839), .A2(new_n841), .ZN(new_n845));
  OAI21_X1  g0645(.A(KEYINPUT40), .B1(new_n845), .B2(new_n812), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  AND2_X1   g0647(.A1(new_n428), .A2(new_n841), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n847), .A2(new_n848), .ZN(new_n851));
  NOR3_X1   g0651(.A1(new_n850), .A2(new_n851), .A3(new_n623), .ZN(new_n852));
  OAI22_X1  g0652(.A1(new_n838), .A2(new_n852), .B1(new_n252), .B2(new_n655), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n853), .B1(new_n838), .B2(new_n852), .ZN(new_n854));
  NOR3_X1   g0654(.A1(new_n217), .A2(new_n324), .A3(new_n507), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n433), .B(KEYINPUT101), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT35), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n855), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n859), .B1(new_n858), .B2(new_n857), .ZN(new_n860));
  XNOR2_X1  g0660(.A(new_n860), .B(KEYINPUT36), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n216), .B(G77), .C1(new_n386), .C2(new_n358), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n329), .A2(G68), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n252), .B(G13), .C1(new_n862), .C2(new_n863), .ZN(new_n864));
  OR3_X1    g0664(.A1(new_n854), .A2(new_n861), .A3(new_n864), .ZN(G367));
  OAI21_X1  g0665(.A(new_n667), .B1(new_n220), .B2(new_n242), .ZN(new_n866));
  INV_X1    g0666(.A(new_n671), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n228), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n658), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  XNOR2_X1  g0669(.A(new_n869), .B(KEYINPUT112), .ZN(new_n870));
  INV_X1    g0670(.A(new_n698), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n746), .A2(G150), .B1(new_n871), .B2(G50), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n714), .A2(G137), .ZN(new_n873));
  INV_X1    g0673(.A(new_n694), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n310), .B1(new_n874), .B2(G58), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n872), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n691), .A2(new_n205), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n684), .A2(G159), .B1(G68), .B2(new_n678), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n878), .B(new_n879), .C1(new_n683), .C2(new_n753), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT46), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n881), .B1(new_n694), .B2(new_n507), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n874), .A2(KEYINPUT46), .A3(G116), .ZN(new_n883));
  OAI211_X1 g0683(.A(new_n882), .B(new_n883), .C1(new_n685), .C2(new_n488), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT113), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  OAI22_X1  g0686(.A1(new_n683), .A2(new_n707), .B1(new_n677), .B2(new_n277), .ZN(new_n887));
  INV_X1    g0687(.A(G283), .ZN(new_n888));
  OAI22_X1  g0688(.A1(new_n697), .A2(new_n518), .B1(new_n698), .B2(new_n888), .ZN(new_n889));
  NOR3_X1   g0689(.A1(new_n887), .A2(new_n670), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n884), .A2(new_n885), .ZN(new_n891));
  AOI22_X1  g0691(.A1(G97), .A2(new_n712), .B1(new_n714), .B2(G317), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n880), .B1(new_n886), .B2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT47), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n894), .A2(new_n895), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n666), .ZN(new_n898));
  OR2_X1    g0698(.A1(new_n540), .A2(new_n605), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n564), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n900), .B1(new_n563), .B2(new_n899), .ZN(new_n901));
  OAI221_X1 g0701(.A(new_n870), .B1(new_n896), .B2(new_n898), .C1(new_n901), .C2(new_n663), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n442), .A2(new_n604), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n472), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n471), .A2(new_n442), .A3(new_n604), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g0706(.A1(KEYINPUT110), .A2(KEYINPUT44), .ZN(new_n907));
  NOR3_X1   g0707(.A1(new_n906), .A2(new_n615), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(KEYINPUT110), .A2(KEYINPUT44), .ZN(new_n909));
  XOR2_X1   g0709(.A(new_n908), .B(new_n909), .Z(new_n910));
  NAND2_X1  g0710(.A1(new_n906), .A2(new_n615), .ZN(new_n911));
  XOR2_X1   g0711(.A(new_n911), .B(KEYINPUT45), .Z(new_n912));
  NAND2_X1  g0712(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  XOR2_X1   g0713(.A(new_n913), .B(new_n613), .Z(new_n914));
  NAND2_X1  g0714(.A1(new_n505), .A2(new_n614), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT111), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n505), .A2(KEYINPUT111), .A3(new_n614), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n917), .B(new_n918), .C1(new_n612), .C2(new_n614), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n610), .B(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n653), .ZN(new_n921));
  OR2_X1    g0721(.A1(new_n914), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(new_n653), .ZN(new_n923));
  XOR2_X1   g0723(.A(new_n618), .B(KEYINPUT41), .Z(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n657), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  XOR2_X1   g0726(.A(new_n906), .B(KEYINPUT108), .Z(new_n927));
  NOR2_X1   g0727(.A1(new_n613), .A2(new_n927), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n928), .B(KEYINPUT109), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n901), .A2(KEYINPUT43), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n929), .B(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(new_n927), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n498), .A2(new_n504), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n604), .B1(new_n934), .B2(new_n733), .ZN(new_n935));
  INV_X1    g0735(.A(new_n906), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n936), .A2(new_n915), .ZN(new_n937));
  XOR2_X1   g0737(.A(new_n937), .B(KEYINPUT42), .Z(new_n938));
  NOR2_X1   g0738(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n939), .B1(KEYINPUT43), .B2(new_n901), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n931), .B(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n902), .B1(new_n926), .B2(new_n941), .ZN(G387));
  OR2_X1    g0742(.A1(new_n612), .A2(new_n663), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n673), .A2(new_n619), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n944), .B1(G107), .B2(new_n220), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n867), .B1(new_n233), .B2(G45), .ZN(new_n946));
  OAI221_X1 g0746(.A(new_n444), .B1(new_n358), .B2(new_n205), .C1(new_n619), .C2(KEYINPUT114), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n947), .B1(KEYINPUT114), .B2(new_n619), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n249), .A2(G50), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(KEYINPUT50), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n945), .B1(new_n946), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n658), .B1(new_n952), .B2(new_n668), .ZN(new_n953));
  XOR2_X1   g0753(.A(new_n953), .B(KEYINPUT115), .Z(new_n954));
  INV_X1    g0754(.A(new_n670), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n955), .B1(G77), .B2(new_n874), .ZN(new_n956));
  OAI221_X1 g0756(.A(new_n956), .B1(new_n340), .B2(new_n691), .C1(new_n322), .C2(new_n701), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(KEYINPUT116), .ZN(new_n958));
  AOI22_X1  g0758(.A1(new_n746), .A2(G50), .B1(new_n871), .B2(G68), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n678), .A2(new_n243), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n959), .B(new_n960), .C1(new_n702), .C2(new_n683), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n961), .B1(new_n768), .B2(new_n684), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n958), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n670), .B1(G326), .B2(new_n714), .ZN(new_n964));
  OAI22_X1  g0764(.A1(new_n694), .A2(new_n488), .B1(new_n677), .B2(new_n888), .ZN(new_n965));
  AOI22_X1  g0765(.A1(new_n746), .A2(G317), .B1(new_n871), .B2(G303), .ZN(new_n966));
  OAI221_X1 g0766(.A(new_n966), .B1(new_n707), .B2(new_n685), .C1(new_n706), .C2(new_n683), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT48), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n965), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(new_n968), .B2(new_n967), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT49), .ZN(new_n971));
  OAI221_X1 g0771(.A(new_n964), .B1(new_n507), .B2(new_n691), .C1(new_n970), .C2(new_n971), .ZN(new_n972));
  AND2_X1   g0772(.A1(new_n970), .A2(new_n971), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n963), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n954), .B1(new_n666), .B2(new_n974), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n920), .A2(new_n657), .B1(new_n943), .B2(new_n975), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n921), .A2(KEYINPUT117), .A3(new_n618), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n977), .B1(new_n653), .B2(new_n920), .ZN(new_n978));
  AOI21_X1  g0778(.A(KEYINPUT117), .B1(new_n921), .B2(new_n618), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n976), .B1(new_n978), .B2(new_n979), .ZN(G393));
  AND2_X1   g0780(.A1(new_n922), .A2(new_n618), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n914), .A2(new_n921), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  OR2_X1    g0783(.A1(new_n914), .A2(new_n656), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n667), .B1(new_n340), .B2(new_n220), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n867), .A2(new_n240), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n658), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n683), .A2(new_n322), .B1(new_n702), .B2(new_n697), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT51), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n698), .A2(new_n249), .B1(new_n694), .B2(new_n358), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n990), .A2(new_n955), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n677), .A2(new_n205), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n992), .B1(new_n684), .B2(G50), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n748), .B1(new_n701), .B2(new_n753), .ZN(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n989), .A2(new_n991), .A3(new_n993), .A4(new_n995), .ZN(new_n996));
  AOI22_X1  g0796(.A1(G317), .A2(new_n682), .B1(new_n746), .B2(G311), .ZN(new_n997));
  XOR2_X1   g0797(.A(new_n997), .B(KEYINPUT52), .Z(new_n998));
  AOI211_X1 g0798(.A(new_n271), .B(new_n692), .C1(G283), .C2(new_n874), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n998), .B(new_n999), .C1(new_n706), .C2(new_n701), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n871), .A2(G294), .B1(new_n678), .B2(G116), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n518), .B2(new_n685), .ZN(new_n1002));
  XOR2_X1   g0802(.A(new_n1002), .B(KEYINPUT118), .Z(new_n1003));
  OAI21_X1  g0803(.A(new_n996), .B1(new_n1000), .B2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n987), .B1(new_n1004), .B2(new_n666), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n932), .B2(new_n663), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n983), .A2(new_n984), .A3(new_n1006), .ZN(G390));
  AOI21_X1  g0807(.A(new_n808), .B1(new_n807), .B2(new_n815), .ZN(new_n1008));
  NOR3_X1   g0808(.A1(new_n821), .A2(new_n822), .A3(KEYINPUT105), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n1008), .A2(new_n1009), .B1(new_n818), .B2(new_n833), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n645), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n644), .B1(new_n576), .B2(new_n578), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n646), .ZN(new_n1013));
  NOR3_X1   g0813(.A1(new_n1011), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n649), .A2(new_n563), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n605), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n832), .B1(new_n1016), .B2(new_n727), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1017), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n817), .B(new_n813), .C1(new_n1018), .C2(new_n831), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n640), .A2(new_n729), .A3(new_n830), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1010), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n841), .A2(G330), .ZN(new_n1022));
  NOR3_X1   g0822(.A1(new_n1022), .A2(new_n730), .A3(new_n831), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n833), .A2(new_n818), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1024), .B1(new_n816), .B2(new_n823), .ZN(new_n1025));
  AOI211_X1 g0825(.A(new_n818), .B(new_n812), .C1(new_n1017), .C2(new_n830), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1023), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1021), .A2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n428), .A2(G330), .A3(new_n841), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n596), .A2(new_n764), .A3(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n737), .A2(new_n832), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n830), .B1(new_n640), .B2(new_n729), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1031), .B1(new_n1032), .B2(new_n1023), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n831), .B1(new_n1022), .B2(new_n730), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1018), .A2(new_n1020), .A3(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1030), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1028), .A2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1021), .A2(new_n1027), .A3(new_n1036), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1038), .A2(new_n618), .A3(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n659), .B1(new_n319), .B2(new_n742), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n271), .B1(new_n874), .B2(G87), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n1042), .B1(new_n340), .B2(new_n698), .C1(new_n507), .C2(new_n697), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n756), .B(new_n1043), .C1(G294), .C2(new_n714), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n683), .A2(new_n888), .ZN(new_n1045));
  AOI211_X1 g0845(.A(new_n992), .B(new_n1045), .C1(G107), .C2(new_n684), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n694), .A2(new_n322), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT53), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n1047), .A2(new_n1048), .B1(new_n702), .B2(new_n677), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(G137), .B2(new_n684), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1051));
  INV_X1    g0851(.A(G128), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1051), .B1(new_n683), .B2(new_n1052), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(KEYINPUT54), .B(G143), .ZN(new_n1054));
  INV_X1    g0854(.A(G132), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n271), .B1(new_n698), .B2(new_n1054), .C1(new_n1055), .C2(new_n697), .ZN(new_n1056));
  INV_X1    g0856(.A(G125), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n329), .A2(new_n691), .B1(new_n701), .B2(new_n1057), .ZN(new_n1058));
  NOR3_X1   g0858(.A1(new_n1053), .A2(new_n1056), .A3(new_n1058), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n1044), .A2(new_n1046), .B1(new_n1050), .B2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1041), .B1(new_n1060), .B2(new_n760), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n816), .A2(new_n823), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1061), .B1(new_n1062), .B2(new_n660), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT119), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1021), .A2(new_n1027), .A3(new_n657), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1040), .A2(new_n1064), .A3(new_n1065), .ZN(G378));
  INV_X1    g0866(.A(KEYINPUT57), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1030), .ZN(new_n1068));
  AND2_X1   g0868(.A1(new_n1039), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n824), .A2(new_n834), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT106), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n824), .A2(KEYINPUT106), .A3(new_n834), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n623), .B1(new_n844), .B2(new_n846), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n332), .B1(new_n585), .B2(new_n586), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n331), .A2(new_n780), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1076), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1081), .B(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1074), .A2(new_n1084), .ZN(new_n1085));
  OR2_X1    g0885(.A1(new_n1074), .A2(new_n1084), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n1072), .A2(new_n1073), .A3(new_n1085), .A4(new_n1086), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1074), .B(new_n1084), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n835), .B2(new_n836), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1067), .B1(new_n1069), .B2(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT121), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1039), .A2(new_n1068), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n1094), .A2(KEYINPUT57), .A3(new_n1087), .A4(new_n1089), .ZN(new_n1095));
  AND2_X1   g0895(.A1(new_n1095), .A2(new_n618), .ZN(new_n1096));
  OAI211_X1 g0896(.A(KEYINPUT121), .B(new_n1067), .C1(new_n1069), .C2(new_n1090), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1093), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1087), .A2(new_n1089), .A3(new_n657), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n659), .B1(new_n329), .B2(new_n742), .ZN(new_n1100));
  OR2_X1    g0900(.A1(new_n670), .A2(G41), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(G77), .B2(new_n874), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n712), .A2(G58), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1102), .B(new_n1103), .C1(new_n888), .C2(new_n701), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n1104), .B(KEYINPUT120), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n277), .A2(new_n697), .B1(new_n698), .B2(new_n242), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1106), .B1(G68), .B2(new_n678), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(G97), .A2(new_n684), .B1(new_n682), .B2(G116), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1105), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT58), .ZN(new_n1110));
  OR2_X1    g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n685), .A2(new_n1055), .B1(new_n683), .B2(new_n1057), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1112), .B1(G150), .B2(new_n678), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1054), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n871), .A2(G137), .B1(new_n874), .B2(new_n1114), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n1113), .B(new_n1115), .C1(new_n1052), .C2(new_n697), .ZN(new_n1116));
  OR2_X1    g0916(.A1(new_n1116), .A2(KEYINPUT59), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(G33), .A2(G41), .ZN(new_n1118));
  INV_X1    g0918(.A(G124), .ZN(new_n1119));
  OAI221_X1 g0919(.A(new_n1118), .B1(new_n691), .B2(new_n702), .C1(new_n1119), .C2(new_n701), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1120), .B1(new_n1116), .B2(KEYINPUT59), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1118), .A2(G50), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n1117), .A2(new_n1121), .B1(new_n1101), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1111), .A2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1124), .B1(new_n1110), .B2(new_n1109), .ZN(new_n1125));
  OAI221_X1 g0925(.A(new_n1100), .B1(new_n760), .B2(new_n1125), .C1(new_n1084), .C2(new_n661), .ZN(new_n1126));
  AND2_X1   g0926(.A1(new_n1099), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1098), .A2(new_n1127), .ZN(G375));
  AND2_X1   g0928(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(new_n656), .B(KEYINPUT122), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n659), .B1(new_n358), .B2(new_n742), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n871), .A2(G107), .B1(new_n874), .B2(G97), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n1134), .B(new_n310), .C1(new_n888), .C2(new_n697), .ZN(new_n1135));
  AOI211_X1 g0935(.A(new_n877), .B(new_n1135), .C1(G303), .C2(new_n714), .ZN(new_n1136));
  OAI221_X1 g0936(.A(new_n960), .B1(new_n683), .B2(new_n488), .C1(new_n507), .C2(new_n685), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n1055), .A2(new_n683), .B1(new_n685), .B2(new_n1054), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n955), .B(new_n1139), .C1(G50), .C2(new_n678), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n746), .A2(G137), .B1(new_n874), .B2(G159), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n1141), .B(new_n1103), .C1(new_n322), .C2(new_n698), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1142), .B1(G128), .B2(new_n714), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n1136), .A2(new_n1138), .B1(new_n1140), .B2(new_n1143), .ZN(new_n1144));
  OAI221_X1 g0944(.A(new_n1133), .B1(new_n760), .B2(new_n1144), .C1(new_n830), .C2(new_n661), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1132), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1129), .A2(new_n1030), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1148), .A2(new_n1037), .A3(new_n925), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1147), .A2(new_n1149), .ZN(G381));
  AND2_X1   g0950(.A1(G375), .A2(KEYINPUT124), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(G375), .A2(KEYINPUT124), .ZN(new_n1152));
  NOR3_X1   g0952(.A1(new_n1151), .A2(new_n1152), .A3(G378), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(G387), .A2(G390), .ZN(new_n1154));
  OR2_X1    g0954(.A1(G393), .A2(G396), .ZN(new_n1155));
  NOR3_X1   g0955(.A1(G381), .A2(new_n1155), .A3(G384), .ZN(new_n1156));
  AOI21_X1  g0956(.A(KEYINPUT123), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1157));
  AND3_X1   g0957(.A1(new_n1154), .A2(KEYINPUT123), .A3(new_n1156), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1153), .B1(new_n1157), .B2(new_n1158), .ZN(G407));
  NAND2_X1  g0959(.A1(new_n603), .A2(G213), .ZN(new_n1160));
  XOR2_X1   g0960(.A(new_n1160), .B(KEYINPUT125), .Z(new_n1161));
  NAND2_X1  g0961(.A1(new_n1153), .A2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(G407), .A2(G213), .A3(new_n1162), .ZN(G409));
  INV_X1    g0963(.A(KEYINPUT61), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1098), .A2(G378), .A3(new_n1127), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1131), .B1(new_n1094), .B2(new_n925), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1126), .B1(new_n1166), .B2(new_n1090), .ZN(new_n1167));
  INV_X1    g0967(.A(G378), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1161), .B1(new_n1165), .B2(new_n1169), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1148), .A2(KEYINPUT60), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT60), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(new_n1129), .B2(new_n1030), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n618), .B(new_n1037), .C1(new_n1171), .C2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(new_n1147), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1175), .A2(new_n762), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1174), .A2(G384), .A3(new_n1147), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n1176), .A2(new_n1177), .B1(G2897), .B2(new_n1161), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1160), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(G2897), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1178), .B1(new_n1180), .B2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1164), .B1(new_n1170), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(KEYINPUT126), .ZN(new_n1186));
  AND2_X1   g0986(.A1(new_n1180), .A2(KEYINPUT62), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1170), .A2(new_n1187), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n1181), .B(new_n1179), .C1(new_n1165), .C2(new_n1169), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1188), .B1(new_n1189), .B2(KEYINPUT62), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT126), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n1191), .B(new_n1164), .C1(new_n1170), .C2(new_n1184), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1186), .A2(new_n1190), .A3(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1154), .ZN(new_n1194));
  XOR2_X1   g0994(.A(G393), .B(G396), .Z(new_n1195));
  NAND2_X1  g0995(.A1(G387), .A2(G390), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1194), .A2(new_n1195), .A3(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1195), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1196), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1198), .B1(new_n1199), .B2(new_n1154), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1197), .A2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1193), .A2(new_n1202), .ZN(new_n1203));
  OR2_X1    g1003(.A1(new_n1189), .A2(KEYINPUT63), .ZN(new_n1204));
  AOI21_X1  g1004(.A(KEYINPUT61), .B1(new_n1197), .B2(new_n1200), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1170), .A2(KEYINPUT63), .A3(new_n1180), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1181), .B1(new_n1165), .B2(new_n1169), .ZN(new_n1207));
  OR2_X1    g1007(.A1(new_n1207), .A2(new_n1184), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1204), .A2(new_n1205), .A3(new_n1206), .A4(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1203), .A2(new_n1209), .ZN(G405));
  INV_X1    g1010(.A(KEYINPUT127), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1165), .ZN(new_n1212));
  AOI21_X1  g1012(.A(G378), .B1(new_n1098), .B2(new_n1127), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1211), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1213), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1215), .A2(KEYINPUT127), .A3(new_n1165), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1179), .B1(new_n1214), .B2(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1214), .A2(new_n1216), .A3(new_n1179), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1218), .A2(new_n1202), .A3(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1219), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1201), .B1(new_n1221), .B2(new_n1217), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1220), .A2(new_n1222), .ZN(G402));
endmodule


