//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 1 1 1 0 1 0 1 1 1 1 0 1 0 1 0 1 1 1 0 1 0 1 1 0 1 0 1 1 0 1 1 1 0 0 0 1 0 0 1 0 1 0 1 1 0 1 0 1 1 1 0 1 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:01 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n728, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n929,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974;
  INV_X1    g000(.A(G104), .ZN(new_n187));
  OAI21_X1  g001(.A(KEYINPUT3), .B1(new_n187), .B2(G107), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT3), .ZN(new_n189));
  INV_X1    g003(.A(G107), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(new_n190), .A3(G104), .ZN(new_n191));
  INV_X1    g005(.A(G101), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n187), .A2(G107), .ZN(new_n193));
  NAND4_X1  g007(.A1(new_n188), .A2(new_n191), .A3(new_n192), .A4(new_n193), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n187), .A2(G107), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n190), .A2(G104), .ZN(new_n196));
  OAI21_X1  g010(.A(G101), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n194), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  NOR2_X1   g013(.A1(KEYINPUT67), .A2(G119), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(KEYINPUT67), .A2(G119), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n201), .A2(G116), .A3(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G119), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n204), .A2(G116), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n203), .A2(KEYINPUT5), .A3(new_n206), .ZN(new_n207));
  AND2_X1   g021(.A1(KEYINPUT67), .A2(G119), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n208), .A2(new_n200), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT5), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n209), .A2(new_n210), .A3(G116), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n207), .A2(G113), .A3(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT68), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n205), .B1(new_n209), .B2(G116), .ZN(new_n214));
  XOR2_X1   g028(.A(KEYINPUT2), .B(G113), .Z(new_n215));
  AOI21_X1  g029(.A(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  AND4_X1   g030(.A1(new_n213), .A2(new_n203), .A3(new_n215), .A4(new_n206), .ZN(new_n217));
  OAI211_X1 g031(.A(new_n199), .B(new_n212), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n214), .A2(new_n215), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n203), .A2(new_n215), .A3(new_n206), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(KEYINPUT68), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n214), .A2(new_n213), .A3(new_n215), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n219), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n188), .A2(new_n191), .A3(new_n193), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G101), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n225), .A2(KEYINPUT4), .A3(new_n194), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT4), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n224), .A2(new_n227), .A3(G101), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n218), .B1(new_n223), .B2(new_n229), .ZN(new_n230));
  XNOR2_X1  g044(.A(G110), .B(G122), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  OAI211_X1 g047(.A(new_n218), .B(new_n231), .C1(new_n223), .C2(new_n229), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n233), .A2(KEYINPUT6), .A3(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT6), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n230), .A2(new_n236), .A3(new_n232), .ZN(new_n237));
  INV_X1    g051(.A(G143), .ZN(new_n238));
  OAI21_X1  g052(.A(KEYINPUT1), .B1(new_n238), .B2(G146), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n238), .A2(G146), .ZN(new_n240));
  INV_X1    g054(.A(G146), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n241), .A2(G143), .ZN(new_n242));
  OAI211_X1 g056(.A(G128), .B(new_n239), .C1(new_n240), .C2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(G125), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n241), .A2(G143), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n238), .A2(G146), .ZN(new_n246));
  INV_X1    g060(.A(G128), .ZN(new_n247));
  OAI211_X1 g061(.A(new_n245), .B(new_n246), .C1(KEYINPUT1), .C2(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n243), .A2(new_n244), .A3(new_n248), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n245), .A2(new_n246), .A3(KEYINPUT0), .A4(G128), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n240), .A2(new_n242), .ZN(new_n251));
  XNOR2_X1  g065(.A(KEYINPUT0), .B(G128), .ZN(new_n252));
  OAI211_X1 g066(.A(new_n250), .B(G125), .C1(new_n251), .C2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n249), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(G953), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G224), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n254), .B(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n235), .A2(new_n237), .A3(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n256), .A2(KEYINPUT85), .A3(KEYINPUT7), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n256), .A2(KEYINPUT7), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT85), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n260), .B1(new_n254), .B2(new_n263), .ZN(new_n264));
  AOI211_X1 g078(.A(new_n262), .B(new_n261), .C1(new_n249), .C2(new_n253), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AND2_X1   g080(.A1(new_n234), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g081(.A(new_n231), .B(KEYINPUT8), .ZN(new_n268));
  INV_X1    g082(.A(new_n218), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n221), .A2(new_n222), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n199), .B1(new_n270), .B2(new_n212), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n268), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(G902), .B1(new_n267), .B2(new_n272), .ZN(new_n273));
  OAI21_X1  g087(.A(G210), .B1(G237), .B2(G902), .ZN(new_n274));
  AND3_X1   g088(.A1(new_n258), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  XOR2_X1   g089(.A(new_n274), .B(KEYINPUT86), .Z(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n277), .B1(new_n258), .B2(new_n273), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n275), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(G214), .B1(G237), .B2(G902), .ZN(new_n281));
  XOR2_X1   g095(.A(new_n281), .B(KEYINPUT84), .Z(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n280), .A2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G469), .ZN(new_n285));
  INV_X1    g099(.A(G902), .ZN(new_n286));
  XNOR2_X1  g100(.A(G110), .B(G140), .ZN(new_n287));
  AND2_X1   g101(.A1(new_n255), .A2(G227), .ZN(new_n288));
  XNOR2_X1  g102(.A(new_n287), .B(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n250), .B1(new_n251), .B2(new_n252), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n226), .A2(new_n292), .A3(new_n228), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT81), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n226), .A2(new_n292), .A3(KEYINPUT81), .A4(new_n228), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n243), .A2(new_n194), .A3(new_n197), .A4(new_n248), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT10), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n298), .B1(KEYINPUT82), .B2(new_n299), .ZN(new_n300));
  XNOR2_X1  g114(.A(KEYINPUT82), .B(KEYINPUT10), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n300), .B1(new_n298), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n297), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G137), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n305), .A2(KEYINPUT11), .A3(G134), .ZN(new_n306));
  INV_X1    g120(.A(G134), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(G137), .ZN(new_n308));
  AND2_X1   g122(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT64), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n305), .A2(G134), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT11), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n310), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  AOI211_X1 g127(.A(KEYINPUT64), .B(KEYINPUT11), .C1(new_n305), .C2(G134), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n309), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G131), .ZN(new_n316));
  INV_X1    g130(.A(G131), .ZN(new_n317));
  OAI211_X1 g131(.A(new_n309), .B(new_n317), .C1(new_n313), .C2(new_n314), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n316), .A2(KEYINPUT65), .A3(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT65), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n315), .A2(new_n320), .A3(G131), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n304), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n297), .A2(new_n303), .A3(new_n322), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n290), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n243), .A2(new_n248), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(new_n198), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(new_n298), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n319), .A2(new_n329), .A3(new_n321), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT12), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n319), .A2(new_n329), .A3(KEYINPUT12), .A4(new_n321), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AND3_X1   g148(.A1(new_n325), .A2(new_n334), .A3(new_n290), .ZN(new_n335));
  OAI211_X1 g149(.A(new_n285), .B(new_n286), .C1(new_n326), .C2(new_n335), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n285), .A2(new_n286), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n325), .A2(new_n334), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(new_n289), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n324), .A2(new_n325), .A3(new_n290), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n340), .A2(new_n341), .A3(G469), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n336), .A2(new_n338), .A3(new_n342), .ZN(new_n343));
  XNOR2_X1  g157(.A(KEYINPUT9), .B(G234), .ZN(new_n344));
  OAI21_X1  g158(.A(G221), .B1(new_n344), .B2(G902), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(KEYINPUT83), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT83), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n343), .A2(new_n348), .A3(new_n345), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n284), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(G140), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(G125), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n244), .A2(G140), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT76), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n352), .A2(new_n353), .A3(new_n354), .A4(KEYINPUT16), .ZN(new_n355));
  AND3_X1   g169(.A1(new_n352), .A2(new_n353), .A3(KEYINPUT16), .ZN(new_n356));
  OAI21_X1  g170(.A(KEYINPUT76), .B1(new_n352), .B2(KEYINPUT16), .ZN(new_n357));
  OAI211_X1 g171(.A(new_n241), .B(new_n355), .C1(new_n356), .C2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n352), .A2(new_n353), .A3(KEYINPUT16), .ZN(new_n360));
  OR3_X1    g174(.A1(new_n244), .A2(KEYINPUT16), .A3(G140), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n360), .A2(new_n361), .A3(KEYINPUT76), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n241), .B1(new_n362), .B2(new_n355), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n359), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(G237), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n365), .A2(new_n255), .A3(G214), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(new_n238), .ZN(new_n367));
  NOR2_X1   g181(.A1(G237), .A2(G953), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n368), .A2(G143), .A3(G214), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(KEYINPUT88), .B1(new_n370), .B2(G131), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT88), .ZN(new_n372));
  AOI211_X1 g186(.A(new_n372), .B(new_n317), .C1(new_n367), .C2(new_n369), .ZN(new_n373));
  OAI21_X1  g187(.A(KEYINPUT17), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  AND4_X1   g188(.A1(G143), .A2(new_n365), .A3(new_n255), .A4(G214), .ZN(new_n375));
  AOI21_X1  g189(.A(G143), .B1(new_n368), .B2(G214), .ZN(new_n376));
  OAI21_X1  g190(.A(G131), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(new_n372), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n370), .A2(KEYINPUT88), .A3(G131), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n367), .A2(new_n317), .A3(new_n369), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(KEYINPUT87), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT87), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n367), .A2(new_n382), .A3(new_n317), .A4(new_n369), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n378), .A2(new_n379), .A3(new_n381), .A4(new_n383), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n364), .B(new_n374), .C1(new_n384), .C2(KEYINPUT17), .ZN(new_n385));
  XNOR2_X1  g199(.A(G113), .B(G122), .ZN(new_n386));
  XNOR2_X1  g200(.A(new_n386), .B(KEYINPUT90), .ZN(new_n387));
  XNOR2_X1  g201(.A(KEYINPUT89), .B(G104), .ZN(new_n388));
  XNOR2_X1  g202(.A(new_n387), .B(new_n388), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n244), .A2(G140), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n351), .A2(G125), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  XNOR2_X1  g206(.A(new_n392), .B(new_n241), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n370), .A2(KEYINPUT18), .A3(G131), .ZN(new_n394));
  NAND2_X1  g208(.A1(KEYINPUT18), .A2(G131), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n367), .A2(new_n369), .A3(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n393), .A2(new_n394), .A3(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n385), .A2(new_n389), .A3(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT19), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n399), .B1(new_n390), .B2(new_n391), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n352), .A2(new_n353), .A3(KEYINPUT19), .ZN(new_n401));
  AOI21_X1  g215(.A(G146), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n355), .B1(new_n356), .B2(new_n357), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n402), .B1(G146), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n384), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n397), .ZN(new_n406));
  INV_X1    g220(.A(new_n389), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n398), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT91), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NOR2_X1   g225(.A1(G475), .A2(G902), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n398), .A2(new_n408), .A3(KEYINPUT91), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(KEYINPUT20), .ZN(new_n415));
  INV_X1    g229(.A(new_n412), .ZN(new_n416));
  AOI211_X1 g230(.A(KEYINPUT20), .B(new_n416), .C1(new_n398), .C2(new_n408), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT92), .ZN(new_n419));
  AND3_X1   g233(.A1(new_n385), .A2(new_n389), .A3(new_n397), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n389), .B1(new_n385), .B2(new_n397), .ZN(new_n421));
  OAI211_X1 g235(.A(new_n419), .B(new_n286), .C1(new_n420), .C2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(G475), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n286), .B1(new_n420), .B2(new_n421), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n423), .B1(new_n424), .B2(KEYINPUT92), .ZN(new_n425));
  AOI22_X1  g239(.A1(new_n415), .A2(new_n418), .B1(new_n422), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n255), .A2(G952), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n427), .B1(G234), .B2(G237), .ZN(new_n428));
  NAND2_X1  g242(.A1(G234), .A2(G237), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n429), .A2(G902), .A3(G953), .ZN(new_n430));
  XOR2_X1   g244(.A(new_n430), .B(KEYINPUT93), .Z(new_n431));
  XNOR2_X1  g245(.A(KEYINPUT21), .B(G898), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n428), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n238), .A2(G128), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n247), .A2(G143), .ZN(new_n436));
  AND2_X1   g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n437), .B(new_n307), .ZN(new_n438));
  XNOR2_X1  g252(.A(G116), .B(G122), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(new_n190), .ZN(new_n440));
  INV_X1    g254(.A(G116), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n441), .A2(KEYINPUT14), .A3(G122), .ZN(new_n442));
  INV_X1    g256(.A(new_n439), .ZN(new_n443));
  OAI211_X1 g257(.A(G107), .B(new_n442), .C1(new_n443), .C2(KEYINPUT14), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n438), .A2(new_n440), .A3(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n435), .ZN(new_n446));
  AND2_X1   g260(.A1(new_n446), .A2(KEYINPUT13), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n436), .B1(new_n446), .B2(KEYINPUT13), .ZN(new_n448));
  OAI21_X1  g262(.A(G134), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n437), .A2(new_n307), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n439), .B(new_n190), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(G217), .ZN(new_n453));
  NOR3_X1   g267(.A1(new_n344), .A2(new_n453), .A3(G953), .ZN(new_n454));
  AND3_X1   g268(.A1(new_n445), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n454), .B1(new_n445), .B2(new_n452), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n457), .A2(G902), .ZN(new_n458));
  INV_X1    g272(.A(G478), .ZN(new_n459));
  OR2_X1    g273(.A1(new_n459), .A2(KEYINPUT15), .ZN(new_n460));
  XOR2_X1   g274(.A(new_n458), .B(new_n460), .Z(new_n461));
  NAND3_X1  g275(.A1(new_n426), .A2(new_n434), .A3(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  AND2_X1   g277(.A1(new_n350), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g278(.A1(G472), .A2(G902), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n319), .A2(new_n292), .A3(new_n321), .ZN(new_n466));
  INV_X1    g280(.A(new_n327), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n311), .A2(new_n308), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(G131), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n467), .A2(new_n318), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n466), .A2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT30), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(KEYINPUT66), .ZN(new_n474));
  INV_X1    g288(.A(new_n223), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n318), .A2(new_n469), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(KEYINPUT69), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT69), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n318), .A2(new_n478), .A3(new_n469), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n477), .A2(new_n467), .A3(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n480), .A2(new_n466), .A3(KEYINPUT30), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT66), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n471), .A2(new_n482), .A3(new_n472), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n474), .A2(new_n475), .A3(new_n481), .A4(new_n483), .ZN(new_n484));
  AND3_X1   g298(.A1(new_n480), .A2(new_n466), .A3(new_n223), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n368), .A2(G210), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n486), .B(KEYINPUT27), .ZN(new_n487));
  XNOR2_X1  g301(.A(KEYINPUT26), .B(G101), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n487), .B(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n485), .A2(new_n490), .ZN(new_n491));
  XOR2_X1   g305(.A(KEYINPUT70), .B(KEYINPUT31), .Z(new_n492));
  NAND3_X1  g306(.A1(new_n484), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(KEYINPUT71), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT71), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n484), .A2(new_n495), .A3(new_n491), .A4(new_n492), .ZN(new_n496));
  AND2_X1   g310(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n223), .B1(new_n466), .B2(new_n470), .ZN(new_n498));
  OAI21_X1  g312(.A(KEYINPUT28), .B1(new_n485), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n480), .A2(new_n466), .A3(new_n223), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT28), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(KEYINPUT72), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT72), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n500), .A2(new_n504), .A3(new_n501), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n499), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(new_n490), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT73), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n484), .A2(new_n491), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(KEYINPUT31), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n506), .A2(KEYINPUT73), .A3(new_n490), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n509), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n465), .B1(new_n497), .B2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT32), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n494), .A2(new_n496), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n517), .A2(new_n511), .A3(new_n512), .A4(new_n509), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n518), .A2(KEYINPUT32), .A3(new_n465), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT29), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n520), .B1(new_n506), .B2(new_n490), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n489), .B1(new_n484), .B2(new_n500), .ZN(new_n522));
  OAI21_X1  g336(.A(KEYINPUT74), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n503), .A2(new_n505), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n223), .B1(new_n480), .B2(new_n466), .ZN(new_n525));
  OAI21_X1  g339(.A(KEYINPUT28), .B1(new_n485), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(KEYINPUT75), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n480), .A2(new_n466), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(new_n475), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(new_n500), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT75), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n530), .A2(new_n531), .A3(KEYINPUT28), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n524), .B1(new_n527), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n490), .A2(new_n520), .ZN(new_n534));
  AOI21_X1  g348(.A(G902), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n523), .A2(new_n535), .ZN(new_n536));
  NOR3_X1   g350(.A1(new_n521), .A2(new_n522), .A3(KEYINPUT74), .ZN(new_n537));
  OAI21_X1  g351(.A(G472), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n516), .A2(new_n519), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n204), .A2(new_n247), .ZN(new_n540));
  OAI211_X1 g354(.A(KEYINPUT23), .B(new_n540), .C1(new_n209), .C2(new_n247), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT23), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n542), .B1(new_n209), .B2(G128), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n540), .B1(new_n209), .B2(new_n247), .ZN(new_n545));
  XOR2_X1   g359(.A(KEYINPUT24), .B(G110), .Z(new_n546));
  OAI22_X1  g360(.A1(new_n544), .A2(G110), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n403), .A2(G146), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n392), .A2(new_n241), .ZN(new_n549));
  AND3_X1   g363(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n544), .A2(G110), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n545), .A2(new_n546), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n551), .B(new_n552), .C1(new_n359), .C2(new_n363), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(KEYINPUT77), .ZN(new_n554));
  AOI22_X1  g368(.A1(new_n548), .A2(new_n358), .B1(new_n545), .B2(new_n546), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT77), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n555), .A2(new_n556), .A3(new_n551), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n550), .B1(new_n554), .B2(new_n557), .ZN(new_n558));
  XNOR2_X1  g372(.A(KEYINPUT22), .B(G137), .ZN(new_n559));
  AND3_X1   g373(.A1(new_n255), .A2(G221), .A3(G234), .ZN(new_n560));
  XOR2_X1   g374(.A(new_n559), .B(new_n560), .Z(new_n561));
  OAI21_X1  g375(.A(KEYINPUT78), .B1(new_n558), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n553), .A2(KEYINPUT77), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n556), .B1(new_n555), .B2(new_n551), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n563), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT78), .ZN(new_n567));
  INV_X1    g381(.A(new_n561), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n563), .B(new_n561), .C1(new_n564), .C2(new_n565), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT79), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n558), .A2(KEYINPUT79), .A3(new_n561), .ZN(new_n573));
  AOI22_X1  g387(.A1(new_n562), .A2(new_n569), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n453), .B1(G234), .B2(new_n286), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n575), .A2(G902), .ZN(new_n576));
  AOI21_X1  g390(.A(KEYINPUT80), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n562), .A2(new_n569), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n572), .A2(new_n573), .ZN(new_n579));
  AND4_X1   g393(.A1(KEYINPUT80), .A2(new_n578), .A3(new_n579), .A4(new_n576), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n578), .A2(new_n579), .A3(new_n286), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(KEYINPUT25), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT25), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n574), .A2(new_n584), .A3(new_n286), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n583), .A2(new_n585), .A3(new_n575), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n581), .A2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  AND3_X1   g402(.A1(new_n464), .A2(new_n539), .A3(new_n588), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n589), .B(new_n192), .ZN(G3));
  OAI21_X1  g404(.A(new_n286), .B1(new_n497), .B2(new_n513), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT94), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n591), .A2(new_n592), .A3(G472), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(G472), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n518), .A2(new_n286), .A3(new_n594), .ZN(new_n595));
  AND2_X1   g409(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n587), .B1(new_n349), .B2(new_n347), .ZN(new_n597));
  AND2_X1   g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AND2_X1   g412(.A1(new_n258), .A2(new_n273), .ZN(new_n599));
  OR2_X1    g413(.A1(new_n599), .A2(new_n274), .ZN(new_n600));
  INV_X1    g414(.A(new_n275), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n282), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(new_n434), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n458), .A2(new_n459), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n459), .A2(new_n286), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n445), .A2(new_n452), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT95), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(KEYINPUT33), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n610), .B1(new_n455), .B2(new_n456), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n457), .A2(KEYINPUT33), .A3(new_n609), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  OAI211_X1 g428(.A(new_n604), .B(new_n606), .C1(new_n614), .C2(new_n459), .ZN(new_n615));
  AND3_X1   g429(.A1(new_n398), .A2(new_n408), .A3(KEYINPUT91), .ZN(new_n616));
  AOI21_X1  g430(.A(KEYINPUT91), .B1(new_n398), .B2(new_n408), .ZN(new_n617));
  NOR3_X1   g431(.A1(new_n616), .A2(new_n617), .A3(new_n416), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT20), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n418), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n425), .A2(new_n422), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n615), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  OR2_X1    g436(.A1(new_n622), .A2(KEYINPUT96), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(KEYINPUT96), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n603), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n598), .A2(new_n625), .ZN(new_n626));
  XOR2_X1   g440(.A(KEYINPUT34), .B(G104), .Z(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G6));
  INV_X1    g442(.A(new_n415), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n414), .A2(KEYINPUT20), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n433), .B(KEYINPUT97), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n424), .A2(KEYINPUT92), .ZN(new_n634));
  AND3_X1   g448(.A1(new_n634), .A2(G475), .A3(new_n422), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n635), .A2(new_n461), .ZN(new_n636));
  AND4_X1   g450(.A1(new_n602), .A2(new_n632), .A3(new_n633), .A4(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n598), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT35), .B(G107), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G9));
  NOR2_X1   g454(.A1(new_n568), .A2(KEYINPUT36), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n558), .B(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n576), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n575), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n645), .B1(new_n582), .B2(KEYINPUT25), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n644), .B1(new_n646), .B2(new_n585), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n647), .A2(new_n462), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n593), .A2(new_n350), .A3(new_n595), .A4(new_n648), .ZN(new_n649));
  XOR2_X1   g463(.A(KEYINPUT37), .B(G110), .Z(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G12));
  AOI21_X1  g465(.A(new_n647), .B1(new_n349), .B2(new_n347), .ZN(new_n652));
  INV_X1    g466(.A(G900), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n428), .B1(new_n431), .B2(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(KEYINPUT98), .ZN(new_n655));
  NOR4_X1   g469(.A1(new_n631), .A2(new_n635), .A3(new_n461), .A4(new_n655), .ZN(new_n656));
  AND2_X1   g470(.A1(new_n656), .A2(new_n602), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n539), .A2(new_n652), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(G128), .ZN(G30));
  AOI21_X1  g473(.A(new_n490), .B1(new_n484), .B2(new_n500), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n286), .B1(new_n530), .B2(new_n489), .ZN(new_n661));
  OAI21_X1  g475(.A(G472), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n516), .A2(new_n519), .A3(new_n662), .ZN(new_n663));
  XOR2_X1   g477(.A(new_n663), .B(KEYINPUT99), .Z(new_n664));
  NAND2_X1  g478(.A1(new_n347), .A2(new_n349), .ZN(new_n665));
  XOR2_X1   g479(.A(new_n655), .B(KEYINPUT39), .Z(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  AND2_X1   g481(.A1(new_n667), .A2(KEYINPUT40), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n279), .B(KEYINPUT38), .ZN(new_n669));
  NOR4_X1   g483(.A1(new_n669), .A2(new_n426), .A3(new_n461), .A4(new_n282), .ZN(new_n670));
  OAI211_X1 g484(.A(new_n670), .B(new_n647), .C1(KEYINPUT40), .C2(new_n667), .ZN(new_n671));
  NOR3_X1   g485(.A1(new_n664), .A2(new_n668), .A3(new_n671), .ZN(new_n672));
  XOR2_X1   g486(.A(new_n672), .B(KEYINPUT100), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G143), .ZN(G45));
  NAND2_X1  g488(.A1(new_n604), .A2(new_n606), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n675), .B1(new_n613), .B2(G478), .ZN(new_n676));
  INV_X1    g490(.A(new_n655), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n417), .B1(new_n414), .B2(KEYINPUT20), .ZN(new_n678));
  OAI211_X1 g492(.A(new_n676), .B(new_n677), .C1(new_n635), .C2(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT101), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n620), .A2(new_n621), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n682), .A2(KEYINPUT101), .A3(new_n676), .A4(new_n677), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n681), .A2(new_n602), .A3(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT102), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n681), .A2(new_n683), .A3(KEYINPUT102), .A4(new_n602), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n539), .A2(new_n686), .A3(new_n652), .A4(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G146), .ZN(G48));
  INV_X1    g503(.A(new_n345), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n286), .B1(new_n326), .B2(new_n335), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(G469), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT103), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n692), .A2(new_n693), .A3(new_n336), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n691), .A2(KEYINPUT103), .A3(G469), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n690), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n539), .A2(new_n625), .A3(new_n588), .A4(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(KEYINPUT104), .ZN(new_n698));
  XNOR2_X1  g512(.A(KEYINPUT41), .B(G113), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(G15));
  NAND4_X1  g514(.A1(new_n539), .A2(new_n588), .A3(new_n637), .A4(new_n696), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G116), .ZN(G18));
  INV_X1    g516(.A(new_n644), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n586), .A2(new_n703), .ZN(new_n704));
  AND4_X1   g518(.A1(new_n463), .A2(new_n704), .A3(new_n602), .A4(new_n696), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n539), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G119), .ZN(G21));
  INV_X1    g521(.A(KEYINPUT106), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n708), .B1(new_n426), .B2(new_n461), .ZN(new_n709));
  INV_X1    g523(.A(new_n461), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n682), .A2(KEYINPUT106), .A3(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n709), .A2(new_n711), .A3(new_n602), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n696), .A2(new_n633), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT105), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n527), .A2(new_n532), .ZN(new_n716));
  INV_X1    g530(.A(new_n524), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n489), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT31), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n719), .B1(new_n484), .B2(new_n491), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n715), .B1(new_n718), .B2(new_n720), .ZN(new_n721));
  OAI211_X1 g535(.A(new_n511), .B(KEYINPUT105), .C1(new_n533), .C2(new_n489), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n721), .A2(new_n517), .A3(new_n722), .ZN(new_n723));
  AOI22_X1  g537(.A1(G472), .A2(new_n591), .B1(new_n723), .B2(new_n465), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n714), .A2(new_n724), .A3(new_n588), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G122), .ZN(G24));
  AND4_X1   g540(.A1(new_n602), .A2(new_n681), .A3(new_n683), .A4(new_n696), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n727), .A2(new_n724), .A3(new_n704), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G125), .ZN(G27));
  INV_X1    g543(.A(KEYINPUT108), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n514), .A2(new_n515), .ZN(new_n731));
  AOI21_X1  g545(.A(KEYINPUT32), .B1(new_n518), .B2(new_n465), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n730), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n516), .A2(new_n519), .A3(KEYINPUT108), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n733), .A2(new_n538), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n681), .A2(new_n683), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n280), .A2(new_n282), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT107), .ZN(new_n738));
  OR2_X1    g552(.A1(new_n343), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n690), .B1(new_n343), .B2(new_n738), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n737), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT42), .ZN(new_n742));
  NOR3_X1   g556(.A1(new_n736), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n735), .A2(new_n588), .A3(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(new_n736), .ZN(new_n745));
  INV_X1    g559(.A(new_n741), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n539), .A2(new_n588), .A3(new_n745), .A4(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(new_n742), .ZN(new_n748));
  AND2_X1   g562(.A1(new_n744), .A2(new_n748), .ZN(new_n749));
  XOR2_X1   g563(.A(KEYINPUT109), .B(G131), .Z(new_n750));
  XNOR2_X1  g564(.A(new_n749), .B(new_n750), .ZN(G33));
  NAND4_X1  g565(.A1(new_n539), .A2(new_n588), .A3(new_n656), .A4(new_n746), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G134), .ZN(G36));
  NAND2_X1  g567(.A1(new_n426), .A2(new_n676), .ZN(new_n754));
  XOR2_X1   g568(.A(new_n754), .B(KEYINPUT43), .Z(new_n755));
  INV_X1    g569(.A(new_n755), .ZN(new_n756));
  NOR3_X1   g570(.A1(new_n596), .A2(new_n647), .A3(new_n756), .ZN(new_n757));
  OR2_X1    g571(.A1(new_n757), .A2(KEYINPUT44), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(KEYINPUT44), .ZN(new_n759));
  INV_X1    g573(.A(new_n336), .ZN(new_n760));
  AND3_X1   g574(.A1(new_n340), .A2(new_n341), .A3(KEYINPUT45), .ZN(new_n761));
  AOI21_X1  g575(.A(KEYINPUT45), .B1(new_n340), .B2(new_n341), .ZN(new_n762));
  NOR3_X1   g576(.A1(new_n761), .A2(new_n762), .A3(new_n285), .ZN(new_n763));
  OR2_X1    g577(.A1(new_n763), .A2(new_n337), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT46), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n760), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n766), .B1(new_n765), .B2(new_n764), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n767), .A2(new_n345), .A3(new_n666), .ZN(new_n768));
  INV_X1    g582(.A(new_n737), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n758), .A2(new_n759), .A3(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G137), .ZN(G39));
  NAND2_X1  g586(.A1(new_n767), .A2(new_n345), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n773), .B1(KEYINPUT110), .B2(KEYINPUT47), .ZN(new_n774));
  AND2_X1   g588(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n775));
  NOR2_X1   g589(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n776));
  OAI211_X1 g590(.A(new_n767), .B(new_n345), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  NOR4_X1   g591(.A1(new_n539), .A2(new_n588), .A3(new_n736), .A4(new_n769), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n774), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G140), .ZN(G42));
  NAND2_X1  g594(.A1(new_n694), .A2(new_n695), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(KEYINPUT112), .ZN(new_n782));
  AOI22_X1  g596(.A1(new_n774), .A2(new_n777), .B1(new_n690), .B2(new_n782), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n755), .A2(new_n724), .A3(new_n588), .A4(new_n428), .ZN(new_n784));
  OR2_X1    g598(.A1(new_n784), .A2(new_n769), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n724), .A2(new_n704), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT115), .ZN(new_n787));
  INV_X1    g601(.A(new_n696), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n787), .B1(new_n788), .B2(new_n769), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n696), .A2(KEYINPUT115), .A3(new_n737), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n789), .A2(new_n428), .A3(new_n790), .ZN(new_n791));
  OR2_X1    g605(.A1(new_n791), .A2(new_n756), .ZN(new_n792));
  OAI22_X1  g606(.A1(new_n783), .A2(new_n785), .B1(new_n786), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n669), .A2(new_n282), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n784), .A2(new_n788), .A3(new_n794), .ZN(new_n795));
  OR2_X1    g609(.A1(new_n795), .A2(KEYINPUT50), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(KEYINPUT50), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n793), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n791), .A2(new_n587), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n664), .A2(new_n426), .A3(new_n615), .A4(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(KEYINPUT116), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n798), .A2(KEYINPUT51), .A3(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n784), .A2(new_n788), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(new_n602), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(KEYINPUT118), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n623), .A2(new_n624), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n664), .A2(new_n806), .A3(new_n799), .ZN(new_n807));
  AND4_X1   g621(.A1(G952), .A2(new_n805), .A3(new_n255), .A4(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(new_n792), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n735), .A2(new_n588), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(KEYINPUT48), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n802), .A2(new_n808), .A3(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT51), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n796), .A2(new_n797), .ZN(new_n815));
  OAI221_X1 g629(.A(new_n815), .B1(new_n786), .B2(new_n792), .C1(new_n783), .C2(new_n785), .ZN(new_n816));
  XOR2_X1   g630(.A(new_n800), .B(KEYINPUT116), .Z(new_n817));
  OAI21_X1  g631(.A(new_n814), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(KEYINPUT117), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT117), .ZN(new_n820));
  OAI211_X1 g634(.A(new_n820), .B(new_n814), .C1(new_n816), .C2(new_n817), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n813), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT114), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT53), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n621), .A2(new_n461), .A3(new_n677), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n769), .A2(new_n825), .A3(new_n631), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n539), .A2(new_n652), .A3(new_n826), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n724), .A2(new_n704), .A3(new_n745), .A4(new_n746), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n752), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n829), .B1(new_n744), .B2(new_n748), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n676), .B1(new_n635), .B2(new_n678), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n283), .B(new_n633), .C1(new_n275), .C2(new_n278), .ZN(new_n832));
  OAI21_X1  g646(.A(KEYINPUT113), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(new_n832), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT113), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n622), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n834), .A2(new_n426), .A3(new_n710), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n833), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n597), .A2(new_n838), .A3(new_n595), .A4(new_n593), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n725), .A2(new_n706), .A3(new_n839), .A4(new_n649), .ZN(new_n840));
  AND4_X1   g654(.A1(new_n539), .A2(new_n588), .A3(new_n637), .A4(new_n696), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n840), .A2(new_n589), .A3(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n830), .A2(new_n842), .A3(new_n698), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n647), .A2(new_n677), .A3(new_n739), .A4(new_n740), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n844), .A2(new_n712), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n663), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n688), .A2(new_n658), .A3(new_n728), .A4(new_n846), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(KEYINPUT52), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n824), .B1(new_n843), .B2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(new_n589), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n725), .A2(new_n839), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n706), .A2(new_n649), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n850), .A2(new_n851), .A3(new_n852), .A4(new_n701), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT104), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n697), .B(new_n854), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n658), .A2(new_n728), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n857), .A2(KEYINPUT52), .A3(new_n688), .A4(new_n846), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT52), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n847), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n856), .A2(new_n861), .A3(KEYINPUT53), .A4(new_n830), .ZN(new_n862));
  AND3_X1   g676(.A1(new_n849), .A2(KEYINPUT54), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(KEYINPUT54), .B1(new_n849), .B2(new_n862), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n823), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n849), .A2(new_n862), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT54), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n849), .A2(KEYINPUT54), .A3(new_n862), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n868), .A2(KEYINPUT114), .A3(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n822), .A2(new_n865), .A3(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n871), .B1(G952), .B2(G953), .ZN(new_n872));
  INV_X1    g686(.A(new_n669), .ZN(new_n873));
  NOR4_X1   g687(.A1(new_n587), .A2(new_n690), .A3(new_n754), .A4(new_n282), .ZN(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n873), .B1(new_n875), .B2(KEYINPUT111), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n782), .B(KEYINPUT49), .ZN(new_n877));
  OR2_X1    g691(.A1(new_n875), .A2(KEYINPUT111), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n664), .A2(new_n876), .A3(new_n877), .A4(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n872), .A2(new_n879), .ZN(G75));
  NOR2_X1   g694(.A1(new_n255), .A2(G952), .ZN(new_n881));
  INV_X1    g695(.A(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n286), .B1(new_n849), .B2(new_n862), .ZN(new_n883));
  AOI21_X1  g697(.A(KEYINPUT56), .B1(new_n883), .B2(G210), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n235), .A2(new_n237), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n885), .B(new_n257), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(KEYINPUT55), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n882), .B1(new_n884), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n883), .A2(new_n276), .ZN(new_n889));
  XOR2_X1   g703(.A(new_n889), .B(KEYINPUT119), .Z(new_n890));
  INV_X1    g704(.A(KEYINPUT56), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n887), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n888), .B1(new_n890), .B2(new_n892), .ZN(G51));
  NOR2_X1   g707(.A1(new_n863), .A2(new_n864), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n337), .B(KEYINPUT57), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n896), .B1(new_n326), .B2(new_n335), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n883), .A2(new_n763), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n881), .B1(new_n897), .B2(new_n898), .ZN(G54));
  NAND3_X1  g713(.A1(new_n883), .A2(KEYINPUT58), .A3(G475), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n616), .A2(new_n617), .ZN(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  OR2_X1    g716(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT120), .ZN(new_n904));
  OR2_X1    g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n903), .A2(new_n904), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n881), .B1(new_n900), .B2(new_n902), .ZN(new_n907));
  AND3_X1   g721(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(G60));
  NAND2_X1  g722(.A1(new_n865), .A2(new_n870), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n605), .B(KEYINPUT59), .ZN(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n614), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n613), .A2(new_n910), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n881), .B1(new_n894), .B2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(KEYINPUT121), .B1(new_n912), .B2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT121), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n910), .B1(new_n865), .B2(new_n870), .ZN(new_n918));
  OAI211_X1 g732(.A(new_n914), .B(new_n917), .C1(new_n918), .C2(new_n614), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n916), .A2(new_n919), .ZN(G63));
  NAND2_X1  g734(.A1(G217), .A2(G902), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT122), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT60), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n866), .A2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(new_n574), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n881), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n926), .B1(new_n642), .B2(new_n924), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT61), .Z(G66));
  INV_X1    g742(.A(G224), .ZN(new_n929));
  OAI21_X1  g743(.A(G953), .B1(new_n432), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n930), .B1(new_n856), .B2(G953), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n885), .B1(G898), .B2(new_n255), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n931), .B(new_n932), .ZN(G69));
  NAND3_X1  g747(.A1(new_n688), .A2(new_n658), .A3(new_n728), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(KEYINPUT124), .Z(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(new_n771), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT126), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n779), .A2(new_n752), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n768), .A2(new_n712), .ZN(new_n939));
  AOI211_X1 g753(.A(new_n749), .B(new_n938), .C1(new_n810), .C2(new_n939), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n937), .A2(new_n255), .A3(new_n940), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n474), .A2(new_n481), .A3(new_n483), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n942), .B(KEYINPUT123), .Z(new_n943));
  NAND2_X1  g757(.A1(new_n400), .A2(new_n401), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n943), .B(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(G900), .A2(G953), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n941), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n622), .B1(new_n426), .B2(new_n710), .ZN(new_n948));
  NOR3_X1   g762(.A1(new_n667), .A2(new_n769), .A3(new_n948), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n949), .A2(new_n539), .A3(new_n588), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT125), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n771), .A2(new_n779), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n673), .A2(new_n935), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n952), .B1(new_n953), .B2(KEYINPUT62), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT62), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n673), .A2(new_n955), .A3(new_n935), .ZN(new_n956));
  AOI21_X1  g770(.A(G953), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n947), .B1(new_n957), .B2(new_n945), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n255), .B1(G227), .B2(G900), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(new_n959), .ZN(new_n961));
  OAI211_X1 g775(.A(new_n947), .B(new_n961), .C1(new_n957), .C2(new_n945), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n960), .A2(new_n962), .ZN(G72));
  NAND2_X1  g777(.A1(G472), .A2(G902), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(KEYINPUT63), .Z(new_n965));
  AND2_X1   g779(.A1(new_n522), .A2(KEYINPUT127), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n510), .B1(new_n522), .B2(KEYINPUT127), .ZN(new_n967));
  OAI211_X1 g781(.A(new_n866), .B(new_n965), .C1(new_n966), .C2(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n968), .A2(new_n882), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n484), .A2(new_n500), .A3(new_n490), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n937), .A2(new_n856), .A3(new_n940), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n970), .B1(new_n971), .B2(new_n965), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n954), .A2(new_n856), .A3(new_n956), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(new_n965), .ZN(new_n974));
  AOI211_X1 g788(.A(new_n969), .B(new_n972), .C1(new_n974), .C2(new_n660), .ZN(G57));
endmodule


