//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 1 0 1 0 1 0 1 0 0 1 0 1 0 1 0 1 0 1 1 1 1 1 1 0 1 1 0 0 0 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n643, new_n644, new_n645,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n805, new_n806,
    new_n807, new_n809, new_n810, new_n811, new_n812, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n862, new_n863, new_n864, new_n866, new_n867, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n877,
    new_n878, new_n879, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n888, new_n889, new_n890, new_n891, new_n892, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n924, new_n925;
  INV_X1    g000(.A(KEYINPUT30), .ZN(new_n202));
  INV_X1    g001(.A(G169gat), .ZN(new_n203));
  INV_X1    g002(.A(G176gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NOR2_X1   g004(.A1(G169gat), .A2(G176gat), .ZN(new_n206));
  AOI21_X1  g005(.A(new_n205), .B1(KEYINPUT23), .B2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n207), .B(KEYINPUT66), .ZN(new_n208));
  OR2_X1    g007(.A1(new_n206), .A2(KEYINPUT23), .ZN(new_n209));
  NAND3_X1  g008(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n210));
  OR2_X1    g009(.A1(new_n210), .A2(KEYINPUT67), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(KEYINPUT67), .ZN(new_n212));
  INV_X1    g011(.A(G183gat), .ZN(new_n213));
  INV_X1    g012(.A(G190gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT24), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n216), .B1(new_n213), .B2(new_n214), .ZN(new_n217));
  NAND4_X1  g016(.A1(new_n211), .A2(new_n212), .A3(new_n215), .A4(new_n217), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n208), .A2(new_n209), .A3(new_n218), .ZN(new_n219));
  OR2_X1    g018(.A1(new_n215), .A2(KEYINPUT65), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n215), .A2(KEYINPUT65), .ZN(new_n221));
  NAND4_X1  g020(.A1(new_n220), .A2(new_n217), .A3(new_n210), .A4(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT25), .ZN(new_n223));
  AND3_X1   g022(.A1(new_n222), .A2(new_n223), .A3(new_n207), .ZN(new_n224));
  AOI22_X1  g023(.A1(new_n219), .A2(KEYINPUT25), .B1(new_n209), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(KEYINPUT27), .B(G183gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(new_n214), .ZN(new_n227));
  XOR2_X1   g026(.A(new_n227), .B(KEYINPUT28), .Z(new_n228));
  INV_X1    g027(.A(KEYINPUT68), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n206), .A2(new_n229), .ZN(new_n230));
  OR2_X1    g029(.A1(new_n230), .A2(KEYINPUT26), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(KEYINPUT26), .ZN(new_n232));
  OAI211_X1 g031(.A(new_n231), .B(new_n232), .C1(new_n203), .C2(new_n204), .ZN(new_n233));
  OAI211_X1 g032(.A(new_n228), .B(new_n233), .C1(new_n213), .C2(new_n214), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n225), .A2(new_n234), .ZN(new_n235));
  AND3_X1   g034(.A1(new_n235), .A2(G226gat), .A3(G233gat), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT29), .ZN(new_n237));
  AOI22_X1  g036(.A1(new_n235), .A2(new_n237), .B1(G226gat), .B2(G233gat), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(G197gat), .B(G204gat), .ZN(new_n240));
  INV_X1    g039(.A(G211gat), .ZN(new_n241));
  INV_X1    g040(.A(G218gat), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n240), .B1(KEYINPUT22), .B2(new_n243), .ZN(new_n244));
  XOR2_X1   g043(.A(G211gat), .B(G218gat), .Z(new_n245));
  XNOR2_X1  g044(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n239), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(G8gat), .B(G36gat), .ZN(new_n248));
  INV_X1    g047(.A(G64gat), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n248), .B(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(G92gat), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n250), .B(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n202), .B1(new_n247), .B2(new_n252), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n247), .A2(new_n252), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n253), .B(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT40), .ZN(new_n256));
  INV_X1    g055(.A(G120gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(G113gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(KEYINPUT69), .B(G113gat), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n258), .B1(new_n259), .B2(new_n257), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT1), .ZN(new_n261));
  XNOR2_X1  g060(.A(G127gat), .B(G134gat), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n260), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n263), .B(KEYINPUT70), .ZN(new_n264));
  INV_X1    g063(.A(new_n262), .ZN(new_n265));
  XNOR2_X1  g064(.A(G113gat), .B(G120gat), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n265), .B1(KEYINPUT1), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n264), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(G155gat), .ZN(new_n269));
  INV_X1    g068(.A(G162gat), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n269), .A2(new_n270), .ZN(new_n273));
  XNOR2_X1  g072(.A(G141gat), .B(G148gat), .ZN(new_n274));
  XOR2_X1   g073(.A(new_n274), .B(KEYINPUT71), .Z(new_n275));
  XNOR2_X1  g074(.A(KEYINPUT72), .B(KEYINPUT2), .ZN(new_n276));
  OAI211_X1 g075(.A(new_n272), .B(new_n273), .C1(new_n275), .C2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n274), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n273), .A2(KEYINPUT2), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n278), .B1(new_n271), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n277), .A2(new_n280), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n268), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT4), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(KEYINPUT74), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n282), .A2(new_n283), .ZN(new_n286));
  OR2_X1    g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n281), .A2(KEYINPUT3), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT3), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n277), .A2(new_n289), .A3(new_n280), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n288), .A2(new_n268), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n285), .A2(new_n286), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n287), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(G225gat), .A2(G233gat), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  XOR2_X1   g095(.A(new_n268), .B(new_n281), .Z(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(new_n294), .ZN(new_n298));
  AND3_X1   g097(.A1(new_n296), .A2(KEYINPUT39), .A3(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(KEYINPUT0), .B(G57gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n300), .B(G85gat), .ZN(new_n301));
  XNOR2_X1  g100(.A(G1gat), .B(G29gat), .ZN(new_n302));
  XOR2_X1   g101(.A(new_n301), .B(new_n302), .Z(new_n303));
  OAI21_X1  g102(.A(new_n303), .B1(new_n296), .B2(KEYINPUT39), .ZN(new_n304));
  OAI211_X1 g103(.A(KEYINPUT78), .B(new_n256), .C1(new_n299), .C2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n291), .A2(new_n294), .ZN(new_n306));
  XNOR2_X1  g105(.A(KEYINPUT73), .B(KEYINPUT5), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n287), .A2(new_n292), .A3(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n282), .B(KEYINPUT4), .ZN(new_n310));
  OAI221_X1 g109(.A(new_n307), .B1(new_n297), .B2(new_n294), .C1(new_n310), .C2(new_n306), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n303), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  OR2_X1    g112(.A1(new_n296), .A2(KEYINPUT39), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n256), .A2(KEYINPUT78), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n296), .A2(KEYINPUT39), .A3(new_n298), .ZN(new_n316));
  NAND4_X1  g115(.A1(new_n314), .A2(new_n303), .A3(new_n315), .A4(new_n316), .ZN(new_n317));
  NAND4_X1  g116(.A1(new_n255), .A2(new_n305), .A3(new_n313), .A4(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n252), .ZN(new_n319));
  INV_X1    g118(.A(new_n246), .ZN(new_n320));
  XNOR2_X1  g119(.A(new_n239), .B(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT37), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n319), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n247), .A2(KEYINPUT37), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n254), .B1(new_n325), .B2(KEYINPUT38), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT6), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n309), .A2(new_n311), .A3(new_n303), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n313), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n312), .A2(KEYINPUT6), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT79), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n324), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT38), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n247), .A2(KEYINPUT79), .A3(KEYINPUT37), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n332), .A2(new_n333), .A3(new_n323), .A4(new_n334), .ZN(new_n335));
  NAND4_X1  g134(.A1(new_n326), .A2(new_n329), .A3(new_n330), .A4(new_n335), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n246), .B1(new_n290), .B2(new_n237), .ZN(new_n337));
  AOI21_X1  g136(.A(KEYINPUT3), .B1(new_n246), .B2(new_n237), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n338), .B1(new_n280), .B2(new_n277), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(G228gat), .A2(G233gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n341), .B(G22gat), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  XNOR2_X1  g142(.A(new_n340), .B(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT77), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(G78gat), .B(G106gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(KEYINPUT76), .B(KEYINPUT31), .ZN(new_n349));
  INV_X1    g148(.A(G50gat), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n349), .B(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n347), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n344), .A2(new_n345), .A3(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n348), .A2(new_n351), .A3(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n351), .B1(new_n348), .B2(new_n353), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n318), .A2(new_n336), .A3(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n235), .B(new_n268), .ZN(new_n360));
  NAND2_X1  g159(.A1(G227gat), .A2(G233gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n361), .B(KEYINPUT64), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT32), .ZN(new_n364));
  OR3_X1    g163(.A1(new_n360), .A2(KEYINPUT34), .A3(new_n362), .ZN(new_n365));
  OAI21_X1  g164(.A(KEYINPUT34), .B1(new_n360), .B2(new_n362), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n364), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  XNOR2_X1  g167(.A(G15gat), .B(G43gat), .ZN(new_n369));
  XNOR2_X1  g168(.A(G71gat), .B(G99gat), .ZN(new_n370));
  XOR2_X1   g169(.A(new_n369), .B(new_n370), .Z(new_n371));
  INV_X1    g170(.A(new_n363), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n371), .B1(new_n372), .B2(KEYINPUT33), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n365), .A2(new_n364), .A3(new_n366), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n368), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n375), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n373), .B1(new_n377), .B2(new_n367), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT36), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n376), .A2(new_n378), .A3(KEYINPUT36), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT75), .ZN(new_n384));
  OR2_X1    g183(.A1(new_n329), .A2(new_n384), .ZN(new_n385));
  AOI22_X1  g184(.A1(new_n329), .A2(new_n384), .B1(KEYINPUT6), .B2(new_n312), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n255), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n359), .B(new_n383), .C1(new_n387), .C2(new_n358), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n379), .A2(new_n357), .ZN(new_n389));
  INV_X1    g188(.A(new_n255), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n329), .A2(new_n330), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n389), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT35), .ZN(new_n393));
  NOR3_X1   g192(.A1(new_n379), .A2(new_n357), .A3(new_n393), .ZN(new_n394));
  AOI22_X1  g193(.A1(new_n392), .A2(new_n393), .B1(new_n387), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n388), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT91), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n249), .A2(G57gat), .ZN(new_n398));
  INV_X1    g197(.A(G57gat), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(G64gat), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(KEYINPUT90), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  AND2_X1   g203(.A1(G71gat), .A2(G78gat), .ZN(new_n405));
  NOR2_X1   g204(.A1(G71gat), .A2(G78gat), .ZN(new_n406));
  OAI22_X1  g205(.A1(new_n402), .A2(KEYINPUT90), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n397), .B1(new_n404), .B2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT90), .ZN(new_n409));
  NAND2_X1  g208(.A1(G71gat), .A2(G78gat), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT9), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  OR2_X1    g211(.A1(G71gat), .A2(G78gat), .ZN(new_n413));
  AOI22_X1  g212(.A1(new_n409), .A2(new_n412), .B1(new_n413), .B2(new_n410), .ZN(new_n414));
  AOI22_X1  g213(.A1(new_n398), .A2(new_n400), .B1(new_n402), .B2(KEYINPUT90), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n414), .A2(new_n415), .A3(KEYINPUT91), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n405), .A2(new_n406), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n401), .A2(KEYINPUT9), .ZN(new_n418));
  AOI22_X1  g217(.A1(new_n408), .A2(new_n416), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n419), .A2(KEYINPUT21), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  OR2_X1    g220(.A1(G15gat), .A2(G22gat), .ZN(new_n422));
  INV_X1    g221(.A(G1gat), .ZN(new_n423));
  NAND2_X1  g222(.A1(G15gat), .A2(G22gat), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n422), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(KEYINPUT85), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT83), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT16), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n427), .B1(new_n428), .B2(G1gat), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n423), .A2(KEYINPUT83), .A3(KEYINPUT16), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n422), .A2(new_n424), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT84), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n426), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  AOI22_X1  g234(.A1(new_n429), .A2(new_n430), .B1(new_n422), .B2(new_n424), .ZN(new_n436));
  INV_X1    g235(.A(G8gat), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n434), .A2(new_n437), .ZN(new_n438));
  OAI22_X1  g237(.A1(new_n436), .A2(new_n438), .B1(KEYINPUT85), .B2(new_n425), .ZN(new_n439));
  OAI21_X1  g238(.A(G8gat), .B1(new_n435), .B2(new_n439), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n433), .B(new_n425), .C1(new_n434), .C2(new_n437), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n419), .A2(KEYINPUT21), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(G183gat), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT92), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n443), .A2(new_n213), .A3(new_n444), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n447), .B1(new_n446), .B2(new_n448), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n421), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n451), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n453), .A2(new_n449), .A3(new_n420), .ZN(new_n454));
  XNOR2_X1  g253(.A(G127gat), .B(G155gat), .ZN(new_n455));
  XNOR2_X1  g254(.A(new_n455), .B(G211gat), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  AND3_X1   g256(.A1(new_n452), .A2(new_n454), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n457), .B1(new_n452), .B2(new_n454), .ZN(new_n459));
  XOR2_X1   g258(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n460));
  NAND2_X1  g259(.A1(G231gat), .A2(G233gat), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n460), .B(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  OR3_X1    g262(.A1(new_n458), .A2(new_n459), .A3(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n463), .B1(new_n458), .B2(new_n459), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(G232gat), .A2(G233gat), .ZN(new_n468));
  XNOR2_X1  g267(.A(new_n468), .B(KEYINPUT93), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(KEYINPUT41), .ZN(new_n470));
  INV_X1    g269(.A(G29gat), .ZN(new_n471));
  INV_X1    g270(.A(G36gat), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT14), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n475), .A2(new_n471), .A3(new_n472), .A4(KEYINPUT80), .ZN(new_n476));
  OAI21_X1  g275(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g277(.A1(G29gat), .A2(G36gat), .ZN(new_n479));
  AOI21_X1  g278(.A(KEYINPUT80), .B1(new_n479), .B2(new_n475), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n474), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(G43gat), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n482), .A2(G50gat), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n350), .A2(G43gat), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT15), .ZN(new_n485));
  NOR3_X1   g284(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n481), .A2(new_n486), .ZN(new_n487));
  XNOR2_X1  g286(.A(G43gat), .B(G50gat), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n473), .B1(new_n488), .B2(KEYINPUT15), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n485), .B1(new_n483), .B2(new_n484), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT81), .ZN(new_n491));
  INV_X1    g290(.A(new_n477), .ZN(new_n492));
  NOR3_X1   g291(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n479), .A2(new_n475), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n495), .A2(KEYINPUT81), .A3(new_n477), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n489), .A2(new_n490), .A3(new_n494), .A4(new_n496), .ZN(new_n497));
  AND2_X1   g296(.A1(new_n487), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(G99gat), .A2(G106gat), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT96), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(KEYINPUT96), .A2(G99gat), .A3(G106gat), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n501), .A2(KEYINPUT8), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(KEYINPUT94), .A2(KEYINPUT7), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT95), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n505), .A2(new_n506), .A3(G85gat), .A4(G92gat), .ZN(new_n507));
  OR2_X1    g306(.A1(new_n506), .A2(KEYINPUT7), .ZN(new_n508));
  NOR2_X1   g307(.A1(G85gat), .A2(G92gat), .ZN(new_n509));
  NAND2_X1  g308(.A1(G85gat), .A2(G92gat), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n509), .B1(new_n504), .B2(new_n510), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n503), .A2(new_n507), .A3(new_n508), .A4(new_n511), .ZN(new_n512));
  XOR2_X1   g311(.A(G99gat), .B(G106gat), .Z(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n504), .A2(new_n510), .ZN(new_n515));
  INV_X1    g314(.A(new_n509), .ZN(new_n516));
  AND3_X1   g315(.A1(new_n508), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n513), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n517), .A2(new_n518), .A3(new_n503), .A4(new_n507), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n514), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n470), .B1(new_n498), .B2(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n521), .B(KEYINPUT97), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n487), .A2(KEYINPUT17), .A3(new_n497), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n487), .A2(new_n497), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT17), .ZN(new_n525));
  AOI21_X1  g324(.A(KEYINPUT82), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT82), .ZN(new_n527));
  AOI211_X1 g326(.A(new_n527), .B(KEYINPUT17), .C1(new_n487), .C2(new_n497), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n520), .B(new_n523), .C1(new_n526), .C2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n522), .A2(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(G134gat), .B(G162gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n469), .A2(KEYINPUT41), .ZN(new_n533));
  XNOR2_X1  g332(.A(G190gat), .B(G218gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n533), .B(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n531), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n522), .A2(new_n536), .A3(new_n529), .ZN(new_n537));
  AND3_X1   g336(.A1(new_n532), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n535), .B1(new_n532), .B2(new_n537), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n467), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n418), .A2(new_n417), .ZN(new_n543));
  NOR3_X1   g342(.A1(new_n404), .A2(new_n407), .A3(new_n397), .ZN(new_n544));
  AOI21_X1  g343(.A(KEYINPUT91), .B1(new_n414), .B2(new_n415), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(new_n520), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n408), .A2(new_n416), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n548), .A2(new_n543), .A3(new_n514), .A4(new_n519), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT10), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n547), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n419), .A2(KEYINPUT10), .A3(new_n519), .A4(new_n514), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(G230gat), .A2(G233gat), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n554), .B1(new_n547), .B2(new_n549), .ZN(new_n556));
  OR2_X1    g355(.A1(new_n556), .A2(KEYINPUT98), .ZN(new_n557));
  XNOR2_X1  g356(.A(G120gat), .B(G148gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(G204gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n559), .B(KEYINPUT99), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n560), .B(new_n204), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n547), .A2(new_n549), .ZN(new_n563));
  INV_X1    g362(.A(new_n554), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n563), .A2(KEYINPUT98), .A3(new_n564), .ZN(new_n565));
  NAND4_X1  g364(.A1(new_n555), .A2(new_n557), .A3(new_n562), .A4(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(KEYINPUT101), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n557), .A2(new_n565), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT100), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n569), .B1(new_n553), .B2(new_n554), .ZN(new_n570));
  AOI211_X1 g369(.A(KEYINPUT100), .B(new_n564), .C1(new_n551), .C2(new_n552), .ZN(new_n571));
  NOR3_X1   g370(.A1(new_n568), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n567), .B1(new_n572), .B2(new_n562), .ZN(new_n573));
  OR2_X1    g372(.A1(new_n570), .A2(new_n571), .ZN(new_n574));
  OAI211_X1 g373(.A(KEYINPUT101), .B(new_n561), .C1(new_n574), .C2(new_n568), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(KEYINPUT11), .B(G169gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(G197gat), .ZN(new_n579));
  XOR2_X1   g378(.A(G113gat), .B(G141gat), .Z(new_n580));
  XOR2_X1   g379(.A(new_n579), .B(new_n580), .Z(new_n581));
  XOR2_X1   g380(.A(new_n581), .B(KEYINPUT12), .Z(new_n582));
  NOR2_X1   g381(.A1(new_n526), .A2(new_n528), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n440), .A2(new_n523), .A3(new_n441), .ZN(new_n584));
  OAI21_X1  g383(.A(KEYINPUT86), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  AND3_X1   g384(.A1(new_n440), .A2(new_n523), .A3(new_n441), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT86), .ZN(new_n587));
  OAI211_X1 g386(.A(new_n586), .B(new_n587), .C1(new_n526), .C2(new_n528), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n442), .A2(new_n524), .ZN(new_n590));
  NAND2_X1  g389(.A1(G229gat), .A2(G233gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(KEYINPUT18), .B1(new_n589), .B2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT18), .ZN(new_n595));
  AOI211_X1 g394(.A(new_n595), .B(new_n592), .C1(new_n585), .C2(new_n588), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT88), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n498), .A2(new_n440), .A3(new_n441), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n590), .A2(new_n599), .ZN(new_n600));
  XOR2_X1   g399(.A(new_n591), .B(KEYINPUT87), .Z(new_n601));
  XOR2_X1   g400(.A(new_n601), .B(KEYINPUT13), .Z(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n598), .B1(new_n600), .B2(new_n603), .ZN(new_n604));
  AOI211_X1 g403(.A(KEYINPUT88), .B(new_n602), .C1(new_n590), .C2(new_n599), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n582), .B1(new_n597), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n589), .A2(new_n593), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n609), .A2(new_n595), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n589), .A2(KEYINPUT18), .A3(new_n593), .ZN(new_n611));
  NAND4_X1  g410(.A1(new_n610), .A2(new_n582), .A3(new_n611), .A4(new_n607), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT89), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND4_X1  g413(.A1(new_n597), .A2(KEYINPUT89), .A3(new_n582), .A4(new_n607), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n608), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND4_X1  g416(.A1(new_n396), .A2(new_n542), .A3(new_n577), .A4(new_n617), .ZN(new_n618));
  OR2_X1    g417(.A1(new_n618), .A2(KEYINPUT102), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(KEYINPUT102), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n385), .A2(new_n386), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(G1gat), .ZN(G1324gat));
  AOI21_X1  g424(.A(new_n390), .B1(new_n619), .B2(new_n620), .ZN(new_n626));
  NAND2_X1  g425(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n428), .A2(new_n437), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT42), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  OR2_X1    g430(.A1(new_n626), .A2(new_n437), .ZN(new_n632));
  NAND4_X1  g431(.A1(new_n626), .A2(KEYINPUT42), .A3(new_n627), .A4(new_n628), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n631), .A2(new_n632), .A3(new_n633), .ZN(G1325gat));
  INV_X1    g433(.A(new_n379), .ZN(new_n635));
  AOI21_X1  g434(.A(G15gat), .B1(new_n621), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n383), .A2(KEYINPUT103), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT103), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n381), .A2(new_n638), .A3(new_n382), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n640), .B1(new_n619), .B2(new_n620), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n636), .B1(G15gat), .B2(new_n641), .ZN(G1326gat));
  NAND2_X1  g441(.A1(new_n621), .A2(new_n357), .ZN(new_n643));
  XOR2_X1   g442(.A(KEYINPUT43), .B(G22gat), .Z(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(KEYINPUT104), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n643), .B(new_n645), .ZN(G1327gat));
  INV_X1    g445(.A(new_n540), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n396), .A2(KEYINPUT44), .A3(new_n647), .ZN(new_n648));
  XOR2_X1   g447(.A(new_n576), .B(KEYINPUT105), .Z(new_n649));
  NAND3_X1  g448(.A1(new_n649), .A2(new_n466), .A3(new_n617), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(KEYINPUT106), .ZN(new_n651));
  OAI211_X1 g450(.A(new_n640), .B(new_n359), .C1(new_n387), .C2(new_n358), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n540), .B1(new_n652), .B2(new_n395), .ZN(new_n653));
  OAI211_X1 g452(.A(new_n648), .B(new_n651), .C1(new_n653), .C2(KEYINPUT44), .ZN(new_n654));
  OAI21_X1  g453(.A(G29gat), .B1(new_n654), .B2(new_n622), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT45), .ZN(new_n656));
  AOI211_X1 g455(.A(new_n576), .B(new_n616), .C1(new_n388), .C2(new_n395), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n657), .A2(new_n466), .A3(new_n647), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n658), .A2(new_n622), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n656), .B1(new_n659), .B2(new_n471), .ZN(new_n660));
  NOR4_X1   g459(.A1(new_n658), .A2(KEYINPUT45), .A3(G29gat), .A4(new_n622), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n655), .B1(new_n660), .B2(new_n661), .ZN(G1328gat));
  INV_X1    g461(.A(new_n658), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n663), .A2(new_n472), .A3(new_n255), .ZN(new_n664));
  AND2_X1   g463(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n665));
  NOR2_X1   g464(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n664), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  OAI21_X1  g466(.A(G36gat), .B1(new_n654), .B2(new_n390), .ZN(new_n668));
  OAI211_X1 g467(.A(new_n667), .B(new_n668), .C1(new_n665), .C2(new_n664), .ZN(G1329gat));
  OAI21_X1  g468(.A(KEYINPUT108), .B1(new_n654), .B2(new_n640), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n359), .B1(new_n387), .B2(new_n358), .ZN(new_n671));
  INV_X1    g470(.A(new_n639), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n638), .B1(new_n381), .B2(new_n382), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n395), .B1(new_n671), .B2(new_n674), .ZN(new_n675));
  AOI21_X1  g474(.A(KEYINPUT44), .B1(new_n675), .B2(new_n647), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT44), .ZN(new_n677));
  AOI211_X1 g476(.A(new_n677), .B(new_n540), .C1(new_n388), .C2(new_n395), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT108), .ZN(new_n680));
  NAND4_X1  g479(.A1(new_n679), .A2(new_n680), .A3(new_n674), .A4(new_n651), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n670), .A2(new_n681), .A3(G43gat), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n635), .A2(new_n482), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n658), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n682), .A2(KEYINPUT47), .A3(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT47), .ZN(new_n687));
  INV_X1    g486(.A(new_n654), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n482), .B1(new_n688), .B2(new_n674), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n687), .B1(new_n689), .B2(new_n684), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n686), .A2(new_n690), .ZN(G1330gat));
  OAI21_X1  g490(.A(G50gat), .B1(new_n654), .B2(new_n358), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n663), .A2(new_n350), .A3(new_n357), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT48), .ZN(new_n694));
  AND3_X1   g493(.A1(new_n692), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n694), .B1(new_n692), .B2(new_n693), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n695), .A2(new_n696), .ZN(G1331gat));
  NAND2_X1  g496(.A1(new_n542), .A2(new_n616), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n698), .B1(new_n652), .B2(new_n395), .ZN(new_n699));
  INV_X1    g498(.A(new_n649), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n622), .B(KEYINPUT109), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(new_n399), .ZN(G1332gat));
  NAND3_X1  g503(.A1(new_n699), .A2(new_n255), .A3(new_n700), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT49), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n706), .A2(new_n249), .ZN(new_n707));
  OR3_X1    g506(.A1(new_n705), .A2(KEYINPUT110), .A3(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(KEYINPUT110), .B1(new_n705), .B2(new_n707), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n710), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n711));
  NAND4_X1  g510(.A1(new_n708), .A2(new_n706), .A3(new_n709), .A4(new_n249), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(G1333gat));
  NAND4_X1  g512(.A1(new_n699), .A2(G71gat), .A3(new_n674), .A4(new_n700), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n701), .A2(new_n379), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n714), .B1(G71gat), .B2(new_n715), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g516(.A1(new_n701), .A2(new_n358), .ZN(new_n718));
  XOR2_X1   g517(.A(KEYINPUT111), .B(G78gat), .Z(new_n719));
  XNOR2_X1  g518(.A(new_n718), .B(new_n719), .ZN(G1335gat));
  NOR2_X1   g519(.A1(new_n467), .A2(new_n617), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n679), .A2(new_n576), .A3(new_n721), .ZN(new_n722));
  OAI21_X1  g521(.A(G85gat), .B1(new_n722), .B2(new_n622), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n653), .A2(KEYINPUT51), .A3(new_n721), .ZN(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n675), .A2(new_n647), .A3(new_n721), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT51), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n576), .B1(new_n725), .B2(new_n729), .ZN(new_n730));
  OR2_X1    g529(.A1(new_n622), .A2(G85gat), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n723), .B1(new_n730), .B2(new_n731), .ZN(G1336gat));
  INV_X1    g531(.A(new_n721), .ZN(new_n733));
  NOR4_X1   g532(.A1(new_n676), .A2(new_n678), .A3(new_n577), .A4(new_n733), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n251), .B1(new_n734), .B2(new_n255), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n390), .A2(G92gat), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  AOI211_X1 g536(.A(new_n649), .B(new_n737), .C1(new_n724), .C2(new_n728), .ZN(new_n738));
  OAI21_X1  g537(.A(KEYINPUT52), .B1(new_n735), .B2(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(G92gat), .B1(new_n722), .B2(new_n390), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT52), .ZN(new_n741));
  OAI211_X1 g540(.A(new_n700), .B(new_n736), .C1(new_n725), .C2(new_n729), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n740), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n739), .A2(new_n743), .ZN(G1337gat));
  OAI21_X1  g543(.A(G99gat), .B1(new_n722), .B2(new_n640), .ZN(new_n745));
  OR2_X1    g544(.A1(new_n379), .A2(G99gat), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n745), .B1(new_n730), .B2(new_n746), .ZN(G1338gat));
  INV_X1    g546(.A(G106gat), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n748), .B1(new_n734), .B2(new_n357), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n358), .A2(G106gat), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  AOI211_X1 g550(.A(new_n649), .B(new_n751), .C1(new_n724), .C2(new_n728), .ZN(new_n752));
  OAI21_X1  g551(.A(KEYINPUT53), .B1(new_n749), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(G106gat), .B1(new_n722), .B2(new_n358), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT53), .ZN(new_n755));
  OAI211_X1 g554(.A(new_n700), .B(new_n750), .C1(new_n725), .C2(new_n729), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n754), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n753), .A2(new_n757), .ZN(G1339gat));
  NAND2_X1  g557(.A1(new_n589), .A2(new_n590), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n759), .A2(G229gat), .A3(G233gat), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n600), .A2(new_n603), .ZN(new_n761));
  INV_X1    g560(.A(new_n761), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n581), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  NOR3_X1   g563(.A1(new_n594), .A2(new_n596), .A3(new_n606), .ZN(new_n765));
  AOI21_X1  g564(.A(KEYINPUT89), .B1(new_n765), .B2(new_n582), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n612), .A2(new_n613), .ZN(new_n767));
  OAI211_X1 g566(.A(new_n576), .B(new_n764), .C1(new_n766), .C2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(new_n566), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT54), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n770), .B1(new_n570), .B2(new_n571), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n551), .A2(new_n564), .A3(new_n552), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n555), .A2(KEYINPUT54), .A3(new_n772), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n771), .A2(new_n561), .A3(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT55), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n769), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n771), .A2(KEYINPUT55), .A3(new_n561), .A4(new_n773), .ZN(new_n777));
  AND2_X1   g576(.A1(new_n777), .A2(KEYINPUT112), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n777), .A2(KEYINPUT112), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n776), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n768), .B1(new_n616), .B2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT113), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  OAI211_X1 g582(.A(new_n768), .B(KEYINPUT113), .C1(new_n616), .C2(new_n780), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n783), .A2(new_n540), .A3(new_n784), .ZN(new_n785));
  AOI211_X1 g584(.A(new_n763), .B(new_n540), .C1(new_n614), .C2(new_n615), .ZN(new_n786));
  INV_X1    g585(.A(new_n780), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n785), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(new_n466), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n467), .A2(new_n540), .A3(new_n577), .A4(new_n616), .ZN(new_n791));
  AOI211_X1 g590(.A(new_n379), .B(new_n357), .C1(new_n790), .C2(new_n791), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n702), .A2(new_n255), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  OR3_X1    g593(.A1(new_n794), .A2(new_n259), .A3(new_n616), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n622), .A2(new_n255), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n792), .A2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(new_n617), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT114), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n799), .A2(new_n800), .A3(G113gat), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n800), .B1(new_n799), .B2(G113gat), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n795), .B1(new_n802), .B2(new_n803), .ZN(G1340gat));
  OAI21_X1  g603(.A(G120gat), .B1(new_n797), .B2(new_n649), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n576), .A2(new_n257), .ZN(new_n806));
  XOR2_X1   g605(.A(new_n806), .B(KEYINPUT115), .Z(new_n807));
  OAI21_X1  g606(.A(new_n805), .B1(new_n794), .B2(new_n807), .ZN(G1341gat));
  INV_X1    g607(.A(G127gat), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n797), .A2(new_n809), .A3(new_n466), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n794), .A2(new_n466), .ZN(new_n811));
  XOR2_X1   g610(.A(new_n811), .B(KEYINPUT116), .Z(new_n812));
  AOI21_X1  g611(.A(new_n810), .B1(new_n812), .B2(new_n809), .ZN(G1342gat));
  NAND2_X1  g612(.A1(new_n798), .A2(new_n647), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT117), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n814), .A2(new_n815), .A3(G134gat), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n815), .B1(new_n814), .B2(G134gat), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n794), .A2(G134gat), .ZN(new_n819));
  AOI21_X1  g618(.A(KEYINPUT56), .B1(new_n819), .B2(new_n647), .ZN(new_n820));
  AND3_X1   g619(.A1(new_n819), .A2(KEYINPUT56), .A3(new_n647), .ZN(new_n821));
  OAI22_X1  g620(.A1(new_n817), .A2(new_n818), .B1(new_n820), .B2(new_n821), .ZN(G1343gat));
  NOR2_X1   g621(.A1(new_n616), .A2(new_n780), .ZN(new_n823));
  AOI221_X4 g622(.A(new_n763), .B1(new_n573), .B2(new_n575), .C1(new_n614), .C2(new_n615), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n540), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n467), .B1(new_n825), .B2(new_n788), .ZN(new_n826));
  NOR4_X1   g625(.A1(new_n466), .A2(new_n617), .A3(new_n647), .A4(new_n576), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n357), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT57), .ZN(new_n829));
  OR3_X1    g628(.A1(new_n828), .A2(KEYINPUT118), .A3(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(KEYINPUT118), .B1(new_n828), .B2(new_n829), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n358), .B1(new_n790), .B2(new_n791), .ZN(new_n832));
  OAI211_X1 g631(.A(new_n830), .B(new_n831), .C1(new_n832), .C2(KEYINPUT57), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n640), .A2(new_n796), .ZN(new_n834));
  INV_X1    g633(.A(new_n834), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n833), .A2(G141gat), .A3(new_n617), .A4(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT58), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(KEYINPUT119), .ZN(new_n838));
  INV_X1    g637(.A(G141gat), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n832), .A2(new_n640), .A3(new_n793), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n839), .B1(new_n840), .B2(new_n616), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n836), .A2(new_n838), .A3(new_n841), .ZN(new_n842));
  OR2_X1    g641(.A1(new_n837), .A2(KEYINPUT119), .ZN(new_n843));
  XNOR2_X1  g642(.A(new_n842), .B(new_n843), .ZN(G1344gat));
  NAND2_X1  g643(.A1(new_n832), .A2(new_n640), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n845), .A2(new_n255), .A3(new_n702), .ZN(new_n846));
  INV_X1    g645(.A(G148gat), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n846), .A2(new_n847), .A3(new_n576), .ZN(new_n848));
  NAND2_X1  g647(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n467), .B1(new_n785), .B2(new_n788), .ZN(new_n850));
  OAI211_X1 g649(.A(KEYINPUT57), .B(new_n357), .C1(new_n850), .C2(new_n827), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT120), .ZN(new_n852));
  AOI22_X1  g651(.A1(new_n781), .A2(new_n540), .B1(new_n787), .B2(new_n786), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n791), .B1(new_n853), .B2(new_n467), .ZN(new_n854));
  AOI211_X1 g653(.A(new_n852), .B(KEYINPUT57), .C1(new_n854), .C2(new_n357), .ZN(new_n855));
  AOI21_X1  g654(.A(KEYINPUT120), .B1(new_n828), .B2(new_n829), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n851), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  AND3_X1   g656(.A1(new_n857), .A2(new_n576), .A3(new_n835), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n833), .A2(new_n835), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n847), .B1(new_n859), .B2(new_n576), .ZN(new_n860));
  OAI221_X1 g659(.A(new_n848), .B1(new_n849), .B2(new_n858), .C1(new_n860), .C2(KEYINPUT59), .ZN(G1345gat));
  NOR2_X1   g660(.A1(new_n840), .A2(new_n466), .ZN(new_n862));
  XNOR2_X1  g661(.A(new_n862), .B(KEYINPUT121), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n466), .A2(new_n269), .ZN(new_n864));
  AOI22_X1  g663(.A1(new_n863), .A2(new_n269), .B1(new_n859), .B2(new_n864), .ZN(G1346gat));
  AOI21_X1  g664(.A(G162gat), .B1(new_n846), .B2(new_n647), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n859), .A2(new_n647), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n866), .B1(new_n867), .B2(G162gat), .ZN(G1347gat));
  AND2_X1   g667(.A1(new_n702), .A2(new_n255), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n792), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(G169gat), .B1(new_n870), .B2(new_n616), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n792), .A2(new_n622), .A3(new_n255), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n872), .A2(G169gat), .ZN(new_n873));
  AND3_X1   g672(.A1(new_n873), .A2(KEYINPUT122), .A3(new_n617), .ZN(new_n874));
  AOI21_X1  g673(.A(KEYINPUT122), .B1(new_n873), .B2(new_n617), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n871), .B1(new_n874), .B2(new_n875), .ZN(G1348gat));
  NOR3_X1   g675(.A1(new_n870), .A2(new_n204), .A3(new_n649), .ZN(new_n877));
  INV_X1    g676(.A(new_n872), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(new_n576), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n877), .B1(new_n879), .B2(new_n204), .ZN(G1349gat));
  INV_X1    g679(.A(new_n870), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n213), .B1(new_n881), .B2(new_n467), .ZN(new_n882));
  INV_X1    g681(.A(new_n226), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n872), .A2(new_n466), .A3(new_n883), .ZN(new_n884));
  OR3_X1    g683(.A1(new_n882), .A2(new_n884), .A3(KEYINPUT60), .ZN(new_n885));
  OAI21_X1  g684(.A(KEYINPUT60), .B1(new_n882), .B2(new_n884), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(G1350gat));
  AOI21_X1  g686(.A(new_n214), .B1(new_n881), .B2(new_n647), .ZN(new_n888));
  XOR2_X1   g687(.A(KEYINPUT123), .B(KEYINPUT61), .Z(new_n889));
  OR2_X1    g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n878), .A2(new_n214), .A3(new_n647), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n888), .A2(new_n889), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(G1351gat));
  NOR3_X1   g692(.A1(new_n845), .A2(new_n623), .A3(new_n390), .ZN(new_n894));
  INV_X1    g693(.A(G197gat), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n894), .A2(new_n895), .A3(new_n617), .ZN(new_n896));
  XNOR2_X1  g695(.A(new_n896), .B(KEYINPUT124), .ZN(new_n897));
  AND3_X1   g696(.A1(new_n702), .A2(new_n255), .A3(new_n640), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n857), .A2(new_n617), .A3(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT125), .ZN(new_n900));
  OR2_X1    g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n899), .A2(new_n900), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n901), .A2(G197gat), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n897), .A2(new_n903), .ZN(G1352gat));
  INV_X1    g703(.A(G204gat), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n894), .A2(new_n905), .A3(new_n576), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT62), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n907), .A2(KEYINPUT126), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n907), .A2(KEYINPUT126), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n906), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  AND3_X1   g709(.A1(new_n857), .A2(new_n700), .A3(new_n898), .ZN(new_n911));
  OAI221_X1 g710(.A(new_n910), .B1(new_n905), .B2(new_n911), .C1(new_n908), .C2(new_n906), .ZN(G1353gat));
  NAND3_X1  g711(.A1(new_n857), .A2(new_n467), .A3(new_n898), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT127), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND4_X1  g714(.A1(new_n857), .A2(KEYINPUT127), .A3(new_n467), .A4(new_n898), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n915), .A2(G211gat), .A3(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT63), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND4_X1  g718(.A1(new_n915), .A2(KEYINPUT63), .A3(G211gat), .A4(new_n916), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n894), .A2(new_n241), .A3(new_n467), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(G1354gat));
  NAND3_X1  g722(.A1(new_n894), .A2(new_n242), .A3(new_n647), .ZN(new_n924));
  AND3_X1   g723(.A1(new_n857), .A2(new_n647), .A3(new_n898), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n924), .B1(new_n925), .B2(new_n242), .ZN(G1355gat));
endmodule


