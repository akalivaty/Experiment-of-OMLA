//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 1 1 0 0 1 1 0 1 0 0 1 0 0 0 1 0 0 1 1 0 1 0 0 0 1 1 0 0 0 0 1 1 1 0 1 0 1 0 1 0 1 1 1 0 1 0 0 0 0 0 1 1 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:56 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n203), .A2(G50), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  OR3_X1    g0014(.A1(new_n213), .A2(new_n207), .A3(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n216));
  INV_X1    g0016(.A(G238), .ZN(new_n217));
  INV_X1    g0017(.A(G87), .ZN(new_n218));
  INV_X1    g0018(.A(G250), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n216), .B1(new_n202), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n221));
  INV_X1    g0021(.A(G232), .ZN(new_n222));
  INV_X1    g0022(.A(G97), .ZN(new_n223));
  INV_X1    g0023(.A(G257), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n221), .B1(new_n201), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n209), .B1(new_n220), .B2(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n212), .B(new_n215), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(new_n222), .ZN(new_n230));
  XOR2_X1   g0030(.A(KEYINPUT2), .B(G226), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G264), .B(G270), .Z(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XOR2_X1   g0036(.A(G107), .B(G116), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT64), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G87), .B(G97), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G58), .B(G77), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  INV_X1    g0044(.A(G33), .ZN(new_n245));
  NOR2_X1   g0045(.A1(new_n245), .A2(KEYINPUT3), .ZN(new_n246));
  INV_X1    g0046(.A(KEYINPUT3), .ZN(new_n247));
  NOR2_X1   g0047(.A1(new_n247), .A2(G33), .ZN(new_n248));
  OAI21_X1  g0048(.A(KEYINPUT66), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n247), .A2(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n245), .A2(KEYINPUT3), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT66), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n250), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n249), .A2(new_n253), .ZN(new_n254));
  AND2_X1   g0054(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n255));
  NOR2_X1   g0055(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n254), .A2(G222), .A3(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n254), .A2(G223), .A3(G1698), .ZN(new_n259));
  INV_X1    g0059(.A(G77), .ZN(new_n260));
  OAI211_X1 g0060(.A(new_n258), .B(new_n259), .C1(new_n260), .C2(new_n254), .ZN(new_n261));
  INV_X1    g0061(.A(G41), .ZN(new_n262));
  OAI211_X1 g0062(.A(G1), .B(G13), .C1(new_n245), .C2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n261), .A2(new_n264), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n266));
  INV_X1    g0066(.A(G274), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT65), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  OAI211_X1 g0070(.A(new_n206), .B(KEYINPUT65), .C1(G41), .C2(G45), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n270), .A2(new_n271), .A3(new_n263), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n268), .B1(new_n273), .B2(G226), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n265), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G200), .ZN(new_n276));
  NAND3_X1  g0076(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(new_n214), .ZN(new_n278));
  OAI21_X1  g0078(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n279));
  INV_X1    g0079(.A(G150), .ZN(new_n280));
  NOR2_X1   g0080(.A1(G20), .A2(G33), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n279), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  AND2_X1   g0083(.A1(KEYINPUT8), .A2(G58), .ZN(new_n284));
  NOR2_X1   g0084(.A1(KEYINPUT8), .A2(G58), .ZN(new_n285));
  OR2_X1    g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n245), .A2(G20), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n278), .B1(new_n283), .B2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G13), .ZN(new_n291));
  NOR3_X1   g0091(.A1(new_n291), .A2(new_n207), .A3(G1), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n292), .A2(new_n278), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n206), .A2(G20), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n293), .A2(G50), .A3(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n292), .ZN(new_n296));
  OAI211_X1 g0096(.A(new_n290), .B(new_n295), .C1(G50), .C2(new_n296), .ZN(new_n297));
  XNOR2_X1  g0097(.A(new_n297), .B(KEYINPUT9), .ZN(new_n298));
  INV_X1    g0098(.A(G190), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n276), .B(new_n298), .C1(new_n299), .C2(new_n275), .ZN(new_n300));
  XNOR2_X1  g0100(.A(new_n300), .B(KEYINPUT10), .ZN(new_n301));
  INV_X1    g0101(.A(new_n275), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n297), .B1(new_n302), .B2(G169), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n275), .A2(G179), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n301), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  XNOR2_X1  g0108(.A(KEYINPUT67), .B(G1698), .ZN(new_n309));
  INV_X1    g0109(.A(G226), .ZN(new_n310));
  INV_X1    g0110(.A(G1698), .ZN(new_n311));
  OAI22_X1  g0111(.A1(new_n309), .A2(new_n310), .B1(new_n222), .B2(new_n311), .ZN(new_n312));
  AOI22_X1  g0112(.A1(new_n254), .A2(new_n312), .B1(G33), .B2(G97), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n313), .A2(new_n263), .ZN(new_n314));
  INV_X1    g0114(.A(new_n268), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n315), .B1(new_n272), .B2(new_n217), .ZN(new_n316));
  OR3_X1    g0116(.A1(new_n314), .A2(KEYINPUT13), .A3(new_n316), .ZN(new_n317));
  OAI21_X1  g0117(.A(KEYINPUT13), .B1(new_n314), .B2(new_n316), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n317), .A2(new_n318), .A3(G190), .ZN(new_n319));
  OR2_X1    g0119(.A1(new_n293), .A2(KEYINPUT68), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n293), .A2(KEYINPUT68), .ZN(new_n321));
  AND2_X1   g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n322), .A2(G68), .A3(new_n294), .ZN(new_n323));
  AOI22_X1  g0123(.A1(new_n281), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n324), .B1(new_n288), .B2(new_n260), .ZN(new_n325));
  AND2_X1   g0125(.A1(new_n325), .A2(new_n278), .ZN(new_n326));
  OR2_X1    g0126(.A1(new_n326), .A2(KEYINPUT11), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(KEYINPUT11), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n292), .A2(new_n202), .ZN(new_n329));
  XNOR2_X1  g0129(.A(new_n329), .B(KEYINPUT12), .ZN(new_n330));
  AND4_X1   g0130(.A1(new_n323), .A2(new_n327), .A3(new_n328), .A4(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n319), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(G200), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n333), .B1(new_n317), .B2(new_n318), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n317), .A2(new_n318), .A3(G179), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(KEYINPUT70), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT70), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n317), .A2(new_n318), .A3(new_n338), .A4(G179), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(G169), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n341), .B1(new_n317), .B2(new_n318), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT69), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n343), .A2(KEYINPUT14), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n343), .A2(KEYINPUT14), .ZN(new_n346));
  AND2_X1   g0146(.A1(new_n342), .A2(new_n346), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n340), .B(new_n345), .C1(new_n347), .C2(new_n344), .ZN(new_n348));
  INV_X1    g0148(.A(new_n331), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n335), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n322), .A2(G77), .A3(new_n294), .ZN(new_n351));
  XNOR2_X1  g0151(.A(KEYINPUT15), .B(G87), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n353), .A2(new_n287), .B1(G20), .B2(G77), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n354), .B1(new_n282), .B2(new_n286), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n355), .A2(new_n278), .B1(new_n260), .B2(new_n292), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n351), .A2(new_n356), .ZN(new_n357));
  AND3_X1   g0157(.A1(new_n250), .A2(new_n251), .A3(new_n252), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n252), .B1(new_n250), .B2(new_n251), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(G107), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n263), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  OAI22_X1  g0162(.A1(new_n309), .A2(new_n222), .B1(new_n217), .B2(new_n311), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n362), .B1(new_n360), .B2(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n268), .B1(new_n273), .B2(G244), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n357), .B1(G200), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n367), .B1(new_n299), .B2(new_n366), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n366), .A2(new_n341), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n369), .B(new_n357), .C1(G179), .C2(new_n366), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n308), .A2(new_n350), .A3(new_n368), .A4(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n286), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(new_n294), .ZN(new_n373));
  INV_X1    g0173(.A(new_n293), .ZN(new_n374));
  OAI22_X1  g0174(.A1(new_n373), .A2(new_n374), .B1(new_n296), .B2(new_n372), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT73), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n377), .B1(new_n245), .B2(KEYINPUT3), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n247), .A2(KEYINPUT73), .A3(G33), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n378), .A2(new_n251), .A3(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT74), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT7), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n382), .A2(G20), .ZN(new_n383));
  AND3_X1   g0183(.A1(new_n380), .A2(new_n381), .A3(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n381), .B1(new_n380), .B2(new_n383), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(KEYINPUT7), .B1(new_n360), .B2(new_n207), .ZN(new_n387));
  OAI21_X1  g0187(.A(G68), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(G159), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n282), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(G58), .A2(G68), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n207), .B1(new_n203), .B2(new_n391), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(KEYINPUT16), .B1(new_n388), .B2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT72), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(KEYINPUT72), .B1(new_n390), .B2(new_n392), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT71), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n399), .B1(new_n247), .B2(G33), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n245), .A2(KEYINPUT71), .A3(KEYINPUT3), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(new_n250), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n403), .A2(new_n382), .A3(new_n207), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n246), .B1(new_n400), .B2(new_n401), .ZN(new_n405));
  OAI21_X1  g0205(.A(KEYINPUT7), .B1(new_n405), .B2(G20), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n404), .A2(G68), .A3(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n398), .A2(new_n407), .A3(KEYINPUT16), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(new_n278), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n376), .B1(new_n394), .B2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(G223), .ZN(new_n411));
  OAI22_X1  g0211(.A1(new_n309), .A2(new_n411), .B1(new_n310), .B2(new_n311), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n405), .ZN(new_n413));
  NAND2_X1  g0213(.A1(G33), .A2(G87), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n264), .ZN(new_n416));
  INV_X1    g0216(.A(G179), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n270), .A2(G232), .A3(new_n263), .A4(new_n271), .ZN(new_n419));
  AOI21_X1  g0219(.A(KEYINPUT75), .B1(new_n419), .B2(new_n315), .ZN(new_n420));
  INV_X1    g0220(.A(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n419), .A2(KEYINPUT75), .A3(new_n315), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n419), .A2(new_n315), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n424), .B1(new_n415), .B2(new_n264), .ZN(new_n425));
  OAI22_X1  g0225(.A1(new_n418), .A2(new_n423), .B1(new_n425), .B2(G169), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n410), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT18), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n393), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n249), .A2(new_n207), .A3(new_n253), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(new_n382), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n433), .B1(new_n384), .B2(new_n385), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n431), .B1(new_n434), .B2(G68), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n278), .B(new_n408), .C1(new_n435), .C2(KEYINPUT16), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n426), .B1(new_n436), .B2(new_n376), .ZN(new_n437));
  OAI21_X1  g0237(.A(KEYINPUT76), .B1(new_n437), .B2(KEYINPUT18), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT76), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n428), .A2(new_n439), .A3(new_n429), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n430), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  AND2_X1   g0241(.A1(new_n299), .A2(KEYINPUT77), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n299), .A2(KEYINPUT77), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  AOI22_X1  g0244(.A1(new_n412), .A2(new_n405), .B1(G33), .B2(G87), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n444), .B1(new_n445), .B2(new_n263), .ZN(new_n446));
  OAI21_X1  g0246(.A(KEYINPUT78), .B1(new_n423), .B2(new_n446), .ZN(new_n447));
  AND3_X1   g0247(.A1(new_n419), .A2(KEYINPUT75), .A3(new_n315), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n448), .A2(new_n420), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT78), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n449), .A2(new_n416), .A3(new_n450), .A4(new_n444), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n445), .A2(new_n263), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n333), .B1(new_n452), .B2(new_n424), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n447), .A2(new_n451), .A3(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n454), .A2(new_n436), .A3(new_n376), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT17), .ZN(new_n456));
  XNOR2_X1  g0256(.A(new_n455), .B(new_n456), .ZN(new_n457));
  OR2_X1    g0257(.A1(new_n441), .A2(new_n457), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n371), .A2(new_n458), .ZN(new_n459));
  OR3_X1    g0259(.A1(new_n296), .A2(KEYINPUT79), .A3(G97), .ZN(new_n460));
  OAI21_X1  g0260(.A(KEYINPUT79), .B1(new_n296), .B2(G97), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n206), .A2(G33), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n293), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n462), .B1(new_n223), .B2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT6), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n223), .A2(new_n361), .ZN(new_n468));
  NOR2_X1   g0268(.A1(G97), .A2(G107), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n361), .A2(KEYINPUT6), .A3(G97), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n472), .A2(G20), .B1(G77), .B2(new_n281), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n474), .B1(new_n434), .B2(G107), .ZN(new_n475));
  INV_X1    g0275(.A(new_n278), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n466), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n402), .A2(G244), .A3(new_n250), .A4(new_n257), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT4), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  OAI211_X1 g0280(.A(G250), .B(G1698), .C1(new_n358), .C2(new_n359), .ZN(new_n481));
  AND2_X1   g0281(.A1(KEYINPUT4), .A2(G244), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n257), .B(new_n482), .C1(new_n358), .C2(new_n359), .ZN(new_n483));
  NAND2_X1  g0283(.A1(G33), .A2(G283), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n480), .A2(new_n481), .A3(new_n483), .A4(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(new_n264), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n206), .B(G45), .C1(new_n262), .C2(KEYINPUT5), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT80), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(G45), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n490), .A2(G1), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT5), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(G41), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n491), .A2(KEYINPUT80), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n262), .A2(KEYINPUT5), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n489), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n496), .A2(G257), .A3(new_n263), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n487), .A2(new_n488), .B1(KEYINPUT5), .B2(new_n262), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n498), .A2(G274), .A3(new_n263), .A4(new_n494), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n486), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n341), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n500), .B1(new_n485), .B2(new_n264), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n417), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n477), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n380), .A2(new_n383), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(KEYINPUT74), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n380), .A2(new_n381), .A3(new_n383), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n508), .A2(new_n509), .B1(new_n432), .B2(new_n382), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n473), .B1(new_n510), .B2(new_n361), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n465), .B1(new_n511), .B2(new_n278), .ZN(new_n512));
  AOI211_X1 g0312(.A(G190), .B(new_n500), .C1(new_n264), .C2(new_n485), .ZN(new_n513));
  AOI21_X1  g0313(.A(G200), .B1(new_n486), .B2(new_n501), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n506), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(KEYINPUT81), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT81), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n506), .A2(new_n515), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT24), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n402), .A2(new_n207), .A3(G87), .A4(new_n250), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(KEYINPUT22), .ZN(new_n523));
  NOR3_X1   g0323(.A1(new_n218), .A2(KEYINPUT22), .A3(G20), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n524), .B1(new_n358), .B2(new_n359), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT23), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n527), .B1(new_n207), .B2(G107), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n361), .A2(KEYINPUT23), .A3(G20), .ZN(new_n529));
  NAND2_X1  g0329(.A1(G33), .A2(G116), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n528), .A2(new_n529), .B1(new_n531), .B2(new_n207), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n521), .B1(new_n526), .B2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(new_n532), .ZN(new_n534));
  AOI211_X1 g0334(.A(KEYINPUT24), .B(new_n534), .C1(new_n523), .C2(new_n525), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n278), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(new_n464), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT25), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n538), .B1(new_n296), .B2(G107), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n292), .A2(KEYINPUT25), .A3(new_n361), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n537), .A2(G107), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n536), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(KEYINPUT84), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT84), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n536), .A2(new_n544), .A3(new_n541), .ZN(new_n545));
  NOR3_X1   g0345(.A1(new_n255), .A2(new_n256), .A3(new_n219), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n224), .A2(new_n311), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n405), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(G33), .A2(G294), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n264), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n264), .B1(new_n498), .B2(new_n494), .ZN(new_n552));
  AOI21_X1  g0352(.A(KEYINPUT85), .B1(new_n552), .B2(G264), .ZN(new_n553));
  AND4_X1   g0353(.A1(KEYINPUT85), .A2(new_n496), .A3(G264), .A4(new_n263), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n499), .B(new_n551), .C1(new_n553), .C2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(G169), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT86), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n263), .B1(new_n548), .B2(new_n549), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n496), .A2(G264), .A3(new_n263), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT85), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n552), .A2(KEYINPUT85), .A3(G264), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n558), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n563), .A2(G179), .A3(new_n499), .ZN(new_n564));
  AND3_X1   g0364(.A1(new_n556), .A2(new_n557), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n557), .B1(new_n556), .B2(new_n564), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n543), .B(new_n545), .C1(new_n565), .C2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n555), .A2(G200), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n563), .A2(G190), .A3(new_n499), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n568), .A2(new_n536), .A3(new_n569), .A4(new_n541), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(G116), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n572), .B1(new_n206), .B2(G33), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n320), .A2(new_n321), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n572), .A2(G20), .ZN(new_n575));
  NOR3_X1   g0375(.A1(new_n575), .A2(G1), .A3(new_n291), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n484), .B(new_n207), .C1(G33), .C2(new_n223), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n577), .A2(KEYINPUT20), .A3(new_n278), .A4(new_n575), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n577), .A2(new_n278), .A3(new_n575), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT20), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n576), .B1(new_n578), .B2(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n341), .B1(new_n574), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n496), .A2(G270), .A3(new_n263), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT83), .ZN(new_n585));
  XNOR2_X1  g0385(.A(new_n584), .B(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(G303), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n257), .A2(G257), .B1(G264), .B2(G1698), .ZN(new_n588));
  OAI22_X1  g0388(.A1(new_n254), .A2(new_n587), .B1(new_n588), .B2(new_n403), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n264), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n499), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n583), .B(KEYINPUT21), .C1(new_n586), .C2(new_n591), .ZN(new_n592));
  XNOR2_X1  g0392(.A(new_n584), .B(KEYINPUT83), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n574), .A2(new_n582), .ZN(new_n594));
  INV_X1    g0394(.A(new_n499), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n595), .B1(new_n589), .B2(new_n264), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n593), .A2(G179), .A3(new_n594), .A4(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n592), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n593), .A2(new_n596), .ZN(new_n599));
  AOI21_X1  g0399(.A(KEYINPUT21), .B1(new_n599), .B2(new_n583), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n309), .A2(new_n217), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n531), .B1(new_n602), .B2(new_n405), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n405), .A2(G244), .A3(G1698), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n603), .A2(KEYINPUT82), .A3(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(KEYINPUT82), .B1(new_n603), .B2(new_n604), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n264), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n491), .A2(new_n219), .ZN(new_n609));
  AOI22_X1  g0409(.A1(new_n609), .A2(new_n263), .B1(G274), .B2(new_n491), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n608), .A2(new_n417), .A3(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n405), .A2(new_n207), .A3(G68), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n287), .A2(G97), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT19), .ZN(new_n614));
  NAND3_X1  g0414(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n207), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n469), .A2(new_n218), .ZN(new_n617));
  AOI22_X1  g0417(.A1(new_n613), .A2(new_n614), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n612), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n278), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n352), .A2(new_n292), .ZN(new_n621));
  AND2_X1   g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n622), .B1(new_n352), .B2(new_n464), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n602), .A2(new_n405), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n624), .A2(new_n604), .A3(new_n530), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT82), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n263), .B1(new_n627), .B2(new_n605), .ZN(new_n628));
  INV_X1    g0428(.A(new_n610), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n611), .B(new_n623), .C1(new_n630), .C2(G169), .ZN(new_n631));
  OAI21_X1  g0431(.A(G200), .B1(new_n628), .B2(new_n629), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n608), .A2(G190), .A3(new_n610), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n537), .A2(G87), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n632), .A2(new_n633), .A3(new_n622), .A4(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(G200), .B1(new_n586), .B2(new_n591), .ZN(new_n636));
  INV_X1    g0436(.A(new_n594), .ZN(new_n637));
  INV_X1    g0437(.A(new_n444), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n593), .A2(new_n638), .A3(new_n596), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n636), .A2(new_n637), .A3(new_n639), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n601), .A2(new_n631), .A3(new_n635), .A4(new_n640), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n571), .A2(new_n641), .ZN(new_n642));
  AND3_X1   g0442(.A1(new_n459), .A2(new_n520), .A3(new_n642), .ZN(G372));
  NAND3_X1  g0443(.A1(new_n620), .A2(new_n634), .A3(new_n621), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(KEYINPUT88), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT88), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n620), .A2(new_n634), .A3(new_n646), .A4(new_n621), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  AND3_X1   g0448(.A1(new_n632), .A2(new_n633), .A3(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(KEYINPUT87), .B1(new_n630), .B2(G169), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n608), .A2(new_n610), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT87), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n651), .A2(new_n652), .A3(new_n341), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n611), .A2(new_n623), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n649), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT26), .ZN(new_n658));
  INV_X1    g0458(.A(new_n506), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n657), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n655), .B1(new_n650), .B2(new_n653), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n659), .A2(new_n631), .A3(new_n635), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n661), .B1(new_n662), .B2(KEYINPUT26), .ZN(new_n663));
  INV_X1    g0463(.A(new_n570), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n516), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n657), .A2(new_n665), .ZN(new_n666));
  AOI22_X1  g0466(.A1(new_n556), .A2(new_n564), .B1(new_n536), .B2(new_n541), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n601), .A2(new_n668), .A3(KEYINPUT89), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT89), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n583), .B1(new_n586), .B2(new_n591), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT21), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n673), .A2(new_n592), .A3(new_n597), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n670), .B1(new_n674), .B2(new_n667), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n669), .A2(new_n675), .ZN(new_n676));
  OAI211_X1 g0476(.A(new_n660), .B(new_n663), .C1(new_n666), .C2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n459), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n428), .A2(new_n429), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n437), .A2(KEYINPUT18), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n335), .A2(new_n370), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n682), .B1(new_n348), .B2(new_n349), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n681), .B1(new_n683), .B2(new_n457), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n305), .B1(new_n684), .B2(new_n301), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n678), .A2(new_n685), .ZN(G369));
  INV_X1    g0486(.A(KEYINPUT94), .ZN(new_n687));
  AND3_X1   g0487(.A1(new_n536), .A2(new_n544), .A3(new_n541), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n544), .B1(new_n536), .B2(new_n541), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n555), .A2(new_n417), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n341), .B1(new_n563), .B2(new_n499), .ZN(new_n692));
  OAI21_X1  g0492(.A(KEYINPUT86), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n556), .A2(new_n564), .A3(new_n557), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n664), .B1(new_n690), .B2(new_n695), .ZN(new_n696));
  NOR3_X1   g0496(.A1(new_n291), .A2(G1), .A3(G20), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT27), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g0499(.A(new_n699), .B(KEYINPUT90), .ZN(new_n700));
  INV_X1    g0500(.A(G213), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n701), .B1(new_n697), .B2(new_n698), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT91), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n700), .A2(KEYINPUT91), .A3(new_n702), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n708), .A2(G343), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n690), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n696), .A2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n567), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(new_n709), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g0514(.A(new_n714), .B(KEYINPUT93), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n674), .A2(new_n594), .A3(new_n709), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT92), .ZN(new_n717));
  INV_X1    g0517(.A(new_n709), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n718), .A2(new_n637), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n640), .A2(new_n673), .A3(new_n592), .A4(new_n597), .ZN(new_n720));
  OAI211_X1 g0520(.A(new_n716), .B(new_n717), .C1(new_n719), .C2(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n719), .A2(KEYINPUT92), .A3(new_n674), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(G330), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n687), .B1(new_n715), .B2(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n714), .A2(KEYINPUT93), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT93), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n728), .B1(new_n711), .B2(new_n713), .ZN(new_n729));
  OAI211_X1 g0529(.A(new_n725), .B(new_n687), .C1(new_n727), .C2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n726), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  XNOR2_X1  g0533(.A(new_n709), .B(KEYINPUT95), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(new_n668), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n601), .A2(new_n709), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n736), .B1(new_n715), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n733), .A2(new_n738), .ZN(G399));
  INV_X1    g0539(.A(new_n210), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(G41), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n617), .A2(G116), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n742), .A2(G1), .A3(new_n743), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n744), .B1(new_n213), .B2(new_n742), .ZN(new_n745));
  XOR2_X1   g0545(.A(KEYINPUT96), .B(KEYINPUT28), .Z(new_n746));
  XNOR2_X1  g0546(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n593), .A2(G179), .A3(new_n596), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n651), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT30), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(KEYINPUT97), .ZN(new_n751));
  AND3_X1   g0551(.A1(new_n504), .A2(new_n563), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n749), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n750), .A2(KEYINPUT97), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  OAI211_X1 g0555(.A(new_n749), .B(new_n752), .C1(KEYINPUT97), .C2(new_n750), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  AOI21_X1  g0557(.A(G179), .B1(new_n593), .B2(new_n596), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n758), .A2(new_n502), .A3(new_n555), .A4(new_n651), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n760), .A2(KEYINPUT31), .A3(new_n735), .ZN(new_n761));
  AOI21_X1  g0561(.A(KEYINPUT31), .B1(new_n760), .B2(new_n709), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n635), .A2(new_n631), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n720), .ZN(new_n765));
  NAND4_X1  g0565(.A1(new_n520), .A2(new_n696), .A3(new_n765), .A4(new_n734), .ZN(new_n766));
  INV_X1    g0566(.A(KEYINPUT98), .ZN(new_n767));
  AND2_X1   g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n766), .A2(new_n767), .ZN(new_n769));
  OAI211_X1 g0569(.A(new_n761), .B(new_n763), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G330), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n658), .B1(new_n657), .B2(new_n659), .ZN(new_n772));
  INV_X1    g0572(.A(new_n661), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n773), .B1(new_n662), .B2(KEYINPUT26), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  OAI211_X1 g0575(.A(new_n657), .B(new_n665), .C1(new_n712), .C2(new_n674), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n709), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(KEYINPUT29), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n677), .A2(new_n734), .ZN(new_n779));
  XOR2_X1   g0579(.A(KEYINPUT99), .B(KEYINPUT29), .Z(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n778), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n771), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n747), .B1(new_n784), .B2(G1), .ZN(G364));
  NOR2_X1   g0585(.A1(new_n291), .A2(G20), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n206), .B1(new_n786), .B2(G45), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n741), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n725), .A2(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(G330), .B1(new_n721), .B2(new_n722), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(G13), .A2(G33), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(G20), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n723), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n789), .ZN(new_n797));
  OAI21_X1  g0597(.A(G20), .B1(KEYINPUT100), .B2(G169), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(KEYINPUT100), .A2(G169), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n214), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NOR3_X1   g0602(.A1(new_n207), .A2(new_n417), .A3(new_n333), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(G190), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  XOR2_X1   g0606(.A(KEYINPUT33), .B(G317), .Z(new_n807));
  INV_X1    g0607(.A(G283), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n207), .A2(G179), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n809), .A2(new_n299), .A3(G200), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n806), .A2(new_n807), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n809), .A2(G190), .A3(G200), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  AOI211_X1 g0613(.A(new_n254), .B(new_n811), .C1(G303), .C2(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(G179), .A2(G200), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(G190), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(G20), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(G294), .ZN(new_n819));
  NOR3_X1   g0619(.A1(new_n207), .A2(new_n417), .A3(G200), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(new_n299), .ZN(new_n821));
  INV_X1    g0621(.A(G311), .ZN(new_n822));
  OAI22_X1  g0622(.A1(new_n818), .A2(new_n819), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n804), .A2(new_n444), .ZN(new_n824));
  AND2_X1   g0624(.A1(new_n824), .A2(G326), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n638), .A2(new_n820), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n823), .B(new_n825), .C1(G322), .C2(new_n827), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n815), .A2(G20), .A3(new_n299), .ZN(new_n829));
  OR2_X1    g0629(.A1(new_n829), .A2(KEYINPUT101), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(KEYINPUT101), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(G329), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n814), .A2(new_n828), .A3(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n832), .A2(new_n389), .ZN(new_n836));
  XNOR2_X1  g0636(.A(new_n836), .B(KEYINPUT32), .ZN(new_n837));
  INV_X1    g0637(.A(new_n824), .ZN(new_n838));
  INV_X1    g0638(.A(G50), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n838), .A2(new_n839), .B1(new_n260), .B2(new_n821), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n813), .A2(G87), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n841), .B1(new_n361), .B2(new_n810), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n360), .B1(new_n827), .B2(G58), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n805), .A2(G68), .B1(G97), .B2(new_n817), .ZN(new_n845));
  NAND4_X1  g0645(.A1(new_n837), .A2(new_n843), .A3(new_n844), .A4(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n802), .B1(new_n835), .B2(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n801), .A2(new_n795), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n254), .A2(G355), .A3(new_n210), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n740), .A2(new_n405), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n850), .B1(G45), .B2(new_n213), .ZN(new_n851));
  AND2_X1   g0651(.A1(new_n243), .A2(G45), .ZN(new_n852));
  OAI221_X1 g0652(.A(new_n849), .B1(G116), .B2(new_n210), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  AOI211_X1 g0653(.A(new_n797), .B(new_n847), .C1(new_n848), .C2(new_n853), .ZN(new_n854));
  AOI22_X1  g0654(.A1(new_n790), .A2(new_n792), .B1(new_n796), .B2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(G396));
  INV_X1    g0656(.A(new_n771), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n709), .A2(new_n357), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n368), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(new_n370), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n709), .A2(new_n370), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  XNOR2_X1  g0664(.A(new_n779), .B(new_n864), .ZN(new_n865));
  OR3_X1    g0665(.A1(new_n857), .A2(KEYINPUT104), .A3(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(KEYINPUT104), .B1(new_n857), .B2(new_n865), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n789), .B1(new_n857), .B2(new_n865), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n802), .A2(new_n794), .ZN(new_n870));
  XOR2_X1   g0670(.A(new_n870), .B(KEYINPUT102), .Z(new_n871));
  OAI21_X1  g0671(.A(new_n789), .B1(new_n871), .B2(G77), .ZN(new_n872));
  XOR2_X1   g0672(.A(new_n872), .B(KEYINPUT103), .Z(new_n873));
  AOI22_X1  g0673(.A1(new_n827), .A2(G143), .B1(G150), .B2(new_n805), .ZN(new_n874));
  INV_X1    g0674(.A(new_n821), .ZN(new_n875));
  AOI22_X1  g0675(.A1(new_n824), .A2(G137), .B1(new_n875), .B2(G159), .ZN(new_n876));
  AND2_X1   g0676(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  OR2_X1    g0677(.A1(new_n877), .A2(KEYINPUT34), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n874), .A2(KEYINPUT34), .A3(new_n876), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n405), .B1(new_n202), .B2(new_n810), .ZN(new_n880));
  OAI22_X1  g0680(.A1(new_n818), .A2(new_n201), .B1(new_n839), .B2(new_n812), .ZN(new_n881));
  AOI211_X1 g0681(.A(new_n880), .B(new_n881), .C1(new_n833), .C2(G132), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n878), .A2(new_n879), .A3(new_n882), .ZN(new_n883));
  OAI22_X1  g0683(.A1(new_n810), .A2(new_n218), .B1(new_n812), .B2(new_n361), .ZN(new_n884));
  AOI211_X1 g0684(.A(new_n254), .B(new_n884), .C1(G97), .C2(new_n817), .ZN(new_n885));
  AOI22_X1  g0685(.A1(new_n805), .A2(G283), .B1(new_n875), .B2(G116), .ZN(new_n886));
  AOI22_X1  g0686(.A1(new_n827), .A2(G294), .B1(G303), .B2(new_n824), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n833), .A2(G311), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n885), .A2(new_n886), .A3(new_n887), .A4(new_n888), .ZN(new_n889));
  AND2_X1   g0689(.A1(new_n883), .A2(new_n889), .ZN(new_n890));
  OAI221_X1 g0690(.A(new_n873), .B1(new_n802), .B2(new_n890), .C1(new_n864), .C2(new_n794), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n869), .A2(new_n891), .ZN(G384));
  NAND3_X1  g0692(.A1(new_n459), .A2(new_n778), .A3(new_n781), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(new_n685), .ZN(new_n894));
  XOR2_X1   g0694(.A(new_n894), .B(KEYINPUT107), .Z(new_n895));
  AOI21_X1  g0695(.A(KEYINPUT16), .B1(new_n398), .B2(new_n407), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n376), .B1(new_n409), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n708), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n899), .B1(new_n441), .B2(new_n457), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT16), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n510), .A2(new_n202), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n901), .B1(new_n902), .B2(new_n431), .ZN(new_n903));
  AND2_X1   g0703(.A1(new_n408), .A2(new_n278), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n375), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n426), .A2(new_n707), .ZN(new_n906));
  AOI22_X1  g0706(.A1(new_n905), .A2(new_n454), .B1(new_n906), .B2(new_n897), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT37), .ZN(new_n908));
  OAI21_X1  g0708(.A(KEYINPUT106), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n906), .A2(new_n897), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n455), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT106), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n911), .A2(new_n912), .A3(KEYINPUT37), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n410), .A2(new_n708), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n428), .A2(new_n914), .A3(new_n455), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n909), .B(new_n913), .C1(KEYINPUT37), .C2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n900), .A2(KEYINPUT38), .A3(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT38), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n915), .B(new_n908), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n455), .A2(new_n456), .ZN(new_n920));
  AOI21_X1  g0720(.A(KEYINPUT17), .B1(new_n905), .B2(new_n454), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n914), .B1(new_n922), .B2(new_n681), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n918), .B1(new_n919), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n917), .A2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT39), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n348), .A2(new_n349), .A3(new_n718), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n900), .A2(new_n916), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n918), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n917), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n927), .B(new_n929), .C1(new_n932), .C2(new_n926), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n681), .A2(new_n708), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n718), .A2(new_n331), .ZN(new_n935));
  AND2_X1   g0735(.A1(new_n348), .A2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n935), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n936), .B1(new_n350), .B2(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n677), .A2(new_n734), .A3(new_n864), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n938), .B1(new_n939), .B2(new_n862), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n934), .B1(new_n940), .B2(new_n932), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n933), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n895), .B(new_n942), .ZN(new_n943));
  AOI211_X1 g0743(.A(new_n335), .B(new_n935), .C1(new_n348), .C2(new_n349), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n864), .B1(new_n944), .B2(new_n936), .ZN(new_n945));
  NAND4_X1  g0745(.A1(new_n642), .A2(KEYINPUT98), .A3(new_n520), .A4(new_n734), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n766), .A2(new_n767), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n762), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n760), .A2(KEYINPUT31), .A3(new_n709), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n945), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT40), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n951), .B1(new_n917), .B2(new_n924), .ZN(new_n952));
  AOI21_X1  g0752(.A(KEYINPUT109), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  OAI211_X1 g0753(.A(new_n763), .B(new_n949), .C1(new_n768), .C2(new_n769), .ZN(new_n954));
  INV_X1    g0754(.A(new_n945), .ZN(new_n955));
  AND4_X1   g0755(.A1(KEYINPUT109), .A2(new_n954), .A3(new_n952), .A4(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n953), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n932), .A2(new_n954), .A3(new_n955), .ZN(new_n958));
  XNOR2_X1  g0758(.A(KEYINPUT108), .B(KEYINPUT40), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n957), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n954), .A2(new_n459), .ZN(new_n962));
  AND2_X1   g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n961), .A2(new_n962), .ZN(new_n964));
  NOR3_X1   g0764(.A1(new_n963), .A2(new_n964), .A3(new_n724), .ZN(new_n965));
  OAI22_X1  g0765(.A1(new_n943), .A2(new_n965), .B1(new_n206), .B2(new_n786), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n966), .B1(new_n943), .B2(new_n965), .ZN(new_n967));
  NOR3_X1   g0767(.A1(new_n214), .A2(new_n207), .A3(new_n572), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n472), .B(KEYINPUT105), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT35), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n968), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n972), .B1(new_n971), .B2(new_n970), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT36), .ZN(new_n974));
  NAND4_X1  g0774(.A1(new_n203), .A2(G50), .A3(G77), .A4(new_n391), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n839), .A2(G68), .ZN(new_n976));
  AOI211_X1 g0776(.A(new_n206), .B(G13), .C1(new_n975), .C2(new_n976), .ZN(new_n977));
  OR3_X1    g0777(.A1(new_n967), .A2(new_n974), .A3(new_n977), .ZN(G367));
  OAI211_X1 g0778(.A(new_n506), .B(new_n515), .C1(new_n734), .C2(new_n512), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n506), .B1(new_n979), .B2(new_n567), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(new_n734), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n735), .A2(new_n659), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(new_n979), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n715), .A2(new_n737), .A3(new_n983), .ZN(new_n984));
  XOR2_X1   g0784(.A(KEYINPUT110), .B(KEYINPUT42), .Z(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n981), .B1(new_n984), .B2(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n987), .B1(new_n984), .B2(new_n986), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT43), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n718), .A2(new_n648), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(new_n661), .ZN(new_n991));
  INV_X1    g0791(.A(new_n657), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n991), .B1(new_n992), .B2(new_n990), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n988), .A2(new_n989), .A3(new_n994), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n993), .A2(KEYINPUT43), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n993), .A2(KEYINPUT43), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n984), .A2(new_n986), .ZN(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  OAI211_X1 g0800(.A(new_n997), .B(new_n998), .C1(new_n1000), .C2(new_n987), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n995), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n983), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n733), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1002), .A2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(KEYINPUT111), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT111), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n995), .A2(new_n1001), .A3(new_n1008), .A4(new_n1004), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  XOR2_X1   g0810(.A(new_n741), .B(KEYINPUT41), .Z(new_n1011));
  INV_X1    g0811(.A(KEYINPUT114), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT113), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1012), .B1(new_n725), .B2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n1012), .B2(new_n725), .ZN(new_n1015));
  OR3_X1    g0815(.A1(new_n727), .A2(new_n729), .A3(new_n737), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n737), .B1(new_n727), .B2(new_n729), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1015), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  AND2_X1   g0818(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1014), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1018), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1021), .A2(new_n783), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT115), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n733), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT112), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n738), .A2(new_n1025), .A3(new_n983), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n736), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1017), .A2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(KEYINPUT112), .B1(new_n1028), .B2(new_n1003), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1026), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(KEYINPUT45), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT45), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1026), .A2(new_n1029), .A3(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT44), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n738), .B2(new_n983), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1028), .A2(KEYINPUT44), .A3(new_n1003), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n1036), .A2(new_n1037), .B1(new_n732), .B2(KEYINPUT115), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1024), .B1(new_n1034), .B2(new_n1038), .ZN(new_n1039));
  AND3_X1   g0839(.A1(new_n1026), .A2(new_n1029), .A3(new_n1032), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1032), .B1(new_n1026), .B2(new_n1029), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n1038), .B(new_n1024), .C1(new_n1040), .C2(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n1042), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1022), .B1(new_n1039), .B2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1011), .B1(new_n1044), .B2(new_n784), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n787), .B(KEYINPUT116), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n1006), .B(new_n1010), .C1(new_n1045), .C2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n994), .A2(new_n795), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n850), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n848), .B1(new_n210), .B2(new_n352), .C1(new_n1049), .C2(new_n235), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n797), .B1(new_n1050), .B2(KEYINPUT117), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(KEYINPUT117), .B2(new_n1050), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n806), .A2(new_n819), .B1(new_n821), .B2(new_n808), .ZN(new_n1053));
  AOI211_X1 g0853(.A(new_n405), .B(new_n1053), .C1(G107), .C2(new_n817), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n833), .A2(G317), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n813), .A2(G116), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT46), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n810), .A2(new_n223), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n826), .A2(new_n587), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n1058), .B(new_n1059), .C1(G311), .C2(new_n824), .ZN(new_n1060));
  NAND4_X1  g0860(.A1(new_n1054), .A2(new_n1055), .A3(new_n1057), .A4(new_n1060), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n833), .A2(G137), .B1(G58), .B2(new_n813), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n1062), .A2(KEYINPUT118), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1062), .A2(KEYINPUT118), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n810), .A2(new_n260), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n821), .A2(new_n839), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n1065), .B(new_n1066), .C1(G143), .C2(new_n824), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n360), .B1(new_n827), .B2(G150), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n805), .A2(G159), .B1(G68), .B2(new_n817), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n1064), .A2(new_n1067), .A3(new_n1068), .A4(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1061), .B1(new_n1063), .B2(new_n1070), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT47), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1052), .B1(new_n1072), .B2(new_n801), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1048), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1047), .A2(new_n1074), .ZN(G387));
  OAI211_X1 g0875(.A(new_n1018), .B(new_n1046), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n254), .A2(new_n210), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n1077), .A2(new_n743), .B1(G107), .B2(new_n210), .ZN(new_n1078));
  OR2_X1    g0878(.A1(new_n232), .A2(new_n490), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n743), .B(new_n490), .C1(new_n202), .C2(new_n260), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(KEYINPUT119), .B(KEYINPUT50), .ZN(new_n1081));
  NOR3_X1   g0881(.A1(new_n286), .A2(new_n1081), .A3(G50), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1081), .B1(new_n286), .B2(G50), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1049), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1078), .B1(new_n1079), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n848), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n789), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n805), .A2(new_n372), .B1(new_n875), .B2(G68), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT120), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n824), .A2(G159), .B1(G77), .B2(new_n813), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n827), .A2(G50), .B1(new_n353), .B2(new_n817), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n403), .B(new_n1058), .C1(new_n833), .C2(G150), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n1090), .A2(new_n1091), .A3(new_n1092), .A4(new_n1093), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n827), .A2(G317), .B1(G303), .B2(new_n875), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(G322), .A2(new_n824), .B1(new_n805), .B2(G311), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1095), .A2(KEYINPUT48), .A3(new_n1096), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n813), .A2(G294), .B1(new_n817), .B2(G283), .ZN(new_n1098));
  AND2_X1   g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  AND2_X1   g0899(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1099), .B1(KEYINPUT48), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT49), .ZN(new_n1102));
  AND2_X1   g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n403), .B1(new_n572), .B2(new_n810), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(new_n833), .B2(G326), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1105), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1094), .B1(new_n1103), .B2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1088), .B1(new_n1107), .B2(new_n801), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n795), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1108), .B1(new_n715), .B2(new_n1109), .ZN(new_n1110));
  AND2_X1   g0910(.A1(new_n1021), .A2(new_n783), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n741), .B1(new_n1021), .B2(new_n783), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n1076), .B(new_n1110), .C1(new_n1111), .C2(new_n1112), .ZN(G393));
  NOR2_X1   g0913(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1038), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n1023), .B(new_n733), .C1(new_n1114), .C2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1022), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1116), .A2(new_n1117), .A3(new_n1042), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1044), .A2(new_n1118), .A3(new_n741), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1116), .A2(new_n1042), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1003), .A2(new_n795), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n848), .B1(new_n223), .B2(new_n210), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1122), .B1(new_n240), .B2(new_n850), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n827), .A2(G311), .B1(G317), .B2(new_n824), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1124), .B(KEYINPUT52), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n833), .A2(G322), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n875), .A2(G294), .B1(new_n813), .B2(G283), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n805), .A2(G303), .B1(G116), .B2(new_n817), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n810), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n254), .B1(G107), .B2(new_n1129), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1126), .A2(new_n1127), .A3(new_n1128), .A4(new_n1130), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n827), .A2(G159), .B1(G150), .B2(new_n824), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n1132), .B(KEYINPUT51), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n833), .A2(G143), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n813), .A2(G68), .B1(new_n817), .B2(G77), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n805), .A2(G50), .B1(new_n875), .B2(new_n372), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n403), .B1(G87), .B2(new_n1129), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n1134), .A2(new_n1135), .A3(new_n1136), .A4(new_n1137), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n1125), .A2(new_n1131), .B1(new_n1133), .B2(new_n1138), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n797), .B(new_n1123), .C1(new_n1139), .C2(new_n801), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n1120), .A2(new_n1046), .B1(new_n1121), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1119), .A2(new_n1141), .ZN(G390));
  INV_X1    g0942(.A(new_n917), .ZN(new_n1143));
  AOI21_X1  g0943(.A(KEYINPUT38), .B1(new_n900), .B2(new_n916), .ZN(new_n1144));
  NOR3_X1   g0944(.A1(new_n1143), .A2(new_n1144), .A3(new_n926), .ZN(new_n1145));
  AOI21_X1  g0945(.A(KEYINPUT39), .B1(new_n917), .B2(new_n924), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n1145), .A2(new_n1146), .B1(new_n940), .B2(new_n929), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n861), .B1(new_n777), .B2(new_n860), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n928), .B(new_n925), .C1(new_n1148), .C2(new_n938), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n938), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n770), .A2(G330), .A3(new_n864), .A4(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1147), .A2(new_n1149), .A3(new_n1151), .ZN(new_n1152));
  AND2_X1   g0952(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n950), .A2(G330), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1152), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1151), .A2(new_n1148), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n724), .B1(new_n948), .B2(new_n949), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1150), .B1(new_n1157), .B2(new_n864), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT121), .ZN(new_n1160));
  AOI211_X1 g0960(.A(new_n724), .B(new_n863), .C1(new_n948), .C2(new_n761), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1160), .B1(new_n1161), .B2(new_n1150), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n770), .A2(G330), .A3(new_n864), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1163), .A2(KEYINPUT121), .A3(new_n938), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1162), .A2(new_n1154), .A3(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n939), .A2(new_n862), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1159), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  AND3_X1   g0967(.A1(new_n954), .A2(new_n459), .A3(G330), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n894), .A2(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1155), .B1(new_n1167), .B2(new_n1170), .ZN(new_n1171));
  AND3_X1   g0971(.A1(new_n1147), .A2(new_n1149), .A3(new_n1151), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1154), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1166), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1163), .A2(new_n938), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n1176), .A2(new_n1160), .B1(G330), .B2(new_n950), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1175), .B1(new_n1177), .B2(new_n1164), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1174), .B(new_n1169), .C1(new_n1178), .C2(new_n1159), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1171), .A2(new_n741), .A3(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n793), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n789), .B1(new_n871), .B2(new_n372), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n360), .B1(G137), .B2(new_n805), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(KEYINPUT54), .B(G143), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(new_n1184), .B(KEYINPUT122), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(new_n875), .ZN(new_n1186));
  INV_X1    g0986(.A(G125), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1183), .B(new_n1186), .C1(new_n1187), .C2(new_n832), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n827), .A2(G132), .B1(G50), .B2(new_n1129), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n812), .A2(new_n280), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(KEYINPUT123), .B(KEYINPUT53), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n1190), .B(new_n1191), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n824), .A2(G128), .B1(G159), .B2(new_n817), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1189), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n805), .A2(G107), .B1(new_n875), .B2(G97), .ZN(new_n1195));
  OAI221_X1 g0995(.A(new_n1195), .B1(new_n572), .B2(new_n826), .C1(new_n808), .C2(new_n838), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n833), .A2(G294), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n1129), .A2(G68), .B1(new_n817), .B2(G77), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1197), .A2(new_n360), .A3(new_n841), .A4(new_n1198), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n1188), .A2(new_n1194), .B1(new_n1196), .B2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1182), .B1(new_n1200), .B2(new_n801), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n1174), .A2(new_n1046), .B1(new_n1181), .B2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1180), .A2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1203), .A2(KEYINPUT124), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT124), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1180), .A2(new_n1205), .A3(new_n1202), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1204), .A2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(G378));
  NAND4_X1  g1008(.A1(new_n957), .A2(G330), .A3(new_n942), .A4(new_n960), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n954), .A2(new_n952), .A3(new_n955), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT109), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n950), .A2(KEYINPUT109), .A3(new_n952), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n960), .A2(new_n1212), .A3(G330), .A4(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n942), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1209), .A2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n708), .A2(new_n297), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(new_n1218), .B(KEYINPUT55), .ZN(new_n1219));
  XNOR2_X1  g1019(.A(new_n307), .B(new_n1219), .ZN(new_n1220));
  XOR2_X1   g1020(.A(KEYINPUT125), .B(KEYINPUT56), .Z(new_n1221));
  XOR2_X1   g1021(.A(new_n1220), .B(new_n1221), .Z(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1217), .A2(new_n1223), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1209), .A2(new_n1216), .A3(new_n1222), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1224), .A2(new_n1046), .A3(new_n1225), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n789), .B1(new_n870), .B2(G50), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n403), .A2(new_n262), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n245), .A2(new_n262), .ZN(new_n1229));
  AND3_X1   g1029(.A1(new_n1228), .A2(new_n839), .A3(new_n1229), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n806), .A2(new_n223), .B1(new_n352), .B2(new_n821), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(new_n827), .A2(G107), .B1(G58), .B2(new_n1129), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1228), .B1(new_n833), .B2(G283), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n813), .A2(G77), .B1(new_n817), .B2(G68), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1232), .A2(new_n1233), .A3(new_n1234), .ZN(new_n1235));
  AOI211_X1 g1035(.A(new_n1231), .B(new_n1235), .C1(G116), .C2(new_n824), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1230), .B1(new_n1236), .B2(KEYINPUT58), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n827), .A2(G128), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n805), .A2(G132), .B1(G150), .B2(new_n817), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1185), .A2(new_n813), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n824), .A2(G125), .B1(new_n875), .B2(G137), .ZN(new_n1241));
  AND4_X1   g1041(.A1(new_n1238), .A2(new_n1239), .A3(new_n1240), .A4(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1243), .A2(KEYINPUT59), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n810), .A2(new_n389), .ZN(new_n1245));
  AOI211_X1 g1045(.A(new_n1229), .B(new_n1245), .C1(new_n833), .C2(G124), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT59), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1246), .B1(new_n1242), .B2(new_n1247), .ZN(new_n1248));
  OAI221_X1 g1048(.A(new_n1237), .B1(KEYINPUT58), .B2(new_n1236), .C1(new_n1244), .C2(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1227), .B1(new_n1249), .B2(new_n801), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1250), .B1(new_n1222), .B2(new_n794), .ZN(new_n1251));
  AND2_X1   g1051(.A1(new_n1226), .A2(new_n1251), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1169), .B1(new_n1167), .B2(new_n1155), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1253), .A2(new_n1224), .A3(KEYINPUT57), .A4(new_n1225), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1254), .A2(new_n741), .ZN(new_n1255));
  AND3_X1   g1055(.A1(new_n1209), .A2(new_n1216), .A3(new_n1222), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1222), .B1(new_n1209), .B2(new_n1216), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(KEYINPUT57), .B1(new_n1258), .B2(new_n1253), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1252), .B1(new_n1255), .B2(new_n1259), .ZN(G375));
  INV_X1    g1060(.A(new_n1167), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n938), .A2(new_n793), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n789), .B1(new_n871), .B2(G68), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(new_n827), .A2(G137), .B1(G132), .B2(new_n824), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1264), .B1(new_n839), .B2(new_n818), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n833), .A2(G128), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n403), .B1(G58), .B2(new_n1129), .ZN(new_n1267));
  AOI22_X1  g1067(.A1(new_n875), .A2(G150), .B1(new_n813), .B2(G159), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1185), .A2(new_n805), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1266), .A2(new_n1267), .A3(new_n1268), .A4(new_n1269), .ZN(new_n1270));
  AOI22_X1  g1070(.A1(new_n875), .A2(G107), .B1(new_n813), .B2(G97), .ZN(new_n1271));
  OAI221_X1 g1071(.A(new_n1271), .B1(new_n826), .B2(new_n808), .C1(new_n572), .C2(new_n806), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(new_n824), .A2(G294), .B1(new_n353), .B2(new_n817), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n254), .A2(new_n1065), .ZN(new_n1274));
  OAI211_X1 g1074(.A(new_n1273), .B(new_n1274), .C1(new_n587), .C2(new_n832), .ZN(new_n1275));
  OAI22_X1  g1075(.A1(new_n1265), .A2(new_n1270), .B1(new_n1272), .B2(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1263), .B1(new_n1276), .B2(new_n801), .ZN(new_n1277));
  AOI22_X1  g1077(.A1(new_n1261), .A2(new_n1046), .B1(new_n1262), .B2(new_n1277), .ZN(new_n1278));
  AOI211_X1 g1078(.A(new_n1169), .B(new_n1159), .C1(new_n1165), .C2(new_n1166), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1169), .B1(new_n1178), .B2(new_n1159), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1011), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1278), .B1(new_n1279), .B2(new_n1282), .ZN(G381));
  INV_X1    g1083(.A(G375), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1203), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(G384), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(G393), .A2(G396), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1119), .A2(new_n1141), .A3(new_n1287), .A4(new_n1288), .ZN(new_n1289));
  OR4_X1    g1089(.A1(G387), .A2(new_n1286), .A3(new_n1289), .A4(G381), .ZN(G407));
  OAI211_X1 g1090(.A(G407), .B(G213), .C1(G343), .C2(new_n1286), .ZN(G409));
  XNOR2_X1  g1091(.A(G393), .B(G396), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1119), .A2(new_n1141), .A3(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1292), .B1(new_n1119), .B2(new_n1141), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1010), .A2(new_n1006), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1117), .B1(new_n1116), .B2(new_n1042), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1281), .B1(new_n1297), .B2(new_n783), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1046), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1296), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1074), .ZN(new_n1301));
  OAI22_X1  g1101(.A1(new_n1294), .A2(new_n1295), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1292), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(G390), .A2(new_n1303), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1304), .A2(new_n1047), .A3(new_n1074), .A4(new_n1293), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT61), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1302), .A2(new_n1305), .A3(new_n1306), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1279), .B1(KEYINPUT60), .B2(new_n1280), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1167), .A2(KEYINPUT60), .A3(new_n1170), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1309), .A2(new_n741), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1278), .B1(new_n1308), .B2(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1311), .A2(new_n1287), .ZN(new_n1312));
  OAI211_X1 g1112(.A(new_n1278), .B(G384), .C1(new_n1308), .C2(new_n1310), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(new_n701), .A2(G343), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1314), .A2(KEYINPUT126), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1312), .A2(new_n1313), .A3(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1314), .A2(G2897), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1317), .ZN(new_n1319));
  NAND4_X1  g1119(.A1(new_n1312), .A2(new_n1313), .A3(new_n1315), .A4(new_n1319), .ZN(new_n1320));
  AND3_X1   g1120(.A1(new_n1258), .A2(new_n1281), .A3(new_n1253), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1226), .A2(new_n1251), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1285), .B1(new_n1321), .B2(new_n1322), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1323), .B1(new_n1207), .B2(G375), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1314), .ZN(new_n1325));
  AOI22_X1  g1125(.A1(new_n1318), .A2(new_n1320), .B1(new_n1324), .B2(new_n1325), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1307), .B1(new_n1326), .B2(KEYINPUT127), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1328), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1324), .A2(new_n1325), .A3(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT63), .ZN(new_n1331));
  OR2_X1    g1131(.A1(new_n1330), .A2(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1330), .A2(new_n1331), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1318), .A2(new_n1320), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1324), .A2(new_n1325), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT127), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1336), .A2(new_n1337), .ZN(new_n1338));
  NAND4_X1  g1138(.A1(new_n1327), .A2(new_n1332), .A3(new_n1333), .A4(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1330), .A2(KEYINPUT62), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT62), .ZN(new_n1341));
  NAND4_X1  g1141(.A1(new_n1324), .A2(new_n1341), .A3(new_n1325), .A4(new_n1329), .ZN(new_n1342));
  NAND4_X1  g1142(.A1(new_n1340), .A2(new_n1336), .A3(new_n1306), .A4(new_n1342), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1302), .A2(new_n1305), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1343), .A2(new_n1344), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1339), .A2(new_n1345), .ZN(G405));
  NAND2_X1  g1146(.A1(G378), .A2(new_n1284), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(G375), .A2(new_n1285), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1347), .A2(new_n1348), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1349), .A2(new_n1329), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1347), .A2(new_n1328), .A3(new_n1348), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1350), .A2(new_n1351), .ZN(new_n1352));
  XNOR2_X1  g1152(.A(new_n1352), .B(new_n1344), .ZN(G402));
endmodule


