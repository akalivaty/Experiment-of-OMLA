

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768;

  NAND2_X2 U375 ( .A1(n693), .A2(n692), .ZN(n698) );
  OR2_X1 U376 ( .A1(n629), .A2(G902), .ZN(n428) );
  NOR2_X1 U377 ( .A1(n767), .A2(n766), .ZN(n575) );
  XNOR2_X1 U378 ( .A(n461), .B(n460), .ZN(n684) );
  XNOR2_X1 U379 ( .A(n427), .B(n458), .ZN(n714) );
  XNOR2_X1 U380 ( .A(n409), .B(KEYINPUT0), .ZN(n609) );
  INV_X1 U381 ( .A(G953), .ZN(n744) );
  INV_X1 U382 ( .A(n481), .ZN(n587) );
  AND2_X1 U383 ( .A1(n618), .A2(n449), .ZN(n619) );
  NOR2_X1 U384 ( .A1(n573), .A2(n595), .ZN(n565) );
  XOR2_X1 U385 ( .A(n623), .B(KEYINPUT64), .Z(n352) );
  AND2_X1 U386 ( .A1(n356), .A2(n622), .ZN(n353) );
  INV_X2 U387 ( .A(n613), .ZN(n693) );
  XNOR2_X2 U388 ( .A(n545), .B(n544), .ZN(n613) );
  XNOR2_X2 U389 ( .A(n520), .B(n521), .ZN(n546) );
  XNOR2_X2 U390 ( .A(n509), .B(n491), .ZN(n520) );
  XNOR2_X2 U391 ( .A(n583), .B(n582), .ZN(n697) );
  XNOR2_X2 U392 ( .A(n619), .B(KEYINPUT32), .ZN(n765) );
  NOR2_X2 U393 ( .A1(n613), .A2(n612), .ZN(n649) );
  NOR2_X1 U394 ( .A1(n684), .A2(n608), .ZN(n425) );
  NOR2_X1 U395 ( .A1(G902), .A2(n724), .ZN(n554) );
  AND2_X1 U396 ( .A1(n362), .A2(n361), .ZN(n360) );
  NOR2_X1 U397 ( .A1(n714), .A2(n365), .ZN(n596) );
  INV_X1 U398 ( .A(n697), .ZN(n451) );
  XNOR2_X1 U399 ( .A(n428), .B(n373), .ZN(n557) );
  OR2_X1 U400 ( .A1(n355), .A2(n494), .ZN(n495) );
  XNOR2_X1 U401 ( .A(n752), .B(n463), .ZN(n724) );
  INV_X1 U402 ( .A(G122), .ZN(n426) );
  NAND2_X1 U403 ( .A1(n450), .A2(n628), .ZN(n454) );
  AND2_X1 U404 ( .A1(n680), .A2(n494), .ZN(n450) );
  NAND2_X1 U405 ( .A1(n364), .A2(n353), .ZN(n363) );
  NAND2_X1 U406 ( .A1(n360), .A2(n357), .ZN(n364) );
  NAND2_X1 U407 ( .A1(n359), .A2(n358), .ZN(n357) );
  NAND2_X1 U408 ( .A1(n414), .A2(n379), .ZN(n356) );
  AND2_X1 U409 ( .A1(n442), .A2(n368), .ZN(n657) );
  NAND2_X1 U410 ( .A1(n388), .A2(n611), .ZN(n614) );
  XNOR2_X1 U411 ( .A(n609), .B(n366), .ZN(n365) );
  NAND2_X1 U412 ( .A1(n367), .A2(n483), .ZN(n409) );
  AND2_X1 U413 ( .A1(n479), .A2(n386), .ZN(n367) );
  NAND2_X1 U414 ( .A1(n587), .A2(n561), .ZN(n483) );
  XNOR2_X1 U415 ( .A(n747), .B(n485), .ZN(n355) );
  XNOR2_X1 U416 ( .A(n406), .B(n404), .ZN(n747) );
  XNOR2_X1 U417 ( .A(n496), .B(G140), .ZN(n497) );
  XNOR2_X1 U418 ( .A(n426), .B(G107), .ZN(n504) );
  XOR2_X1 U419 ( .A(KEYINPUT70), .B(G137), .Z(n547) );
  XNOR2_X1 U420 ( .A(G125), .B(G146), .ZN(n429) );
  XNOR2_X1 U421 ( .A(G146), .B(G140), .ZN(n550) );
  XOR2_X1 U422 ( .A(G134), .B(G131), .Z(n521) );
  XNOR2_X1 U423 ( .A(n355), .B(n354), .ZN(n637) );
  INV_X1 U424 ( .A(KEYINPUT84), .ZN(n354) );
  INV_X1 U425 ( .A(n649), .ZN(n358) );
  NOR2_X1 U426 ( .A1(n437), .A2(KEYINPUT83), .ZN(n359) );
  NAND2_X1 U427 ( .A1(n437), .A2(KEYINPUT83), .ZN(n361) );
  NAND2_X1 U428 ( .A1(n649), .A2(KEYINPUT83), .ZN(n362) );
  XNOR2_X2 U429 ( .A(n363), .B(n352), .ZN(n675) );
  NOR2_X1 U430 ( .A1(n365), .A2(n615), .ZN(n600) );
  INV_X1 U431 ( .A(KEYINPUT89), .ZN(n366) );
  XNOR2_X1 U432 ( .A(n553), .B(n552), .ZN(n463) );
  AND2_X1 U433 ( .A1(KEYINPUT44), .A2(KEYINPUT67), .ZN(n418) );
  NOR2_X1 U434 ( .A1(n576), .A2(n473), .ZN(n472) );
  XNOR2_X1 U435 ( .A(n513), .B(n462), .ZN(n570) );
  XNOR2_X1 U436 ( .A(G478), .B(KEYINPUT102), .ZN(n462) );
  OR2_X1 U437 ( .A1(n644), .A2(G902), .ZN(n440) );
  XNOR2_X1 U438 ( .A(n543), .B(n372), .ZN(n544) );
  NAND2_X1 U439 ( .A1(n669), .A2(n396), .ZN(n604) );
  NAND2_X1 U440 ( .A1(n620), .A2(n419), .ZN(n417) );
  OR2_X1 U441 ( .A1(n415), .A2(n657), .ZN(n414) );
  INV_X1 U442 ( .A(n547), .ZN(n456) );
  XOR2_X1 U443 ( .A(KEYINPUT91), .B(KEYINPUT90), .Z(n535) );
  XNOR2_X1 U444 ( .A(n520), .B(n486), .ZN(n485) );
  XNOR2_X1 U445 ( .A(n452), .B(n429), .ZN(n486) );
  XNOR2_X1 U446 ( .A(n487), .B(n492), .ZN(n452) );
  XNOR2_X1 U447 ( .A(n394), .B(n387), .ZN(n393) );
  NAND2_X1 U448 ( .A1(n474), .A2(n472), .ZN(n394) );
  XNOR2_X1 U449 ( .A(n584), .B(KEYINPUT108), .ZN(n403) );
  INV_X1 U450 ( .A(KEYINPUT1), .ZN(n580) );
  NAND2_X1 U451 ( .A1(n613), .A2(n430), .ZN(n578) );
  AND2_X1 U452 ( .A1(n446), .A2(n692), .ZN(n430) );
  INV_X1 U453 ( .A(KEYINPUT66), .ZN(n453) );
  NAND2_X1 U454 ( .A1(n465), .A2(n464), .ZN(n589) );
  NAND2_X1 U455 ( .A1(n467), .A2(n466), .ZN(n464) );
  AND2_X1 U456 ( .A1(n469), .A2(n468), .ZN(n465) );
  AND2_X1 U457 ( .A1(n470), .A2(KEYINPUT39), .ZN(n466) );
  NAND2_X1 U458 ( .A1(n557), .A2(n570), .ZN(n396) );
  XNOR2_X1 U459 ( .A(n530), .B(n529), .ZN(n555) );
  XNOR2_X1 U460 ( .A(KEYINPUT107), .B(KEYINPUT30), .ZN(n529) );
  NOR2_X1 U461 ( .A1(n698), .A2(n583), .ZN(n601) );
  XNOR2_X1 U462 ( .A(n615), .B(n420), .ZN(n617) );
  INV_X1 U463 ( .A(KEYINPUT6), .ZN(n420) );
  XNOR2_X1 U464 ( .A(n528), .B(n476), .ZN(n475) );
  XNOR2_X1 U465 ( .A(n527), .B(n369), .ZN(n528) );
  XNOR2_X1 U466 ( .A(n524), .B(n477), .ZN(n476) );
  XNOR2_X1 U467 ( .A(G110), .B(G119), .ZN(n538) );
  XNOR2_X1 U468 ( .A(n389), .B(n510), .ZN(n511) );
  XNOR2_X1 U469 ( .A(n631), .B(n630), .ZN(n632) );
  BUF_X1 U470 ( .A(n728), .Z(n735) );
  AND2_X1 U471 ( .A1(n368), .A2(n418), .ZN(n413) );
  XNOR2_X1 U472 ( .A(n565), .B(n439), .ZN(n438) );
  INV_X1 U473 ( .A(KEYINPUT47), .ZN(n439) );
  XNOR2_X1 U474 ( .A(n488), .B(KEYINPUT17), .ZN(n487) );
  INV_X1 U475 ( .A(KEYINPUT18), .ZN(n488) );
  INV_X1 U476 ( .A(KEYINPUT38), .ZN(n436) );
  NOR2_X1 U477 ( .A1(G953), .A2(G237), .ZN(n526) );
  INV_X1 U478 ( .A(KEYINPUT4), .ZN(n491) );
  XNOR2_X1 U479 ( .A(n435), .B(KEYINPUT97), .ZN(n434) );
  INV_X1 U480 ( .A(KEYINPUT12), .ZN(n435) );
  XNOR2_X1 U481 ( .A(G122), .B(G131), .ZN(n499) );
  NAND2_X1 U482 ( .A1(G237), .A2(G234), .ZN(n514) );
  OR2_X1 U483 ( .A1(G902), .A2(G237), .ZN(n519) );
  INV_X1 U484 ( .A(KEYINPUT103), .ZN(n460) );
  AND2_X1 U485 ( .A1(n682), .A2(n446), .ZN(n470) );
  OR2_X1 U486 ( .A1(n470), .A2(KEYINPUT39), .ZN(n468) );
  XNOR2_X1 U487 ( .A(n525), .B(KEYINPUT95), .ZN(n477) );
  XNOR2_X1 U488 ( .A(G113), .B(G101), .ZN(n525) );
  XNOR2_X1 U489 ( .A(n478), .B(G104), .ZN(n498) );
  INV_X1 U490 ( .A(G113), .ZN(n478) );
  XNOR2_X1 U491 ( .A(n407), .B(G119), .ZN(n527) );
  XNOR2_X1 U492 ( .A(G116), .B(KEYINPUT3), .ZN(n407) );
  XOR2_X1 U493 ( .A(KEYINPUT16), .B(KEYINPUT71), .Z(n493) );
  XNOR2_X1 U494 ( .A(n448), .B(n536), .ZN(n455) );
  XNOR2_X1 U495 ( .A(n456), .B(n535), .ZN(n448) );
  XNOR2_X1 U496 ( .A(n509), .B(n370), .ZN(n389) );
  XNOR2_X1 U497 ( .A(n432), .B(KEYINPUT99), .ZN(n431) );
  INV_X1 U498 ( .A(KEYINPUT7), .ZN(n432) );
  XNOR2_X1 U499 ( .A(n546), .B(n547), .ZN(n752) );
  XOR2_X1 U500 ( .A(G107), .B(G104), .Z(n549) );
  XNOR2_X1 U501 ( .A(n405), .B(G110), .ZN(n553) );
  XNOR2_X1 U502 ( .A(G101), .B(KEYINPUT87), .ZN(n405) );
  NAND2_X1 U503 ( .A1(n393), .A2(n380), .ZN(n590) );
  AND2_X1 U504 ( .A1(n393), .A2(n375), .ZN(n755) );
  NOR2_X1 U505 ( .A1(n696), .A2(n578), .ZN(n563) );
  XNOR2_X1 U506 ( .A(n614), .B(KEYINPUT105), .ZN(n442) );
  XNOR2_X1 U507 ( .A(n553), .B(n498), .ZN(n404) );
  XNOR2_X1 U508 ( .A(n408), .B(n527), .ZN(n406) );
  XNOR2_X1 U509 ( .A(n504), .B(n493), .ZN(n408) );
  XNOR2_X1 U510 ( .A(n637), .B(n636), .ZN(n638) );
  NOR2_X1 U511 ( .A1(n589), .A2(n396), .ZN(n569) );
  NAND2_X1 U512 ( .A1(n398), .A2(n397), .ZN(n672) );
  AND2_X1 U513 ( .A1(n399), .A2(n384), .ZN(n398) );
  NAND2_X1 U514 ( .A1(n402), .A2(n401), .ZN(n397) );
  NOR2_X1 U515 ( .A1(n617), .A2(n693), .ZN(n449) );
  XNOR2_X1 U516 ( .A(n396), .B(n395), .ZN(n664) );
  INV_X1 U517 ( .A(KEYINPUT106), .ZN(n395) );
  AND2_X1 U518 ( .A1(n568), .A2(n381), .ZN(n662) );
  XNOR2_X1 U519 ( .A(n392), .B(n391), .ZN(n612) );
  INV_X1 U520 ( .A(KEYINPUT82), .ZN(n391) );
  NOR2_X1 U521 ( .A1(n614), .A2(n617), .ZN(n392) );
  XNOR2_X1 U522 ( .A(n644), .B(n643), .ZN(n645) );
  XNOR2_X1 U523 ( .A(n736), .B(n737), .ZN(n422) );
  INV_X1 U524 ( .A(n729), .ZN(n730) );
  INV_X1 U525 ( .A(KEYINPUT60), .ZN(n423) );
  INV_X1 U526 ( .A(n587), .ZN(n433) );
  BUF_X1 U527 ( .A(n697), .Z(n388) );
  NOR2_X1 U528 ( .A1(n693), .A2(n615), .ZN(n368) );
  AND2_X1 U529 ( .A1(G210), .A2(n526), .ZN(n369) );
  XNOR2_X1 U530 ( .A(KEYINPUT100), .B(KEYINPUT101), .ZN(n370) );
  INV_X1 U531 ( .A(n562), .ZN(n446) );
  XOR2_X1 U532 ( .A(n594), .B(KEYINPUT88), .Z(n371) );
  XNOR2_X1 U533 ( .A(KEYINPUT25), .B(KEYINPUT75), .ZN(n372) );
  XOR2_X1 U534 ( .A(n503), .B(G475), .Z(n373) );
  XOR2_X1 U535 ( .A(G143), .B(KEYINPUT11), .Z(n374) );
  AND2_X1 U536 ( .A1(n674), .A2(n673), .ZN(n375) );
  NOR2_X1 U537 ( .A1(n697), .A2(n698), .ZN(n376) );
  AND2_X1 U538 ( .A1(n457), .A2(n617), .ZN(n377) );
  NOR2_X1 U539 ( .A1(n657), .A2(n765), .ZN(n378) );
  AND2_X1 U540 ( .A1(n411), .A2(n410), .ZN(n379) );
  AND2_X1 U541 ( .A1(n375), .A2(KEYINPUT2), .ZN(n380) );
  AND2_X1 U542 ( .A1(n597), .A2(n433), .ZN(n381) );
  AND2_X1 U543 ( .A1(n519), .A2(G210), .ZN(n382) );
  XOR2_X1 U544 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n383) );
  INV_X1 U545 ( .A(n429), .ZN(n496) );
  AND2_X1 U546 ( .A1(n451), .A2(n400), .ZN(n384) );
  AND2_X1 U547 ( .A1(n483), .A2(n482), .ZN(n385) );
  AND2_X1 U548 ( .A1(n482), .A2(n371), .ZN(n386) );
  INV_X1 U549 ( .A(KEYINPUT39), .ZN(n471) );
  INV_X1 U550 ( .A(n681), .ZN(n484) );
  XNOR2_X1 U551 ( .A(KEYINPUT48), .B(KEYINPUT81), .ZN(n387) );
  INV_X1 U552 ( .A(KEYINPUT67), .ZN(n419) );
  XNOR2_X1 U553 ( .A(G902), .B(KEYINPUT15), .ZN(n625) );
  XNOR2_X1 U554 ( .A(n434), .B(n374), .ZN(n443) );
  NAND2_X1 U555 ( .A1(n451), .A2(n377), .ZN(n427) );
  XNOR2_X1 U556 ( .A(n443), .B(n501), .ZN(n441) );
  XNOR2_X1 U557 ( .A(n390), .B(KEYINPUT22), .ZN(n616) );
  NAND2_X1 U558 ( .A1(n459), .A2(n610), .ZN(n390) );
  INV_X1 U559 ( .A(n403), .ZN(n402) );
  NAND2_X1 U560 ( .A1(n403), .A2(KEYINPUT36), .ZN(n399) );
  NAND2_X1 U561 ( .A1(n579), .A2(KEYINPUT36), .ZN(n400) );
  NOR2_X1 U562 ( .A1(n579), .A2(KEYINPUT36), .ZN(n401) );
  NAND2_X1 U563 ( .A1(n481), .A2(n480), .ZN(n479) );
  NAND2_X1 U564 ( .A1(n765), .A2(n418), .ZN(n410) );
  AND2_X1 U565 ( .A1(n412), .A2(n417), .ZN(n411) );
  NAND2_X1 U566 ( .A1(n442), .A2(n413), .ZN(n412) );
  NAND2_X1 U567 ( .A1(n416), .A2(n419), .ZN(n415) );
  INV_X1 U568 ( .A(n765), .ZN(n416) );
  NAND2_X1 U569 ( .A1(n728), .A2(G478), .ZN(n731) );
  XNOR2_X2 U570 ( .A(n454), .B(n453), .ZN(n728) );
  NAND2_X1 U571 ( .A1(n728), .A2(G210), .ZN(n639) );
  XNOR2_X1 U572 ( .A(n421), .B(n642), .ZN(G51) );
  NAND2_X1 U573 ( .A1(n640), .A2(n732), .ZN(n421) );
  NOR2_X1 U574 ( .A1(n422), .A2(n738), .ZN(G66) );
  XNOR2_X1 U575 ( .A(n424), .B(n423), .ZN(G60) );
  NAND2_X1 U576 ( .A1(n635), .A2(n732), .ZN(n424) );
  XNOR2_X1 U577 ( .A(n441), .B(n500), .ZN(n502) );
  XNOR2_X1 U578 ( .A(n425), .B(KEYINPUT104), .ZN(n459) );
  XNOR2_X1 U579 ( .A(n508), .B(n431), .ZN(n510) );
  NAND2_X1 U580 ( .A1(n675), .A2(n624), .ZN(n680) );
  NOR2_X1 U581 ( .A1(G902), .A2(n737), .ZN(n545) );
  INV_X1 U582 ( .A(n698), .ZN(n457) );
  NAND2_X1 U583 ( .A1(n682), .A2(n681), .ZN(n685) );
  XNOR2_X1 U584 ( .A(n481), .B(n436), .ZN(n682) );
  NAND2_X1 U585 ( .A1(n607), .A2(n606), .ZN(n437) );
  NAND2_X1 U586 ( .A1(n566), .A2(n438), .ZN(n445) );
  XNOR2_X1 U587 ( .A(n511), .B(n512), .ZN(n729) );
  XNOR2_X2 U588 ( .A(n440), .B(G472), .ZN(n615) );
  XNOR2_X1 U589 ( .A(n498), .B(n499), .ZN(n500) );
  XNOR2_X2 U590 ( .A(n554), .B(G469), .ZN(n583) );
  NAND2_X1 U591 ( .A1(n444), .A2(n564), .ZN(n573) );
  XNOR2_X1 U592 ( .A(n563), .B(KEYINPUT28), .ZN(n444) );
  NAND2_X1 U593 ( .A1(n445), .A2(n567), .ZN(n447) );
  XNOR2_X1 U594 ( .A(n575), .B(KEYINPUT46), .ZN(n474) );
  XNOR2_X1 U595 ( .A(n447), .B(KEYINPUT72), .ZN(n576) );
  NAND2_X1 U596 ( .A1(n571), .A2(n570), .ZN(n461) );
  XNOR2_X1 U597 ( .A(n753), .B(n455), .ZN(n541) );
  NAND2_X1 U598 ( .A1(n675), .A2(n755), .ZN(n627) );
  XNOR2_X1 U599 ( .A(n546), .B(n475), .ZN(n644) );
  XNOR2_X2 U600 ( .A(n495), .B(n382), .ZN(n481) );
  INV_X1 U601 ( .A(KEYINPUT33), .ZN(n458) );
  INV_X1 U602 ( .A(n556), .ZN(n467) );
  NAND2_X1 U603 ( .A1(n556), .A2(n471), .ZN(n469) );
  NOR2_X1 U604 ( .A1(n556), .A2(n562), .ZN(n568) );
  INV_X1 U605 ( .A(n672), .ZN(n473) );
  NAND2_X1 U606 ( .A1(n385), .A2(n479), .ZN(n595) );
  NAND2_X1 U607 ( .A1(n433), .A2(n681), .ZN(n579) );
  NOR2_X1 U608 ( .A1(n484), .A2(n561), .ZN(n480) );
  NAND2_X1 U609 ( .A1(n484), .A2(n561), .ZN(n482) );
  XNOR2_X1 U610 ( .A(n726), .B(n725), .ZN(n727) );
  XNOR2_X1 U611 ( .A(n724), .B(n489), .ZN(n725) );
  BUF_X1 U612 ( .A(n675), .Z(n743) );
  XNOR2_X2 U613 ( .A(n490), .B(G143), .ZN(n509) );
  XNOR2_X2 U614 ( .A(G128), .B(KEYINPUT65), .ZN(n490) );
  XNOR2_X2 U615 ( .A(n497), .B(KEYINPUT10), .ZN(n753) );
  XOR2_X1 U616 ( .A(n723), .B(n722), .Z(n489) );
  INV_X1 U617 ( .A(KEYINPUT62), .ZN(n643) );
  XNOR2_X1 U618 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U619 ( .A(n646), .B(n645), .ZN(n647) );
  XNOR2_X1 U620 ( .A(n639), .B(n638), .ZN(n640) );
  NAND2_X1 U621 ( .A1(G224), .A2(n744), .ZN(n492) );
  INV_X1 U622 ( .A(n625), .ZN(n494) );
  NAND2_X1 U623 ( .A1(n526), .A2(G214), .ZN(n501) );
  XNOR2_X1 U624 ( .A(n502), .B(n753), .ZN(n629) );
  XNOR2_X1 U625 ( .A(KEYINPUT13), .B(KEYINPUT98), .ZN(n503) );
  INV_X1 U626 ( .A(n557), .ZN(n571) );
  XOR2_X1 U627 ( .A(n504), .B(KEYINPUT9), .Z(n507) );
  NAND2_X1 U628 ( .A1(G234), .A2(n744), .ZN(n505) );
  XOR2_X1 U629 ( .A(KEYINPUT8), .B(n505), .Z(n537) );
  NAND2_X1 U630 ( .A1(G217), .A2(n537), .ZN(n506) );
  XNOR2_X1 U631 ( .A(n507), .B(n506), .ZN(n512) );
  XNOR2_X1 U632 ( .A(G116), .B(G134), .ZN(n508) );
  NOR2_X1 U633 ( .A1(n729), .A2(G902), .ZN(n513) );
  NOR2_X1 U634 ( .A1(n571), .A2(n570), .ZN(n597) );
  XOR2_X1 U635 ( .A(KEYINPUT73), .B(KEYINPUT14), .Z(n515) );
  XNOR2_X1 U636 ( .A(n515), .B(n514), .ZN(n516) );
  NAND2_X1 U637 ( .A1(G952), .A2(n516), .ZN(n713) );
  NOR2_X1 U638 ( .A1(G953), .A2(n713), .ZN(n593) );
  NAND2_X1 U639 ( .A1(G902), .A2(n516), .ZN(n591) );
  OR2_X1 U640 ( .A1(n744), .A2(n591), .ZN(n517) );
  NOR2_X1 U641 ( .A1(G900), .A2(n517), .ZN(n518) );
  NOR2_X1 U642 ( .A1(n593), .A2(n518), .ZN(n562) );
  NAND2_X1 U643 ( .A1(G214), .A2(n519), .ZN(n681) );
  XOR2_X1 U644 ( .A(KEYINPUT94), .B(KEYINPUT5), .Z(n523) );
  XNOR2_X1 U645 ( .A(G146), .B(G137), .ZN(n522) );
  XNOR2_X1 U646 ( .A(n523), .B(n522), .ZN(n524) );
  NAND2_X1 U647 ( .A1(n681), .A2(n615), .ZN(n530) );
  XOR2_X1 U648 ( .A(KEYINPUT20), .B(KEYINPUT93), .Z(n532) );
  NAND2_X1 U649 ( .A1(G234), .A2(n625), .ZN(n531) );
  XNOR2_X1 U650 ( .A(n532), .B(n531), .ZN(n542) );
  NAND2_X1 U651 ( .A1(G221), .A2(n542), .ZN(n533) );
  XNOR2_X1 U652 ( .A(KEYINPUT21), .B(n533), .ZN(n608) );
  INV_X1 U653 ( .A(n608), .ZN(n692) );
  XNOR2_X1 U654 ( .A(G128), .B(KEYINPUT92), .ZN(n534) );
  XNOR2_X1 U655 ( .A(n383), .B(n534), .ZN(n536) );
  NAND2_X1 U656 ( .A1(n537), .A2(G221), .ZN(n539) );
  XNOR2_X1 U657 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U658 ( .A(n541), .B(n540), .ZN(n737) );
  NAND2_X1 U659 ( .A1(n542), .A2(G217), .ZN(n543) );
  NAND2_X1 U660 ( .A1(G227), .A2(n744), .ZN(n548) );
  XOR2_X1 U661 ( .A(n549), .B(n548), .Z(n551) );
  XNOR2_X1 U662 ( .A(n551), .B(n550), .ZN(n552) );
  NAND2_X1 U663 ( .A1(n555), .A2(n601), .ZN(n556) );
  NOR2_X1 U664 ( .A1(n570), .A2(n557), .ZN(n659) );
  INV_X1 U665 ( .A(n659), .ZN(n669) );
  INV_X1 U666 ( .A(n604), .ZN(n686) );
  NAND2_X1 U667 ( .A1(n686), .A2(KEYINPUT47), .ZN(n558) );
  XNOR2_X1 U668 ( .A(KEYINPUT77), .B(n558), .ZN(n559) );
  NOR2_X1 U669 ( .A1(n662), .A2(n559), .ZN(n560) );
  XNOR2_X1 U670 ( .A(n560), .B(KEYINPUT76), .ZN(n567) );
  XOR2_X1 U671 ( .A(KEYINPUT74), .B(KEYINPUT19), .Z(n561) );
  INV_X1 U672 ( .A(n615), .ZN(n696) );
  INV_X1 U673 ( .A(n583), .ZN(n564) );
  NAND2_X1 U674 ( .A1(n565), .A2(n686), .ZN(n566) );
  XNOR2_X1 U675 ( .A(n569), .B(KEYINPUT40), .ZN(n767) );
  NOR2_X1 U676 ( .A1(n685), .A2(n684), .ZN(n572) );
  XNOR2_X1 U677 ( .A(n572), .B(KEYINPUT41), .ZN(n715) );
  NOR2_X1 U678 ( .A1(n715), .A2(n573), .ZN(n574) );
  XNOR2_X1 U679 ( .A(n574), .B(KEYINPUT42), .ZN(n766) );
  NAND2_X1 U680 ( .A1(n617), .A2(n664), .ZN(n577) );
  OR2_X1 U681 ( .A1(n578), .A2(n577), .ZN(n584) );
  INV_X1 U682 ( .A(KEYINPUT68), .ZN(n581) );
  NOR2_X1 U683 ( .A1(n451), .A2(n584), .ZN(n585) );
  NAND2_X1 U684 ( .A1(n585), .A2(n681), .ZN(n586) );
  XNOR2_X1 U685 ( .A(KEYINPUT43), .B(n586), .ZN(n588) );
  NAND2_X1 U686 ( .A1(n588), .A2(n587), .ZN(n674) );
  OR2_X1 U687 ( .A1(n669), .A2(n589), .ZN(n673) );
  XNOR2_X1 U688 ( .A(n590), .B(KEYINPUT79), .ZN(n624) );
  OR2_X1 U689 ( .A1(n744), .A2(G898), .ZN(n749) );
  NOR2_X1 U690 ( .A1(n749), .A2(n591), .ZN(n592) );
  NOR2_X1 U691 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U692 ( .A(n596), .B(KEYINPUT34), .ZN(n598) );
  NAND2_X1 U693 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X2 U694 ( .A(n599), .B(KEYINPUT35), .ZN(n763) );
  NAND2_X1 U695 ( .A1(n763), .A2(KEYINPUT44), .ZN(n607) );
  NAND2_X1 U696 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U697 ( .A(KEYINPUT96), .B(n602), .ZN(n654) );
  NAND2_X1 U698 ( .A1(n615), .A2(n376), .ZN(n703) );
  NOR2_X1 U699 ( .A1(n609), .A2(n703), .ZN(n603) );
  XNOR2_X1 U700 ( .A(KEYINPUT31), .B(n603), .ZN(n668) );
  NAND2_X1 U701 ( .A1(n654), .A2(n668), .ZN(n605) );
  NAND2_X1 U702 ( .A1(n605), .A2(n604), .ZN(n606) );
  INV_X1 U703 ( .A(n609), .ZN(n610) );
  INV_X1 U704 ( .A(n616), .ZN(n611) );
  NOR2_X1 U705 ( .A1(n616), .A2(n388), .ZN(n618) );
  INV_X1 U706 ( .A(KEYINPUT44), .ZN(n620) );
  NOR2_X1 U707 ( .A1(n763), .A2(KEYINPUT44), .ZN(n621) );
  NAND2_X1 U708 ( .A1(n378), .A2(n621), .ZN(n622) );
  INV_X1 U709 ( .A(KEYINPUT45), .ZN(n623) );
  INV_X1 U710 ( .A(KEYINPUT2), .ZN(n626) );
  NAND2_X1 U711 ( .A1(n627), .A2(n626), .ZN(n628) );
  NAND2_X1 U712 ( .A1(n728), .A2(G475), .ZN(n633) );
  XNOR2_X1 U713 ( .A(KEYINPUT69), .B(KEYINPUT85), .ZN(n631) );
  XNOR2_X1 U714 ( .A(n629), .B(KEYINPUT59), .ZN(n630) );
  XNOR2_X1 U715 ( .A(n633), .B(n632), .ZN(n635) );
  NOR2_X1 U716 ( .A1(G952), .A2(n744), .ZN(n634) );
  XNOR2_X1 U717 ( .A(KEYINPUT86), .B(n634), .ZN(n738) );
  INV_X1 U718 ( .A(n738), .ZN(n732) );
  XOR2_X1 U719 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n636) );
  XOR2_X1 U720 ( .A(KEYINPUT80), .B(KEYINPUT118), .Z(n641) );
  XNOR2_X1 U721 ( .A(n641), .B(KEYINPUT56), .ZN(n642) );
  NAND2_X1 U722 ( .A1(n728), .A2(G472), .ZN(n646) );
  NAND2_X1 U723 ( .A1(n647), .A2(n732), .ZN(n648) );
  XNOR2_X1 U724 ( .A(n648), .B(KEYINPUT63), .ZN(G57) );
  XOR2_X1 U725 ( .A(n649), .B(G101), .Z(G3) );
  XNOR2_X1 U726 ( .A(G104), .B(KEYINPUT109), .ZN(n651) );
  INV_X1 U727 ( .A(n664), .ZN(n666) );
  NOR2_X1 U728 ( .A1(n654), .A2(n666), .ZN(n650) );
  XNOR2_X1 U729 ( .A(n651), .B(n650), .ZN(G6) );
  XOR2_X1 U730 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n653) );
  XNOR2_X1 U731 ( .A(G107), .B(KEYINPUT110), .ZN(n652) );
  XNOR2_X1 U732 ( .A(n653), .B(n652), .ZN(n656) );
  NOR2_X1 U733 ( .A1(n654), .A2(n669), .ZN(n655) );
  XOR2_X1 U734 ( .A(n656), .B(n655), .Z(G9) );
  XNOR2_X1 U735 ( .A(n657), .B(G110), .ZN(n658) );
  XNOR2_X1 U736 ( .A(n658), .B(KEYINPUT111), .ZN(G12) );
  XOR2_X1 U737 ( .A(G128), .B(KEYINPUT29), .Z(n661) );
  NAND2_X1 U738 ( .A1(n565), .A2(n659), .ZN(n660) );
  XNOR2_X1 U739 ( .A(n661), .B(n660), .ZN(G30) );
  XOR2_X1 U740 ( .A(n662), .B(G143), .Z(n663) );
  XNOR2_X1 U741 ( .A(KEYINPUT112), .B(n663), .ZN(G45) );
  NAND2_X1 U742 ( .A1(n664), .A2(n565), .ZN(n665) );
  XNOR2_X1 U743 ( .A(n665), .B(G146), .ZN(G48) );
  NOR2_X1 U744 ( .A1(n666), .A2(n668), .ZN(n667) );
  XOR2_X1 U745 ( .A(G113), .B(n667), .Z(G15) );
  NOR2_X1 U746 ( .A1(n669), .A2(n668), .ZN(n670) );
  XOR2_X1 U747 ( .A(G116), .B(n670), .Z(G18) );
  XOR2_X1 U748 ( .A(G125), .B(KEYINPUT37), .Z(n671) );
  XNOR2_X1 U749 ( .A(n672), .B(n671), .ZN(G27) );
  XNOR2_X1 U750 ( .A(G134), .B(n673), .ZN(G36) );
  XNOR2_X1 U751 ( .A(G140), .B(n674), .ZN(G42) );
  NOR2_X1 U752 ( .A1(KEYINPUT2), .A2(n743), .ZN(n676) );
  XNOR2_X1 U753 ( .A(n676), .B(KEYINPUT78), .ZN(n678) );
  NOR2_X1 U754 ( .A1(n755), .A2(KEYINPUT2), .ZN(n677) );
  NOR2_X1 U755 ( .A1(n678), .A2(n677), .ZN(n679) );
  NAND2_X1 U756 ( .A1(n680), .A2(n679), .ZN(n719) );
  NOR2_X1 U757 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U758 ( .A1(n684), .A2(n683), .ZN(n689) );
  NOR2_X1 U759 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U760 ( .A(n687), .B(KEYINPUT116), .ZN(n688) );
  NOR2_X1 U761 ( .A1(n689), .A2(n688), .ZN(n690) );
  XOR2_X1 U762 ( .A(KEYINPUT117), .B(n690), .Z(n691) );
  NOR2_X1 U763 ( .A1(n714), .A2(n691), .ZN(n710) );
  NOR2_X1 U764 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U765 ( .A(n694), .B(KEYINPUT49), .ZN(n695) );
  NAND2_X1 U766 ( .A1(n696), .A2(n695), .ZN(n701) );
  NAND2_X1 U767 ( .A1(n698), .A2(n388), .ZN(n699) );
  XOR2_X1 U768 ( .A(KEYINPUT50), .B(n699), .Z(n700) );
  NOR2_X1 U769 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U770 ( .A(KEYINPUT113), .B(n702), .ZN(n704) );
  NAND2_X1 U771 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U772 ( .A(n705), .B(KEYINPUT115), .ZN(n707) );
  XOR2_X1 U773 ( .A(KEYINPUT51), .B(KEYINPUT114), .Z(n706) );
  XNOR2_X1 U774 ( .A(n707), .B(n706), .ZN(n708) );
  NOR2_X1 U775 ( .A1(n715), .A2(n708), .ZN(n709) );
  NOR2_X1 U776 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U777 ( .A(n711), .B(KEYINPUT52), .ZN(n712) );
  NOR2_X1 U778 ( .A1(n713), .A2(n712), .ZN(n717) );
  NOR2_X1 U779 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U780 ( .A1(n717), .A2(n716), .ZN(n718) );
  NAND2_X1 U781 ( .A1(n719), .A2(n718), .ZN(n720) );
  NOR2_X1 U782 ( .A1(n720), .A2(G953), .ZN(n721) );
  XNOR2_X1 U783 ( .A(n721), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U784 ( .A1(n735), .A2(G469), .ZN(n726) );
  XOR2_X1 U785 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n723) );
  XNOR2_X1 U786 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n722) );
  NOR2_X1 U787 ( .A1(n738), .A2(n727), .ZN(G54) );
  XNOR2_X1 U788 ( .A(n731), .B(n730), .ZN(n733) );
  NAND2_X1 U789 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U790 ( .A(n734), .B(KEYINPUT121), .ZN(G63) );
  NAND2_X1 U791 ( .A1(G217), .A2(n735), .ZN(n736) );
  XOR2_X1 U792 ( .A(KEYINPUT61), .B(KEYINPUT123), .Z(n740) );
  NAND2_X1 U793 ( .A1(G224), .A2(G953), .ZN(n739) );
  XNOR2_X1 U794 ( .A(n740), .B(n739), .ZN(n741) );
  XNOR2_X1 U795 ( .A(KEYINPUT122), .B(n741), .ZN(n742) );
  NAND2_X1 U796 ( .A1(n742), .A2(G898), .ZN(n746) );
  NAND2_X1 U797 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U798 ( .A1(n746), .A2(n745), .ZN(n751) );
  XNOR2_X1 U799 ( .A(n747), .B(KEYINPUT124), .ZN(n748) );
  NAND2_X1 U800 ( .A1(n749), .A2(n748), .ZN(n750) );
  XOR2_X1 U801 ( .A(n751), .B(n750), .Z(G69) );
  XOR2_X1 U802 ( .A(n752), .B(n753), .Z(n758) );
  INV_X1 U803 ( .A(n758), .ZN(n754) );
  XNOR2_X1 U804 ( .A(n755), .B(n754), .ZN(n756) );
  NOR2_X1 U805 ( .A1(G953), .A2(n756), .ZN(n757) );
  XNOR2_X1 U806 ( .A(KEYINPUT125), .B(n757), .ZN(n762) );
  XOR2_X1 U807 ( .A(G227), .B(n758), .Z(n759) );
  NAND2_X1 U808 ( .A1(n759), .A2(G900), .ZN(n760) );
  NAND2_X1 U809 ( .A1(n760), .A2(G953), .ZN(n761) );
  NAND2_X1 U810 ( .A1(n762), .A2(n761), .ZN(G72) );
  XOR2_X1 U811 ( .A(n763), .B(G122), .Z(G24) );
  XOR2_X1 U812 ( .A(G119), .B(KEYINPUT126), .Z(n764) );
  XNOR2_X1 U813 ( .A(n765), .B(n764), .ZN(G21) );
  XOR2_X1 U814 ( .A(n766), .B(G137), .Z(G39) );
  XNOR2_X1 U815 ( .A(G131), .B(KEYINPUT127), .ZN(n768) );
  XNOR2_X1 U816 ( .A(n768), .B(n767), .ZN(G33) );
endmodule

