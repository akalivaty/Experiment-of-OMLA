//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 1 0 0 0 1 0 1 1 1 1 0 0 1 1 0 0 1 0 0 1 0 1 0 1 1 0 1 1 0 0 0 1 1 0 0 0 1 1 1 0 1 0 1 1 1 1 1 1 1 0 0 1 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:11 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n603, new_n604, new_n605, new_n606, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n616, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n674, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n887, new_n888, new_n889, new_n890, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951;
  INV_X1    g000(.A(G237), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n187), .A2(new_n188), .A3(G210), .ZN(new_n189));
  INV_X1    g003(.A(G101), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n192));
  XOR2_X1   g006(.A(new_n191), .B(new_n192), .Z(new_n193));
  INV_X1    g007(.A(KEYINPUT11), .ZN(new_n194));
  INV_X1    g008(.A(G134), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n194), .B1(new_n195), .B2(G137), .ZN(new_n196));
  INV_X1    g010(.A(G137), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n197), .A2(KEYINPUT11), .A3(G134), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n195), .A2(G137), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n196), .A2(new_n198), .A3(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(KEYINPUT68), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT68), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n196), .A2(new_n198), .A3(new_n202), .A4(new_n199), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n201), .A2(G131), .A3(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT69), .ZN(new_n205));
  AND3_X1   g019(.A1(new_n196), .A2(new_n198), .A3(new_n199), .ZN(new_n206));
  INV_X1    g020(.A(G131), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n204), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G143), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(KEYINPUT66), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT66), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G143), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G146), .ZN(new_n215));
  AND2_X1   g029(.A1(KEYINPUT67), .A2(G146), .ZN(new_n216));
  NOR2_X1   g030(.A1(KEYINPUT67), .A2(G146), .ZN(new_n217));
  OAI21_X1  g031(.A(G143), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n215), .A2(KEYINPUT0), .A3(G128), .A4(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(KEYINPUT0), .A2(G128), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT0), .ZN(new_n221));
  INV_X1    g035(.A(G128), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n221), .A2(new_n222), .A3(KEYINPUT65), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT65), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n224), .B1(KEYINPUT0), .B2(G128), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G146), .ZN(new_n227));
  AND3_X1   g041(.A1(new_n211), .A2(new_n213), .A3(new_n227), .ZN(new_n228));
  NOR3_X1   g042(.A1(new_n216), .A2(new_n217), .A3(G143), .ZN(new_n229));
  OAI211_X1 g043(.A(new_n220), .B(new_n226), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n201), .A2(new_n205), .A3(G131), .A4(new_n203), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n209), .A2(new_n219), .A3(new_n230), .A4(new_n231), .ZN(new_n232));
  XNOR2_X1  g046(.A(KEYINPUT71), .B(G116), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G119), .ZN(new_n234));
  INV_X1    g048(.A(G116), .ZN(new_n235));
  OAI21_X1  g049(.A(KEYINPUT70), .B1(new_n235), .B2(G119), .ZN(new_n236));
  OR3_X1    g050(.A1(new_n235), .A2(KEYINPUT70), .A3(G119), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n234), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  XNOR2_X1  g052(.A(KEYINPUT2), .B(G113), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n239), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n234), .A2(new_n241), .A3(new_n236), .A4(new_n237), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT1), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n215), .A2(new_n245), .A3(G128), .A4(new_n218), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n228), .A2(new_n229), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n222), .B1(new_n218), .B2(KEYINPUT1), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n246), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n206), .A2(new_n207), .ZN(new_n250));
  INV_X1    g064(.A(new_n199), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n195), .A2(G137), .ZN(new_n252));
  OAI21_X1  g066(.A(G131), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n249), .A2(new_n250), .A3(new_n253), .ZN(new_n254));
  AND3_X1   g068(.A1(new_n232), .A2(new_n244), .A3(new_n254), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n244), .B1(new_n232), .B2(new_n254), .ZN(new_n256));
  OAI21_X1  g070(.A(KEYINPUT28), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n232), .A2(new_n244), .A3(new_n254), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT28), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(KEYINPUT72), .B1(new_n257), .B2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT72), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n232), .A2(new_n254), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(new_n243), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(new_n258), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n262), .B1(new_n265), .B2(KEYINPUT28), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n193), .B1(new_n261), .B2(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(KEYINPUT30), .B1(new_n263), .B2(KEYINPUT64), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT64), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT30), .ZN(new_n270));
  AOI211_X1 g084(.A(new_n269), .B(new_n270), .C1(new_n232), .C2(new_n254), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n243), .B1(new_n268), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n193), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n272), .A2(new_n258), .A3(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(KEYINPUT29), .B1(new_n267), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G902), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n257), .A2(new_n260), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n193), .A2(KEYINPUT29), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n276), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(G472), .B1(new_n275), .B2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT73), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n272), .A2(new_n258), .A3(new_n193), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(KEYINPUT31), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n273), .B1(new_n261), .B2(new_n266), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT31), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n272), .A2(new_n286), .A3(new_n258), .A4(new_n193), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n284), .A2(new_n285), .A3(new_n287), .ZN(new_n288));
  NOR2_X1   g102(.A1(G472), .A2(G902), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT32), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  OAI211_X1 g106(.A(KEYINPUT73), .B(G472), .C1(new_n275), .C2(new_n279), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n282), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n288), .A2(KEYINPUT32), .A3(new_n289), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(KEYINPUT74), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT74), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n288), .A2(new_n297), .A3(KEYINPUT32), .A4(new_n289), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  OR2_X1    g113(.A1(new_n294), .A2(new_n299), .ZN(new_n300));
  XNOR2_X1  g114(.A(KEYINPUT9), .B(G234), .ZN(new_n301));
  XNOR2_X1  g115(.A(new_n301), .B(KEYINPUT79), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(new_n276), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(G221), .ZN(new_n304));
  XOR2_X1   g118(.A(new_n304), .B(KEYINPUT80), .Z(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  XOR2_X1   g120(.A(G110), .B(G140), .Z(new_n307));
  INV_X1    g121(.A(G227), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n308), .A2(G953), .ZN(new_n309));
  XNOR2_X1  g123(.A(new_n307), .B(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G104), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G107), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(KEYINPUT83), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT83), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n315), .A2(new_n312), .A3(G107), .ZN(new_n316));
  INV_X1    g130(.A(G107), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G104), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n314), .A2(new_n316), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G101), .ZN(new_n320));
  AND3_X1   g134(.A1(new_n317), .A2(KEYINPUT3), .A3(G104), .ZN(new_n321));
  AOI21_X1  g135(.A(KEYINPUT3), .B1(new_n317), .B2(G104), .ZN(new_n322));
  OAI211_X1 g136(.A(new_n190), .B(new_n313), .C1(new_n321), .C2(new_n322), .ZN(new_n323));
  AND2_X1   g137(.A1(new_n320), .A2(new_n323), .ZN(new_n324));
  AND3_X1   g138(.A1(new_n249), .A2(new_n324), .A3(KEYINPUT10), .ZN(new_n325));
  XNOR2_X1  g139(.A(KEYINPUT67), .B(G146), .ZN(new_n326));
  AOI22_X1  g140(.A1(G146), .A2(new_n214), .B1(new_n326), .B2(G143), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n211), .A2(new_n213), .A3(new_n227), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n222), .B1(new_n328), .B2(KEYINPUT1), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n246), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  AOI21_X1  g144(.A(KEYINPUT10), .B1(new_n330), .B2(new_n324), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n325), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT3), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n318), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n317), .A2(KEYINPUT3), .A3(G104), .ZN(new_n335));
  AOI22_X1  g149(.A1(new_n334), .A2(new_n335), .B1(new_n312), .B2(G107), .ZN(new_n336));
  NAND2_X1  g150(.A1(KEYINPUT81), .A2(G101), .ZN(new_n337));
  OAI211_X1 g151(.A(new_n323), .B(KEYINPUT4), .C1(new_n336), .C2(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n313), .B1(new_n321), .B2(new_n322), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT4), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n339), .A2(KEYINPUT81), .A3(new_n340), .A4(G101), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n338), .A2(new_n219), .A3(new_n341), .A4(new_n230), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(KEYINPUT82), .ZN(new_n343));
  AND2_X1   g157(.A1(new_n230), .A2(new_n219), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT82), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n344), .A2(new_n345), .A3(new_n341), .A4(new_n338), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n209), .A2(new_n231), .ZN(new_n348));
  AND3_X1   g162(.A1(new_n332), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n348), .B1(new_n332), .B2(new_n347), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n311), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT86), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n348), .ZN(new_n354));
  AND2_X1   g168(.A1(new_n346), .A2(new_n343), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n249), .A2(new_n324), .A3(KEYINPUT10), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n330), .A2(new_n324), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n356), .B1(new_n358), .B2(KEYINPUT10), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n354), .B1(new_n355), .B2(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n332), .A2(new_n347), .A3(new_n348), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n362), .A2(KEYINPUT86), .A3(new_n311), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n353), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT85), .ZN(new_n365));
  OAI21_X1  g179(.A(KEYINPUT84), .B1(new_n249), .B2(new_n324), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n320), .A2(new_n323), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n245), .B1(new_n326), .B2(G143), .ZN(new_n368));
  OAI22_X1  g182(.A1(new_n368), .A2(new_n222), .B1(new_n228), .B2(new_n229), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT84), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n367), .A2(new_n369), .A3(new_n370), .A4(new_n246), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n366), .A2(new_n357), .A3(new_n371), .ZN(new_n372));
  AND3_X1   g186(.A1(new_n372), .A2(KEYINPUT12), .A3(new_n354), .ZN(new_n373));
  AOI21_X1  g187(.A(KEYINPUT12), .B1(new_n372), .B2(new_n354), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n365), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n372), .A2(new_n354), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT12), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n372), .A2(KEYINPUT12), .A3(new_n354), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n378), .A2(KEYINPUT85), .A3(new_n379), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n349), .A2(new_n311), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n375), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n364), .A2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(G469), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n383), .A2(new_n384), .A3(new_n276), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n361), .B1(new_n373), .B2(new_n374), .ZN(new_n386));
  AOI22_X1  g200(.A1(new_n386), .A2(new_n311), .B1(new_n381), .B2(new_n360), .ZN(new_n387));
  OAI21_X1  g201(.A(G469), .B1(new_n387), .B2(G902), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n306), .B1(new_n385), .B2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(G214), .B1(G237), .B2(G902), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n344), .A2(G125), .ZN(new_n393));
  INV_X1    g207(.A(G125), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n249), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(G224), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n397), .A2(G953), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n396), .B(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n243), .A2(new_n341), .A3(new_n338), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT5), .ZN(new_n402));
  INV_X1    g216(.A(G119), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n402), .A2(new_n403), .A3(G116), .ZN(new_n404));
  OAI211_X1 g218(.A(G113), .B(new_n404), .C1(new_n238), .C2(new_n402), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n405), .A2(new_n242), .A3(new_n324), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n401), .A2(new_n406), .ZN(new_n407));
  XOR2_X1   g221(.A(G110), .B(G122), .Z(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n408), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n401), .A2(new_n410), .A3(new_n406), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n409), .A2(KEYINPUT6), .A3(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT6), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n407), .A2(new_n413), .A3(new_n408), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n400), .A2(new_n412), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n405), .A2(new_n242), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n367), .A2(KEYINPUT87), .ZN(new_n417));
  OR2_X1    g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n416), .A2(new_n417), .ZN(new_n419));
  XOR2_X1   g233(.A(new_n408), .B(KEYINPUT8), .Z(new_n420));
  NAND3_X1  g234(.A1(new_n418), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n399), .A2(KEYINPUT7), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n393), .A2(new_n422), .A3(new_n395), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n396), .A2(KEYINPUT7), .A3(new_n399), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n421), .A2(new_n423), .A3(new_n424), .A4(new_n411), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n415), .A2(new_n276), .A3(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(G210), .B1(G237), .B2(G902), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n415), .A2(new_n425), .A3(new_n276), .A4(new_n427), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n392), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  AND2_X1   g246(.A1(new_n188), .A2(G952), .ZN(new_n433));
  NAND2_X1  g247(.A1(G234), .A2(G237), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  AND3_X1   g250(.A1(new_n434), .A2(G902), .A3(G953), .ZN(new_n437));
  XNOR2_X1  g251(.A(KEYINPUT21), .B(G898), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n436), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n432), .A2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n210), .A2(G128), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  XNOR2_X1  g257(.A(KEYINPUT66), .B(G143), .ZN(new_n444));
  OAI211_X1 g258(.A(KEYINPUT13), .B(new_n443), .C1(new_n444), .C2(new_n222), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n222), .B1(new_n211), .B2(new_n213), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  OAI211_X1 g261(.A(new_n445), .B(G134), .C1(KEYINPUT13), .C2(new_n447), .ZN(new_n448));
  AND2_X1   g262(.A1(KEYINPUT71), .A2(G116), .ZN(new_n449));
  NOR2_X1   g263(.A1(KEYINPUT71), .A2(G116), .ZN(new_n450));
  OAI21_X1  g264(.A(G122), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  OR2_X1    g265(.A1(new_n235), .A2(G122), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(G107), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n451), .A2(new_n317), .A3(new_n452), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  OAI211_X1 g270(.A(new_n195), .B(new_n443), .C1(new_n444), .C2(new_n222), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n448), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n233), .A2(KEYINPUT14), .A3(G122), .ZN(new_n459));
  OAI211_X1 g273(.A(G107), .B(new_n459), .C1(new_n453), .C2(KEYINPUT14), .ZN(new_n460));
  OAI21_X1  g274(.A(G134), .B1(new_n446), .B2(new_n442), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(new_n457), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n460), .A2(new_n462), .A3(new_n455), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n458), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n302), .A2(G217), .A3(new_n188), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n465), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n458), .A2(new_n467), .A3(new_n463), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n466), .A2(KEYINPUT90), .A3(new_n468), .ZN(new_n469));
  OR3_X1    g283(.A1(new_n464), .A2(KEYINPUT90), .A3(new_n465), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n469), .A2(new_n470), .A3(new_n276), .ZN(new_n471));
  INV_X1    g285(.A(G478), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n472), .A2(KEYINPUT15), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n473), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n469), .A2(new_n470), .A3(new_n276), .A4(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(G475), .ZN(new_n479));
  XNOR2_X1  g293(.A(G113), .B(G122), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n480), .B(new_n312), .ZN(new_n481));
  INV_X1    g295(.A(G140), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(G125), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n394), .A2(G140), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n483), .A2(new_n484), .A3(KEYINPUT76), .A4(KEYINPUT16), .ZN(new_n485));
  AND3_X1   g299(.A1(new_n483), .A2(new_n484), .A3(KEYINPUT16), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT76), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n394), .A2(G140), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT16), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  OAI211_X1 g304(.A(G146), .B(new_n485), .C1(new_n486), .C2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(KEYINPUT77), .ZN(new_n492));
  OAI21_X1  g306(.A(KEYINPUT76), .B1(new_n483), .B2(KEYINPUT16), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n483), .A2(new_n484), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n493), .B1(new_n494), .B2(new_n489), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT77), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n495), .A2(new_n496), .A3(G146), .A4(new_n485), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n492), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n494), .A2(KEYINPUT19), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT89), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n494), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n483), .A2(new_n484), .A3(KEYINPUT89), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n499), .B1(new_n503), .B2(KEYINPUT19), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(new_n326), .ZN(new_n505));
  INV_X1    g319(.A(G214), .ZN(new_n506));
  NOR3_X1   g320(.A1(new_n506), .A2(G237), .A3(G953), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n444), .A2(new_n507), .ZN(new_n508));
  NOR4_X1   g322(.A1(new_n210), .A2(new_n506), .A3(G237), .A4(G953), .ZN(new_n509));
  OAI21_X1  g323(.A(G131), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n507), .A2(G143), .ZN(new_n511));
  OAI211_X1 g325(.A(new_n511), .B(new_n207), .C1(new_n444), .C2(new_n507), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n498), .A2(new_n505), .A3(new_n513), .ZN(new_n514));
  AND2_X1   g328(.A1(KEYINPUT88), .A2(KEYINPUT18), .ZN(new_n515));
  OAI211_X1 g329(.A(G131), .B(new_n515), .C1(new_n508), .C2(new_n509), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(G131), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n511), .B(new_n517), .C1(new_n444), .C2(new_n507), .ZN(new_n518));
  INV_X1    g332(.A(new_n494), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(new_n326), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n227), .B1(new_n501), .B2(new_n502), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n516), .B(new_n518), .C1(new_n521), .C2(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n481), .B1(new_n514), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT17), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n510), .A2(new_n525), .A3(new_n512), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n495), .A2(new_n485), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(new_n227), .ZN(new_n528));
  OAI211_X1 g342(.A(KEYINPUT17), .B(G131), .C1(new_n508), .C2(new_n509), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n526), .A2(new_n528), .A3(new_n491), .A4(new_n529), .ZN(new_n530));
  AND3_X1   g344(.A1(new_n530), .A2(new_n481), .A3(new_n523), .ZN(new_n531));
  OAI211_X1 g345(.A(new_n479), .B(new_n276), .C1(new_n524), .C2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(KEYINPUT20), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n530), .A2(new_n481), .A3(new_n523), .ZN(new_n534));
  INV_X1    g348(.A(new_n523), .ZN(new_n535));
  AOI22_X1  g349(.A1(new_n492), .A2(new_n497), .B1(new_n504), .B2(new_n326), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n535), .B1(new_n536), .B2(new_n513), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n534), .B1(new_n537), .B2(new_n481), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT20), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n538), .A2(new_n539), .A3(new_n479), .A4(new_n276), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n481), .B1(new_n530), .B2(new_n523), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n276), .B1(new_n531), .B2(new_n541), .ZN(new_n542));
  AOI22_X1  g356(.A1(new_n533), .A2(new_n540), .B1(new_n542), .B2(G475), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n478), .A2(new_n543), .ZN(new_n544));
  NOR3_X1   g358(.A1(new_n390), .A2(new_n441), .A3(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT78), .ZN(new_n546));
  OAI21_X1  g360(.A(KEYINPUT75), .B1(new_n403), .B2(G128), .ZN(new_n547));
  OR2_X1    g361(.A1(new_n547), .A2(KEYINPUT23), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(KEYINPUT23), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n548), .B(new_n549), .C1(G119), .C2(new_n222), .ZN(new_n550));
  XNOR2_X1  g364(.A(G119), .B(G128), .ZN(new_n551));
  XOR2_X1   g365(.A(KEYINPUT24), .B(G110), .Z(new_n552));
  OAI22_X1  g366(.A1(new_n550), .A2(G110), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n498), .A2(new_n553), .A3(new_n520), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n528), .A2(new_n491), .ZN(new_n555));
  AOI22_X1  g369(.A1(new_n550), .A2(G110), .B1(new_n551), .B2(new_n552), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  XNOR2_X1  g372(.A(KEYINPUT22), .B(G137), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n559), .B(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n558), .B(new_n562), .ZN(new_n563));
  OR4_X1    g377(.A1(new_n546), .A2(new_n563), .A3(KEYINPUT25), .A4(G902), .ZN(new_n564));
  INV_X1    g378(.A(G217), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n565), .B1(G234), .B2(new_n276), .ZN(new_n566));
  OAI22_X1  g380(.A1(new_n563), .A2(G902), .B1(new_n546), .B2(KEYINPUT25), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n564), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n563), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n566), .A2(G902), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n300), .A2(new_n545), .A3(new_n573), .ZN(new_n574));
  XOR2_X1   g388(.A(KEYINPUT91), .B(G101), .Z(new_n575));
  XNOR2_X1  g389(.A(new_n574), .B(new_n575), .ZN(G3));
  INV_X1    g390(.A(G472), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n577), .B1(new_n288), .B2(new_n276), .ZN(new_n578));
  OR2_X1    g392(.A1(new_n578), .A2(KEYINPUT92), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(KEYINPUT92), .ZN(new_n580));
  AND4_X1   g394(.A1(new_n290), .A2(new_n579), .A3(new_n389), .A4(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n468), .ZN(new_n582));
  OR2_X1    g396(.A1(new_n582), .A2(KEYINPUT93), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(KEYINPUT93), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n583), .A2(KEYINPUT33), .A3(new_n466), .A4(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT33), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n469), .A2(new_n470), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  OAI21_X1  g402(.A(G478), .B1(new_n588), .B2(G902), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT94), .ZN(new_n590));
  OR2_X1    g404(.A1(new_n471), .A2(G478), .ZN(new_n591));
  AND3_X1   g405(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n590), .B1(new_n589), .B2(new_n591), .ZN(new_n593));
  OR2_X1    g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n533), .A2(new_n540), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n542), .A2(G475), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n598), .A2(new_n441), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n581), .A2(new_n573), .A3(new_n599), .ZN(new_n600));
  XOR2_X1   g414(.A(KEYINPUT34), .B(G104), .Z(new_n601));
  XNOR2_X1  g415(.A(new_n600), .B(new_n601), .ZN(G6));
  NOR2_X1   g416(.A1(new_n597), .A2(new_n478), .ZN(new_n603));
  AND2_X1   g417(.A1(new_n440), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n581), .A2(new_n573), .A3(new_n604), .ZN(new_n605));
  XOR2_X1   g419(.A(KEYINPUT35), .B(G107), .Z(new_n606));
  XNOR2_X1  g420(.A(new_n605), .B(new_n606), .ZN(G9));
  AND3_X1   g421(.A1(new_n579), .A2(new_n290), .A3(new_n580), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n562), .A2(KEYINPUT36), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n558), .B(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(new_n570), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n568), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n545), .A2(new_n608), .A3(new_n612), .ZN(new_n613));
  XOR2_X1   g427(.A(KEYINPUT37), .B(G110), .Z(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(G12));
  XOR2_X1   g429(.A(new_n435), .B(KEYINPUT95), .Z(new_n616));
  INV_X1    g430(.A(G900), .ZN(new_n617));
  AND2_X1   g431(.A1(new_n437), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n477), .A2(new_n595), .A3(new_n596), .A4(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(KEYINPUT96), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT96), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n543), .A2(new_n623), .A3(new_n477), .A4(new_n620), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n622), .A2(new_n431), .A3(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT97), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n622), .A2(new_n431), .A3(KEYINPUT97), .A4(new_n624), .ZN(new_n628));
  AND3_X1   g442(.A1(new_n627), .A2(new_n389), .A3(new_n628), .ZN(new_n629));
  OAI211_X1 g443(.A(new_n629), .B(new_n612), .C1(new_n299), .C2(new_n294), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(G128), .ZN(G30));
  XNOR2_X1  g445(.A(new_n619), .B(KEYINPUT39), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n390), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(KEYINPUT40), .ZN(new_n634));
  AND2_X1   g448(.A1(new_n296), .A2(new_n298), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT100), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n273), .B1(new_n272), .B2(new_n258), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n276), .B1(new_n265), .B2(new_n193), .ZN(new_n638));
  OAI21_X1  g452(.A(G472), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n635), .A2(new_n636), .A3(new_n292), .A4(new_n639), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n296), .A2(new_n292), .A3(new_n298), .A4(new_n639), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(KEYINPUT100), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n429), .A2(new_n430), .ZN(new_n644));
  XNOR2_X1  g458(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(KEYINPUT99), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n644), .B(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n597), .A2(new_n477), .ZN(new_n648));
  NOR3_X1   g462(.A1(new_n612), .A2(new_n648), .A3(new_n392), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(KEYINPUT101), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n634), .A2(new_n643), .A3(new_n647), .A4(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(new_n651), .B(KEYINPUT102), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(new_n444), .ZN(G45));
  OAI21_X1  g467(.A(new_n612), .B1(new_n294), .B2(new_n299), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  OAI211_X1 g469(.A(new_n597), .B(new_n620), .C1(new_n592), .C2(new_n593), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n655), .A2(new_n431), .A3(new_n389), .A4(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(G146), .ZN(G48));
  NOR2_X1   g473(.A1(new_n294), .A2(new_n299), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n660), .A2(new_n572), .ZN(new_n661));
  AND2_X1   g475(.A1(new_n375), .A2(new_n380), .ZN(new_n662));
  AOI22_X1  g476(.A1(new_n662), .A2(new_n381), .B1(new_n353), .B2(new_n363), .ZN(new_n663));
  OAI21_X1  g477(.A(G469), .B1(new_n663), .B2(G902), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT103), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n664), .A2(new_n665), .A3(new_n385), .ZN(new_n666));
  OAI211_X1 g480(.A(KEYINPUT103), .B(G469), .C1(new_n663), .C2(G902), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n304), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n661), .A2(new_n599), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(KEYINPUT41), .B(G113), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G15));
  NAND3_X1  g487(.A1(new_n661), .A2(new_n604), .A3(new_n670), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G116), .ZN(G18));
  NOR3_X1   g489(.A1(new_n654), .A2(new_n432), .A3(new_n544), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n669), .A2(new_n439), .ZN(new_n677));
  AOI21_X1  g491(.A(KEYINPUT104), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n676), .A2(KEYINPUT104), .A3(new_n677), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G119), .ZN(G21));
  NAND2_X1  g496(.A1(new_n288), .A2(new_n276), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n277), .A2(new_n273), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n284), .A2(new_n684), .A3(new_n287), .ZN(new_n685));
  AOI22_X1  g499(.A1(new_n683), .A2(G472), .B1(new_n289), .B2(new_n685), .ZN(new_n686));
  AND2_X1   g500(.A1(new_n686), .A2(new_n573), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n648), .A2(KEYINPUT105), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT105), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n597), .A2(new_n689), .A3(new_n477), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n688), .A2(new_n431), .A3(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n677), .A2(new_n687), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G122), .ZN(G24));
  NAND2_X1  g508(.A1(new_n686), .A2(new_n612), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT106), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n686), .A2(KEYINPUT106), .A3(new_n612), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(new_n304), .ZN(new_n700));
  AOI211_X1 g514(.A(new_n432), .B(new_n700), .C1(new_n666), .C2(new_n667), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n699), .A2(new_n701), .A3(new_n657), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G125), .ZN(G27));
  NOR2_X1   g517(.A1(new_n644), .A2(new_n392), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n300), .A2(new_n573), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n385), .A2(new_n388), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(new_n304), .ZN(new_n707));
  NOR4_X1   g521(.A1(new_n705), .A2(KEYINPUT42), .A3(new_n656), .A4(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT42), .ZN(new_n709));
  INV_X1    g523(.A(new_n598), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n700), .B1(new_n385), .B2(new_n388), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(new_n295), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n573), .B1(new_n294), .B2(new_n713), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(new_n704), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n716), .A2(new_n619), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n709), .B1(new_n715), .B2(new_n717), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n708), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G131), .ZN(G33));
  NAND2_X1  g534(.A1(new_n622), .A2(new_n624), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(KEYINPUT107), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n705), .A2(new_n707), .A3(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(new_n195), .ZN(G36));
  INV_X1    g538(.A(KEYINPUT108), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(KEYINPUT43), .ZN(new_n726));
  XOR2_X1   g540(.A(KEYINPUT108), .B(KEYINPUT43), .Z(new_n727));
  AND2_X1   g541(.A1(new_n594), .A2(new_n543), .ZN(new_n728));
  MUX2_X1   g542(.A(new_n726), .B(new_n727), .S(new_n728), .Z(new_n729));
  INV_X1    g543(.A(new_n608), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n729), .A2(new_n730), .A3(new_n612), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(KEYINPUT44), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n704), .ZN(new_n733));
  OR2_X1    g547(.A1(new_n733), .A2(KEYINPUT109), .ZN(new_n734));
  XOR2_X1   g548(.A(new_n387), .B(KEYINPUT45), .Z(new_n735));
  OAI21_X1  g549(.A(G469), .B1(new_n735), .B2(G902), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(KEYINPUT46), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n385), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n736), .A2(KEYINPUT46), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n304), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  OR2_X1    g554(.A1(new_n740), .A2(new_n632), .ZN(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n733), .A2(KEYINPUT109), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n734), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G137), .ZN(G39));
  XOR2_X1   g559(.A(KEYINPUT110), .B(KEYINPUT47), .Z(new_n746));
  NOR2_X1   g560(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n747));
  MUX2_X1   g561(.A(new_n746), .B(new_n747), .S(new_n740), .Z(new_n748));
  NOR3_X1   g562(.A1(new_n716), .A2(new_n573), .A3(new_n619), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n748), .A2(new_n660), .A3(new_n710), .A4(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G140), .ZN(G42));
  XOR2_X1   g565(.A(new_n668), .B(KEYINPUT49), .Z(new_n752));
  NOR2_X1   g566(.A1(new_n752), .A2(new_n572), .ZN(new_n753));
  INV_X1    g567(.A(new_n643), .ZN(new_n754));
  NOR3_X1   g568(.A1(new_n647), .A2(new_n392), .A3(new_n306), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n753), .A2(new_n754), .A3(new_n728), .A4(new_n755), .ZN(new_n756));
  AND2_X1   g570(.A1(new_n729), .A2(new_n616), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n669), .A2(new_n716), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n759), .A2(new_n714), .ZN(new_n760));
  XOR2_X1   g574(.A(new_n760), .B(KEYINPUT48), .Z(new_n761));
  NAND4_X1  g575(.A1(new_n754), .A2(new_n573), .A3(new_n436), .A4(new_n758), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(KEYINPUT120), .ZN(new_n763));
  OAI211_X1 g577(.A(new_n761), .B(new_n433), .C1(new_n598), .C2(new_n763), .ZN(new_n764));
  AND2_X1   g578(.A1(new_n757), .A2(new_n687), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n647), .A2(new_n391), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n765), .A2(new_n670), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(KEYINPUT119), .A2(KEYINPUT50), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g583(.A1(KEYINPUT119), .A2(KEYINPUT50), .ZN(new_n770));
  XOR2_X1   g584(.A(new_n769), .B(new_n770), .Z(new_n771));
  NOR3_X1   g585(.A1(new_n763), .A2(new_n597), .A3(new_n594), .ZN(new_n772));
  INV_X1    g586(.A(new_n759), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n772), .B1(new_n699), .B2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(new_n668), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n775), .A2(new_n305), .ZN(new_n776));
  OAI211_X1 g590(.A(new_n765), .B(new_n704), .C1(new_n748), .C2(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n771), .A2(new_n774), .A3(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT51), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n764), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n765), .A2(new_n701), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n774), .A2(KEYINPUT121), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n774), .B1(KEYINPUT121), .B2(new_n779), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n783), .A2(new_n771), .A3(new_n777), .ZN(new_n784));
  OAI211_X1 g598(.A(new_n780), .B(new_n781), .C1(new_n782), .C2(new_n784), .ZN(new_n785));
  AND3_X1   g599(.A1(new_n686), .A2(KEYINPUT106), .A3(new_n612), .ZN(new_n786));
  AOI21_X1  g600(.A(KEYINPUT106), .B1(new_n686), .B2(new_n612), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n668), .A2(new_n657), .A3(new_n431), .A4(new_n304), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n627), .A2(new_n389), .A3(new_n628), .ZN(new_n790));
  OAI22_X1  g604(.A1(new_n788), .A2(new_n789), .B1(new_n654), .B2(new_n790), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n791), .A2(KEYINPUT112), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT112), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n793), .B1(new_n702), .B2(new_n630), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT52), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n612), .A2(new_n619), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n692), .A2(new_n711), .A3(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n641), .A2(KEYINPUT100), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n641), .A2(KEYINPUT100), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n799), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(KEYINPUT113), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT113), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n643), .A2(new_n804), .A3(new_n799), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n796), .B1(new_n803), .B2(new_n805), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n795), .A2(KEYINPUT114), .A3(new_n658), .A4(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT114), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n791), .A2(KEYINPUT112), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n702), .A2(new_n630), .A3(new_n793), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n809), .A2(new_n810), .A3(new_n658), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n804), .B1(new_n643), .B2(new_n799), .ZN(new_n812));
  AOI211_X1 g626(.A(KEYINPUT113), .B(new_n798), .C1(new_n640), .C2(new_n642), .ZN(new_n813));
  OAI21_X1  g627(.A(KEYINPUT52), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n808), .B1(new_n811), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n812), .A2(new_n813), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n658), .A2(new_n630), .A3(new_n702), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n796), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n807), .A2(new_n815), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(KEYINPUT115), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT115), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n807), .A2(new_n815), .A3(new_n821), .A4(new_n818), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  OAI211_X1 g637(.A(new_n581), .B(new_n573), .C1(new_n599), .C2(new_n604), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n824), .A2(new_n574), .A3(new_n613), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(KEYINPUT111), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT111), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n824), .A2(new_n574), .A3(new_n613), .A4(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n826), .A2(new_n671), .A3(new_n693), .A4(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n708), .A2(new_n723), .A3(new_n718), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n655), .A2(new_n478), .A3(new_n543), .A4(new_n389), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n832), .B1(new_n788), .B2(new_n712), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(new_n717), .ZN(new_n834));
  INV_X1    g648(.A(new_n674), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n835), .B1(new_n679), .B2(new_n680), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n830), .A2(new_n831), .A3(new_n834), .A4(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n823), .A2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT53), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n839), .A2(KEYINPUT116), .A3(new_n840), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n816), .A2(new_n817), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(KEYINPUT52), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(new_n818), .ZN(new_n844));
  XNOR2_X1  g658(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n838), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT116), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n837), .B1(new_n820), .B2(new_n822), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n847), .B1(new_n848), .B2(KEYINPUT53), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n841), .A2(new_n846), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(KEYINPUT54), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n848), .A2(KEYINPUT53), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n838), .A2(new_n844), .ZN(new_n853));
  INV_X1    g667(.A(new_n845), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  OR2_X1    g670(.A1(new_n856), .A2(KEYINPUT54), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n851), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(KEYINPUT118), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT118), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n851), .A2(new_n860), .A3(new_n857), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n785), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(G952), .A2(G953), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n756), .B1(new_n862), .B2(new_n863), .ZN(G75));
  AOI21_X1  g678(.A(new_n276), .B1(new_n852), .B2(new_n855), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(G210), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT56), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n412), .A2(new_n414), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n868), .B(new_n400), .ZN(new_n869));
  XOR2_X1   g683(.A(new_n869), .B(KEYINPUT55), .Z(new_n870));
  INV_X1    g684(.A(KEYINPUT122), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n870), .B1(new_n871), .B2(new_n867), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n866), .A2(new_n867), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n872), .B1(new_n866), .B2(new_n867), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n188), .A2(G952), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(G51));
  XNOR2_X1  g690(.A(new_n856), .B(KEYINPUT54), .ZN(new_n877));
  NAND2_X1  g691(.A1(G469), .A2(G902), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n878), .B(KEYINPUT123), .ZN(new_n879));
  INV_X1    g693(.A(new_n879), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n877), .B1(KEYINPUT57), .B2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT57), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n383), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n865), .A2(G469), .A3(new_n735), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n875), .B1(new_n884), .B2(new_n885), .ZN(G54));
  NAND3_X1  g700(.A1(new_n865), .A2(KEYINPUT58), .A3(G475), .ZN(new_n887));
  INV_X1    g701(.A(new_n538), .ZN(new_n888));
  AND2_X1   g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n887), .A2(new_n888), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n889), .A2(new_n890), .A3(new_n875), .ZN(G60));
  NAND2_X1  g705(.A1(G478), .A2(G902), .ZN(new_n892));
  XOR2_X1   g706(.A(new_n892), .B(KEYINPUT59), .Z(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n877), .A2(new_n587), .A3(new_n585), .A4(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(new_n875), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n859), .A2(new_n861), .A3(new_n894), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n897), .B1(new_n898), .B2(new_n588), .ZN(G63));
  NAND2_X1  g713(.A1(G217), .A2(G902), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(KEYINPUT60), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n901), .B1(new_n852), .B2(new_n855), .ZN(new_n902));
  OR2_X1    g716(.A1(new_n902), .A2(new_n569), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n610), .B(KEYINPUT124), .Z(new_n904));
  NAND2_X1  g718(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n903), .A2(new_n896), .A3(new_n905), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n906), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g721(.A(G953), .B1(new_n438), .B2(new_n397), .ZN(new_n908));
  INV_X1    g722(.A(new_n836), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n909), .A2(new_n829), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n908), .B1(new_n910), .B2(G953), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n868), .B1(G898), .B2(new_n188), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n911), .B(new_n912), .ZN(G69));
  NOR2_X1   g727(.A1(new_n268), .A2(new_n271), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(new_n504), .ZN(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(new_n705), .ZN(new_n917));
  OAI211_X1 g731(.A(new_n917), .B(new_n633), .C1(new_n710), .C2(new_n603), .ZN(new_n918));
  AND3_X1   g732(.A1(new_n744), .A2(new_n750), .A3(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(new_n811), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n652), .A2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n922), .A2(KEYINPUT62), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(KEYINPUT62), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n919), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n916), .B1(new_n926), .B2(new_n188), .ZN(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  OAI21_X1  g742(.A(G953), .B1(new_n308), .B2(new_n617), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(KEYINPUT126), .ZN(new_n930));
  OR2_X1    g744(.A1(new_n929), .A2(KEYINPUT126), .ZN(new_n931));
  NAND2_X1  g745(.A1(G900), .A2(G953), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n741), .A2(new_n691), .A3(new_n714), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n933), .B(KEYINPUT125), .Z(new_n934));
  AND2_X1   g748(.A1(new_n934), .A2(new_n831), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n744), .A2(new_n935), .A3(new_n750), .A4(new_n920), .ZN(new_n936));
  OAI211_X1 g750(.A(new_n916), .B(new_n932), .C1(new_n936), .C2(G953), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n928), .A2(new_n930), .A3(new_n931), .A4(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(new_n937), .ZN(new_n939));
  OAI211_X1 g753(.A(KEYINPUT126), .B(new_n929), .C1(new_n927), .C2(new_n939), .ZN(new_n940));
  AND2_X1   g754(.A1(new_n938), .A2(new_n940), .ZN(G72));
  INV_X1    g755(.A(new_n637), .ZN(new_n942));
  OAI211_X1 g756(.A(new_n919), .B(new_n910), .C1(new_n923), .C2(new_n925), .ZN(new_n943));
  NAND2_X1  g757(.A1(G472), .A2(G902), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(KEYINPUT63), .Z(new_n945));
  AOI21_X1  g759(.A(new_n942), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  AND4_X1   g760(.A1(new_n274), .A2(new_n850), .A3(new_n942), .A4(new_n945), .ZN(new_n947));
  INV_X1    g761(.A(new_n910), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n945), .B1(new_n936), .B2(new_n948), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n274), .B(KEYINPUT127), .Z(new_n950));
  AND2_X1   g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NOR4_X1   g765(.A1(new_n946), .A2(new_n947), .A3(new_n951), .A4(new_n875), .ZN(G57));
endmodule


