//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 0 0 1 0 1 1 0 0 0 1 0 0 1 1 0 0 1 0 1 0 0 1 0 1 1 1 1 0 0 0 1 1 0 1 0 0 1 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:30 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n730, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n950, new_n951, new_n952, new_n953, new_n954, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n970, new_n971,
    new_n972, new_n973, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007;
  INV_X1    g000(.A(KEYINPUT28), .ZN(new_n187));
  INV_X1    g001(.A(G131), .ZN(new_n188));
  INV_X1    g002(.A(G134), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G137), .ZN(new_n190));
  INV_X1    g004(.A(G137), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G134), .ZN(new_n192));
  AOI21_X1  g006(.A(new_n188), .B1(new_n190), .B2(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n193), .B(KEYINPUT64), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT67), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT11), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n196), .B1(new_n189), .B2(G137), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n191), .A2(KEYINPUT11), .A3(G134), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n197), .A2(new_n198), .A3(new_n188), .A4(new_n190), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G143), .ZN(new_n201));
  INV_X1    g015(.A(G143), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G146), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT1), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n201), .A2(new_n203), .A3(new_n204), .A4(G128), .ZN(new_n205));
  INV_X1    g019(.A(G128), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n206), .B1(new_n201), .B2(KEYINPUT1), .ZN(new_n207));
  XNOR2_X1  g021(.A(G143), .B(G146), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n205), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n194), .A2(new_n195), .A3(new_n199), .A4(new_n209), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n193), .A2(KEYINPUT64), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT64), .ZN(new_n212));
  AOI211_X1 g026(.A(new_n212), .B(new_n188), .C1(new_n190), .C2(new_n192), .ZN(new_n213));
  OAI211_X1 g027(.A(new_n209), .B(new_n199), .C1(new_n211), .C2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(KEYINPUT67), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n197), .A2(new_n190), .A3(new_n198), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G131), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(new_n199), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n201), .A2(new_n203), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT0), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n220), .A2(new_n206), .ZN(new_n221));
  NOR2_X1   g035(.A1(KEYINPUT0), .A2(G128), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n219), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n208), .B1(new_n220), .B2(new_n206), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n218), .A2(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n210), .A2(new_n215), .A3(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT2), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n228), .A2(G113), .ZN(new_n229));
  INV_X1    g043(.A(G113), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n230), .A2(KEYINPUT2), .ZN(new_n231));
  NOR2_X1   g045(.A1(G116), .A2(G119), .ZN(new_n232));
  AND2_X1   g046(.A1(G116), .A2(G119), .ZN(new_n233));
  OAI22_X1  g047(.A1(new_n229), .A2(new_n231), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n232), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n230), .A2(KEYINPUT2), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n228), .A2(G113), .ZN(new_n237));
  NAND2_X1  g051(.A1(G116), .A2(G119), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n235), .A2(new_n236), .A3(new_n237), .A4(new_n238), .ZN(new_n239));
  AND3_X1   g053(.A1(new_n234), .A2(new_n239), .A3(KEYINPUT66), .ZN(new_n240));
  AOI21_X1  g054(.A(KEYINPUT66), .B1(new_n234), .B2(new_n239), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n227), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n242), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n244), .A2(new_n210), .A3(new_n215), .A4(new_n226), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n187), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n226), .A2(new_n214), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n187), .B1(new_n247), .B2(new_n242), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n246), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g064(.A(KEYINPUT68), .B(G953), .ZN(new_n251));
  INV_X1    g065(.A(G237), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n251), .A2(G210), .A3(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT70), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XOR2_X1   g069(.A(KEYINPUT26), .B(G101), .Z(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  XNOR2_X1  g072(.A(new_n253), .B(KEYINPUT70), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(new_n256), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  XNOR2_X1  g075(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n258), .A2(new_n260), .A3(new_n262), .ZN(new_n265));
  AND2_X1   g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT29), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(G902), .B1(new_n250), .B2(new_n268), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n210), .A2(new_n215), .A3(KEYINPUT30), .A4(new_n226), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT30), .ZN(new_n271));
  AOI21_X1  g085(.A(KEYINPUT65), .B1(new_n247), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT65), .ZN(new_n273));
  AOI211_X1 g087(.A(new_n273), .B(KEYINPUT30), .C1(new_n226), .C2(new_n214), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n242), .B(new_n270), .C1(new_n272), .C2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(new_n245), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(new_n266), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(new_n267), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n247), .A2(new_n242), .ZN(new_n279));
  OAI211_X1 g093(.A(new_n279), .B(new_n248), .C1(new_n245), .C2(new_n187), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n266), .A2(new_n280), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n269), .B1(new_n278), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(G472), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n264), .A2(new_n265), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n275), .A2(new_n245), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(KEYINPUT31), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT31), .ZN(new_n287));
  NAND4_X1  g101(.A1(new_n275), .A2(new_n284), .A3(new_n287), .A4(new_n245), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n266), .A2(new_n280), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n286), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT32), .ZN(new_n291));
  NOR2_X1   g105(.A1(G472), .A2(G902), .ZN(new_n292));
  AND3_X1   g106(.A1(new_n290), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n291), .B1(new_n290), .B2(new_n292), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n283), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  XNOR2_X1  g109(.A(KEYINPUT74), .B(KEYINPUT22), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n251), .A2(G221), .A3(G234), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(G137), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n251), .A2(new_n191), .A3(G221), .A4(G234), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n296), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n298), .A2(new_n296), .A3(new_n299), .ZN(new_n302));
  AOI21_X1  g116(.A(KEYINPUT75), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(new_n302), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT75), .ZN(new_n305));
  NOR3_X1   g119(.A1(new_n304), .A2(new_n305), .A3(new_n300), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n303), .A2(new_n306), .ZN(new_n307));
  XNOR2_X1  g121(.A(G125), .B(G140), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(KEYINPUT16), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT16), .ZN(new_n310));
  INV_X1    g124(.A(G140), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n310), .A2(new_n311), .A3(G125), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(KEYINPUT72), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT72), .ZN(new_n314));
  NAND4_X1  g128(.A1(new_n314), .A2(new_n310), .A3(new_n311), .A4(G125), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n309), .A2(new_n313), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(new_n200), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n309), .A2(G146), .A3(new_n313), .A4(new_n315), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  XOR2_X1   g133(.A(KEYINPUT24), .B(G110), .Z(new_n320));
  XNOR2_X1  g134(.A(G119), .B(G128), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT71), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT23), .ZN(new_n324));
  INV_X1    g138(.A(G119), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n324), .B1(new_n325), .B2(G128), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n206), .A2(KEYINPUT23), .A3(G119), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n326), .B(new_n327), .C1(G119), .C2(new_n206), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n323), .B1(new_n328), .B2(G110), .ZN(new_n329));
  AND3_X1   g143(.A1(new_n328), .A2(new_n323), .A3(G110), .ZN(new_n330));
  OAI211_X1 g144(.A(new_n319), .B(new_n322), .C1(new_n329), .C2(new_n330), .ZN(new_n331));
  OAI22_X1  g145(.A1(new_n328), .A2(G110), .B1(new_n321), .B2(new_n320), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n308), .A2(new_n200), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n332), .A2(new_n318), .A3(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(KEYINPUT73), .B1(new_n331), .B2(new_n334), .ZN(new_n335));
  AND2_X1   g149(.A1(new_n317), .A2(new_n318), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n322), .B1(new_n330), .B2(new_n329), .ZN(new_n337));
  OAI211_X1 g151(.A(KEYINPUT73), .B(new_n334), .C1(new_n336), .C2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n307), .B1(new_n335), .B2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(G902), .ZN(new_n341));
  OAI211_X1 g155(.A(new_n331), .B(new_n334), .C1(new_n304), .C2(new_n300), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(KEYINPUT25), .ZN(new_n344));
  INV_X1    g158(.A(G217), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n345), .B1(G234), .B2(new_n341), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT25), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n340), .A2(new_n347), .A3(new_n341), .A4(new_n342), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n344), .A2(new_n346), .A3(new_n348), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n346), .A2(G902), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n340), .A2(new_n342), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n295), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(G104), .ZN(new_n356));
  OAI21_X1  g170(.A(KEYINPUT3), .B1(new_n356), .B2(G107), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT3), .ZN(new_n358));
  INV_X1    g172(.A(G107), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n358), .A2(new_n359), .A3(G104), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n356), .A2(G107), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n357), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n362), .A2(KEYINPUT77), .A3(G101), .ZN(new_n363));
  INV_X1    g177(.A(G101), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n357), .A2(new_n360), .A3(new_n364), .A4(new_n361), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(KEYINPUT4), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n362), .A2(KEYINPUT77), .A3(KEYINPUT4), .A4(G101), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(new_n242), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n359), .A2(G104), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n356), .A2(G107), .ZN(new_n372));
  OAI21_X1  g186(.A(G101), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  AND2_X1   g187(.A1(new_n365), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n236), .A2(new_n237), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n235), .A2(new_n238), .ZN(new_n376));
  OAI21_X1  g190(.A(KEYINPUT5), .B1(new_n233), .B2(new_n232), .ZN(new_n377));
  NOR2_X1   g191(.A1(KEYINPUT5), .A2(G119), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n230), .B1(new_n378), .B2(G116), .ZN(new_n379));
  AOI22_X1  g193(.A1(new_n375), .A2(new_n376), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n374), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(KEYINPUT84), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT84), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n374), .A2(new_n380), .A3(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n370), .A2(new_n382), .A3(new_n384), .ZN(new_n385));
  XOR2_X1   g199(.A(G110), .B(G122), .Z(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(new_n386), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n370), .A2(new_n382), .A3(new_n388), .A4(new_n384), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n387), .A2(KEYINPUT6), .A3(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT6), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n385), .A2(new_n391), .A3(new_n386), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n223), .A2(new_n224), .A3(G125), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT85), .ZN(new_n394));
  OR2_X1    g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n393), .B(new_n394), .C1(G125), .C2(new_n209), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(G953), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(G224), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n397), .B(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n390), .A2(new_n392), .A3(new_n400), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n386), .A2(KEYINPUT8), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n365), .A2(new_n373), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n402), .B1(new_n380), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n386), .A2(KEYINPUT8), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n379), .B(KEYINPUT86), .ZN(new_n406));
  AOI22_X1  g220(.A1(new_n406), .A2(new_n377), .B1(new_n375), .B2(new_n376), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n404), .B(new_n405), .C1(new_n407), .C2(new_n403), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT7), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n395), .A2(new_n396), .A3(new_n409), .ZN(new_n410));
  AND2_X1   g224(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  OR2_X1    g225(.A1(new_n397), .A2(new_n399), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n397), .A2(KEYINPUT7), .A3(new_n399), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n411), .A2(new_n389), .A3(new_n412), .A4(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n401), .A2(new_n341), .A3(new_n414), .ZN(new_n415));
  OAI21_X1  g229(.A(G210), .B1(G237), .B2(G902), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT87), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n401), .A2(new_n414), .A3(new_n341), .A4(new_n416), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n418), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(G214), .B1(G237), .B2(G902), .ZN(new_n422));
  OR2_X1    g236(.A1(new_n420), .A2(new_n419), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n421), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(G469), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n204), .B1(G143), .B2(new_n200), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT78), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n206), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n201), .A2(KEYINPUT1), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(KEYINPUT78), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n208), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n205), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n374), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  XNOR2_X1  g247(.A(KEYINPUT79), .B(KEYINPUT10), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n369), .A2(new_n225), .ZN(new_n437));
  INV_X1    g251(.A(new_n218), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n374), .A2(KEYINPUT10), .A3(new_n209), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n436), .A2(new_n437), .A3(new_n438), .A4(new_n439), .ZN(new_n440));
  XNOR2_X1  g254(.A(G110), .B(G140), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n441), .B(KEYINPUT76), .ZN(new_n442));
  AND2_X1   g256(.A1(new_n251), .A2(G227), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n442), .B(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n440), .A2(new_n444), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n403), .B(new_n205), .C1(new_n208), .C2(new_n207), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n438), .B1(new_n433), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(KEYINPUT81), .B1(new_n447), .B2(KEYINPUT12), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n374), .A2(new_n209), .ZN(new_n449));
  OAI211_X1 g263(.A(new_n427), .B(KEYINPUT1), .C1(new_n202), .C2(G146), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(G128), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n427), .B1(new_n201), .B2(KEYINPUT1), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n219), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n403), .B1(new_n453), .B2(new_n205), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n218), .B1(new_n449), .B2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT81), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT12), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n448), .A2(new_n458), .ZN(new_n459));
  OAI211_X1 g273(.A(KEYINPUT12), .B(new_n218), .C1(new_n449), .C2(new_n454), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(KEYINPUT80), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n433), .A2(new_n446), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT80), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n462), .A2(new_n463), .A3(KEYINPUT12), .A4(new_n218), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n445), .B1(new_n459), .B2(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n439), .B1(new_n454), .B2(new_n434), .ZN(new_n467));
  AOI22_X1  g281(.A1(new_n367), .A2(new_n368), .B1(new_n223), .B2(new_n224), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n218), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n444), .B1(new_n440), .B2(new_n469), .ZN(new_n470));
  OAI211_X1 g284(.A(new_n425), .B(new_n341), .C1(new_n466), .C2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT82), .ZN(new_n472));
  NOR3_X1   g286(.A1(new_n467), .A2(new_n218), .A3(new_n468), .ZN(new_n473));
  INV_X1    g287(.A(new_n444), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n440), .A2(KEYINPUT82), .A3(new_n444), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n475), .A2(new_n469), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n473), .B1(new_n459), .B2(new_n465), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n477), .B(G469), .C1(new_n478), .C2(new_n444), .ZN(new_n479));
  NAND2_X1  g293(.A1(G469), .A2(G902), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n471), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(G221), .ZN(new_n482));
  XOR2_X1   g296(.A(KEYINPUT9), .B(G234), .Z(new_n483));
  AOI21_X1  g297(.A(new_n482), .B1(new_n483), .B2(new_n341), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  AND3_X1   g299(.A1(new_n481), .A2(KEYINPUT83), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(KEYINPUT83), .B1(new_n481), .B2(new_n485), .ZN(new_n487));
  NOR3_X1   g301(.A1(new_n424), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(G952), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n489), .A2(G953), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n491), .B1(G234), .B2(G237), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  AOI211_X1 g307(.A(new_n341), .B(new_n251), .C1(G234), .C2(G237), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  XOR2_X1   g309(.A(KEYINPUT21), .B(G898), .Z(new_n496));
  OAI21_X1  g310(.A(new_n493), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  XNOR2_X1  g312(.A(G116), .B(G122), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(new_n359), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  OR2_X1    g315(.A1(new_n501), .A2(KEYINPUT93), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n202), .A2(G128), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n206), .A2(G143), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n505), .B(new_n189), .ZN(new_n506));
  INV_X1    g320(.A(G116), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n507), .A2(KEYINPUT14), .A3(G122), .ZN(new_n508));
  INV_X1    g322(.A(new_n499), .ZN(new_n509));
  OAI211_X1 g323(.A(G107), .B(new_n508), .C1(new_n509), .C2(KEYINPUT14), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n501), .A2(KEYINPUT93), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n502), .A2(new_n506), .A3(new_n510), .A4(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT91), .ZN(new_n513));
  AOI21_X1  g327(.A(KEYINPUT13), .B1(new_n202), .B2(G128), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n513), .B1(new_n514), .B2(new_n503), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n206), .A2(G143), .ZN(new_n516));
  OAI211_X1 g330(.A(KEYINPUT91), .B(new_n516), .C1(new_n504), .C2(KEYINPUT13), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n504), .A2(KEYINPUT13), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n515), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n509), .A2(G107), .ZN(new_n520));
  AOI22_X1  g334(.A1(new_n519), .A2(G134), .B1(new_n520), .B2(new_n500), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n505), .A2(new_n189), .ZN(new_n522));
  AND3_X1   g336(.A1(new_n521), .A2(KEYINPUT92), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(KEYINPUT92), .B1(new_n521), .B2(new_n522), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n512), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n483), .A2(G217), .A3(new_n398), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT94), .ZN(new_n528));
  INV_X1    g342(.A(new_n526), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n512), .B(new_n529), .C1(new_n523), .C2(new_n524), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n527), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  OR3_X1    g345(.A1(new_n525), .A2(new_n528), .A3(new_n526), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n531), .A2(new_n532), .A3(new_n341), .ZN(new_n533));
  INV_X1    g347(.A(G478), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n534), .A2(KEYINPUT15), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n535), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n531), .A2(new_n532), .A3(new_n341), .A4(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  AND2_X1   g353(.A1(KEYINPUT68), .A2(G953), .ZN(new_n540));
  NOR2_X1   g354(.A1(KEYINPUT68), .A2(G953), .ZN(new_n541));
  OAI211_X1 g355(.A(G214), .B(new_n252), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(new_n202), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n251), .A2(G143), .A3(G214), .A4(new_n252), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(G131), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT17), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n543), .A2(new_n544), .A3(new_n188), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n545), .A2(KEYINPUT17), .A3(G131), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n549), .A2(new_n336), .A3(new_n550), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n308), .B(new_n200), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT18), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n553), .A2(new_n188), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n552), .B1(new_n545), .B2(new_n554), .ZN(new_n555));
  AOI211_X1 g369(.A(new_n553), .B(new_n188), .C1(new_n543), .C2(new_n544), .ZN(new_n556));
  OR2_X1    g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  XNOR2_X1  g371(.A(G113), .B(G122), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n558), .B(new_n356), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n551), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n559), .ZN(new_n561));
  NAND2_X1  g375(.A1(KEYINPUT88), .A2(KEYINPUT19), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n308), .A2(new_n562), .ZN(new_n563));
  XOR2_X1   g377(.A(KEYINPUT88), .B(KEYINPUT19), .Z(new_n564));
  OAI21_X1  g378(.A(new_n563), .B1(new_n308), .B2(new_n564), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n318), .B1(new_n565), .B2(G146), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n566), .B1(new_n546), .B2(new_n548), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n555), .A2(new_n556), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n561), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n560), .A2(new_n569), .ZN(new_n570));
  NOR2_X1   g384(.A1(G475), .A2(G902), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT20), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n572), .A2(KEYINPUT89), .A3(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n560), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n559), .B1(new_n551), .B2(new_n557), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n341), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(G475), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT89), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n570), .A2(new_n579), .A3(new_n571), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(KEYINPUT20), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n579), .B1(new_n570), .B2(new_n571), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n574), .B(new_n578), .C1(new_n581), .C2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(KEYINPUT90), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n572), .A2(KEYINPUT89), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n585), .A2(KEYINPUT20), .A3(new_n580), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT90), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n586), .A2(new_n587), .A3(new_n574), .A4(new_n578), .ZN(new_n588));
  AOI211_X1 g402(.A(new_n498), .B(new_n539), .C1(new_n584), .C2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n355), .A2(new_n488), .A3(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(G101), .ZN(G3));
  NAND2_X1  g405(.A1(new_n533), .A2(new_n534), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT33), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n531), .A2(new_n532), .A3(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n526), .B(KEYINPUT96), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n525), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT97), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n525), .A2(KEYINPUT97), .A3(new_n595), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n598), .A2(KEYINPUT33), .A3(new_n530), .A4(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n594), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n341), .A2(G478), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n592), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n584), .A2(new_n603), .A3(new_n588), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(KEYINPUT98), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT98), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  AND2_X1   g422(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n418), .A2(new_n420), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(new_n422), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n611), .A2(new_n498), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n481), .A2(new_n485), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT83), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n481), .A2(KEYINPUT83), .A3(new_n485), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  AND2_X1   g431(.A1(new_n288), .A2(new_n289), .ZN(new_n618));
  AOI21_X1  g432(.A(G902), .B1(new_n618), .B2(new_n286), .ZN(new_n619));
  INV_X1    g433(.A(G472), .ZN(new_n620));
  OAI21_X1  g434(.A(KEYINPUT95), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  AND2_X1   g435(.A1(new_n285), .A2(KEYINPUT31), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n288), .A2(new_n289), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n292), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n290), .A2(new_n341), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT95), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n625), .A2(new_n626), .A3(G472), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n621), .A2(new_n624), .A3(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n617), .A2(new_n628), .ZN(new_n629));
  AND4_X1   g443(.A1(new_n353), .A2(new_n609), .A3(new_n612), .A4(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(KEYINPUT34), .B(G104), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G6));
  INV_X1    g446(.A(new_n539), .ZN(new_n633));
  NOR4_X1   g447(.A1(new_n611), .A2(new_n633), .A3(new_n583), .A4(new_n498), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n629), .A2(new_n353), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(G107), .ZN(new_n636));
  XNOR2_X1  g450(.A(KEYINPUT99), .B(KEYINPUT35), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G9));
  OR2_X1    g452(.A1(new_n335), .A2(new_n339), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n307), .A2(KEYINPUT36), .ZN(new_n640));
  AND2_X1   g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n350), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  AND2_X1   g457(.A1(new_n349), .A2(new_n643), .ZN(new_n644));
  OAI21_X1  g458(.A(KEYINPUT100), .B1(new_n628), .B2(new_n644), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n626), .B1(new_n625), .B2(G472), .ZN(new_n646));
  AOI211_X1 g460(.A(KEYINPUT95), .B(new_n620), .C1(new_n290), .C2(new_n341), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT100), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n349), .A2(new_n643), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n648), .A2(new_n649), .A3(new_n624), .A4(new_n650), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n645), .A2(new_n651), .A3(new_n589), .A4(new_n488), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G110), .ZN(new_n653));
  XNOR2_X1  g467(.A(KEYINPUT101), .B(KEYINPUT37), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G12));
  NAND2_X1  g469(.A1(new_n624), .A2(KEYINPUT32), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n290), .A2(new_n291), .A3(new_n292), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n644), .B1(new_n658), .B2(new_n283), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n486), .A2(new_n487), .ZN(new_n660));
  INV_X1    g474(.A(new_n611), .ZN(new_n661));
  INV_X1    g475(.A(G900), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n492), .B1(new_n494), .B2(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n583), .A2(new_n663), .ZN(new_n664));
  AND2_X1   g478(.A1(new_n664), .A2(new_n539), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n659), .A2(new_n660), .A3(new_n661), .A4(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G128), .ZN(G30));
  XNOR2_X1  g481(.A(new_n663), .B(KEYINPUT39), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n617), .A2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  OR2_X1    g484(.A1(new_n670), .A2(KEYINPUT40), .ZN(new_n671));
  INV_X1    g485(.A(new_n276), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n672), .A2(new_n266), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n243), .A2(new_n245), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n341), .B1(new_n674), .B2(new_n284), .ZN(new_n675));
  OAI21_X1  g489(.A(G472), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  AND2_X1   g490(.A1(new_n658), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n584), .A2(new_n588), .ZN(new_n678));
  INV_X1    g492(.A(new_n422), .ZN(new_n679));
  NOR4_X1   g493(.A1(new_n677), .A2(new_n633), .A3(new_n678), .A4(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n670), .A2(KEYINPUT40), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n421), .A2(new_n423), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(KEYINPUT38), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n683), .A2(new_n650), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n671), .A2(new_n680), .A3(new_n681), .A4(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(KEYINPUT102), .B(G143), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(G45));
  AND4_X1   g501(.A1(new_n295), .A2(new_n615), .A3(new_n616), .A4(new_n650), .ZN(new_n688));
  INV_X1    g502(.A(new_n663), .ZN(new_n689));
  AND4_X1   g503(.A1(new_n584), .A2(new_n603), .A3(new_n588), .A4(new_n689), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n688), .A2(KEYINPUT103), .A3(new_n661), .A4(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n659), .A2(new_n660), .A3(new_n661), .A4(new_n690), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT103), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G146), .ZN(G48));
  NOR2_X1   g510(.A1(new_n466), .A2(new_n470), .ZN(new_n697));
  OAI21_X1  g511(.A(G469), .B1(new_n697), .B2(G902), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n698), .A2(new_n485), .A3(new_n471), .ZN(new_n699));
  AOI211_X1 g513(.A(new_n352), .B(new_n699), .C1(new_n658), .C2(new_n283), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n700), .A2(new_n612), .A3(new_n606), .A4(new_n608), .ZN(new_n701));
  XOR2_X1   g515(.A(KEYINPUT41), .B(G113), .Z(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(KEYINPUT104), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n701), .B(new_n703), .ZN(G15));
  NAND2_X1  g518(.A1(new_n700), .A2(new_n634), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G116), .ZN(G18));
  NOR2_X1   g520(.A1(new_n611), .A2(new_n699), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n659), .A2(new_n589), .A3(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G119), .ZN(G21));
  AOI21_X1  g523(.A(new_n679), .B1(new_n536), .B2(new_n538), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n584), .A2(new_n710), .A3(new_n588), .A4(new_n610), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n711), .A2(new_n498), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n352), .A2(KEYINPUT107), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT107), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n714), .B1(new_n349), .B2(new_n351), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(new_n699), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT106), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n718), .B1(new_n619), .B2(new_n620), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n625), .A2(KEYINPUT106), .A3(G472), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n266), .B1(new_n246), .B2(new_n249), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(new_n288), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n292), .B1(new_n622), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(KEYINPUT105), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT105), .ZN(new_n725));
  OAI211_X1 g539(.A(new_n725), .B(new_n292), .C1(new_n622), .C2(new_n722), .ZN(new_n726));
  AOI22_X1  g540(.A1(new_n719), .A2(new_n720), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n712), .A2(new_n716), .A3(new_n717), .A4(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G122), .ZN(G24));
  NAND4_X1  g543(.A1(new_n727), .A2(new_n690), .A3(new_n650), .A4(new_n707), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G125), .ZN(G27));
  AOI21_X1  g545(.A(new_n679), .B1(new_n421), .B2(new_n423), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n613), .A2(KEYINPUT108), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT108), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n481), .A2(new_n734), .A3(new_n485), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n732), .A2(new_n733), .A3(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT109), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n732), .A2(new_n733), .A3(KEYINPUT109), .A4(new_n735), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT110), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n741), .B1(new_n293), .B2(new_n294), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n656), .A2(KEYINPUT110), .A3(new_n657), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n742), .A2(new_n283), .A3(new_n743), .ZN(new_n744));
  AND2_X1   g558(.A1(new_n744), .A2(new_n716), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n740), .A2(KEYINPUT42), .A3(new_n690), .A4(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(new_n690), .ZN(new_n747));
  AOI211_X1 g561(.A(new_n354), .B(new_n747), .C1(new_n738), .C2(new_n739), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n746), .B1(new_n748), .B2(KEYINPUT42), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G131), .ZN(G33));
  AND3_X1   g564(.A1(new_n481), .A2(new_n734), .A3(new_n485), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n734), .B1(new_n481), .B2(new_n485), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  AOI21_X1  g567(.A(KEYINPUT109), .B1(new_n753), .B2(new_n732), .ZN(new_n754));
  AND4_X1   g568(.A1(KEYINPUT109), .A2(new_n732), .A3(new_n733), .A4(new_n735), .ZN(new_n755));
  OAI211_X1 g569(.A(new_n355), .B(new_n665), .C1(new_n754), .C2(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT111), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n740), .A2(KEYINPUT111), .A3(new_n355), .A4(new_n665), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G134), .ZN(G36));
  AOI22_X1  g575(.A1(new_n448), .A2(new_n458), .B1(new_n461), .B2(new_n464), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n474), .B1(new_n762), .B2(new_n473), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(new_n477), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT45), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n763), .A2(KEYINPUT45), .A3(new_n477), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n766), .A2(G469), .A3(new_n767), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n768), .A2(KEYINPUT46), .A3(new_n480), .ZN(new_n769));
  AOI21_X1  g583(.A(KEYINPUT46), .B1(new_n768), .B2(new_n480), .ZN(new_n770));
  INV_X1    g584(.A(new_n471), .ZN(new_n771));
  NOR3_X1   g585(.A1(new_n769), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n772), .A2(new_n484), .ZN(new_n773));
  INV_X1    g587(.A(new_n668), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(KEYINPUT112), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT112), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n773), .A2(new_n777), .A3(new_n774), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(new_n732), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n678), .A2(new_n603), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT43), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n678), .A2(KEYINPUT43), .A3(new_n603), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n785), .A2(new_n628), .A3(new_n650), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n780), .B1(new_n787), .B2(KEYINPUT44), .ZN(new_n788));
  OAI211_X1 g602(.A(new_n779), .B(new_n788), .C1(KEYINPUT44), .C2(new_n787), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G137), .ZN(G39));
  NAND2_X1  g604(.A1(new_n773), .A2(KEYINPUT47), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT47), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n792), .B1(new_n772), .B2(new_n484), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n780), .A2(new_n295), .A3(new_n353), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n794), .A2(new_n690), .A3(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G140), .ZN(G42));
  AOI21_X1  g611(.A(new_n493), .B1(new_n783), .B2(new_n784), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n780), .A2(new_n699), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n727), .A2(new_n650), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n352), .A2(new_n493), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n799), .A2(new_n677), .A3(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n678), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n804), .A2(new_n805), .A3(new_n603), .ZN(new_n806));
  OR2_X1    g620(.A1(new_n802), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n716), .A2(new_n727), .ZN(new_n808));
  INV_X1    g622(.A(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n798), .A2(new_n809), .A3(new_n679), .ZN(new_n810));
  INV_X1    g624(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n683), .A2(new_n717), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  AOI21_X1  g627(.A(KEYINPUT50), .B1(new_n811), .B2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT50), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n810), .A2(new_n816), .A3(new_n812), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n807), .B1(new_n815), .B2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(new_n698), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n820), .A2(new_n771), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(new_n484), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n791), .A2(new_n793), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(KEYINPUT116), .ZN(new_n824));
  AND3_X1   g638(.A1(new_n798), .A2(new_n809), .A3(new_n732), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT116), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n791), .A2(new_n826), .A3(new_n793), .A4(new_n822), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n824), .A2(new_n825), .A3(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n819), .A2(KEYINPUT51), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(KEYINPUT117), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT117), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n819), .A2(new_n828), .A3(new_n831), .A4(KEYINPUT51), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n823), .A2(new_n825), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n802), .A2(new_n806), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n834), .B(new_n835), .C1(new_n814), .C2(new_n817), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT51), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(KEYINPUT115), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT115), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n836), .A2(new_n840), .A3(new_n837), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n798), .A2(new_n809), .A3(new_n707), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(new_n490), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n798), .A2(new_n745), .A3(new_n799), .ZN(new_n844));
  OR2_X1    g658(.A1(new_n844), .A2(KEYINPUT48), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(KEYINPUT48), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n843), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT118), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n609), .A2(new_n677), .A3(new_n799), .A4(new_n803), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n847), .A2(new_n849), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(KEYINPUT118), .ZN(new_n852));
  AOI22_X1  g666(.A1(new_n839), .A2(new_n841), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n604), .B1(new_n805), .B2(new_n633), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n424), .A2(new_n498), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n629), .A2(new_n353), .A3(new_n854), .A4(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n652), .A2(new_n856), .A3(new_n590), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n701), .A2(new_n705), .A3(new_n708), .A4(new_n728), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n732), .A2(new_n633), .A3(new_n664), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n860), .B(KEYINPUT113), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n801), .A2(new_n747), .ZN(new_n862));
  AOI22_X1  g676(.A1(new_n861), .A2(new_n688), .B1(new_n862), .B2(new_n740), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n859), .A2(new_n760), .A3(new_n749), .A4(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n666), .A2(new_n730), .ZN(new_n866));
  INV_X1    g680(.A(new_n866), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n677), .A2(new_n650), .A3(new_n663), .ZN(new_n868));
  INV_X1    g682(.A(new_n711), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n868), .A2(new_n485), .A3(new_n481), .A4(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n695), .A2(new_n867), .A3(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT52), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n866), .B1(new_n694), .B2(new_n691), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n874), .A2(KEYINPUT52), .A3(new_n870), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n865), .A2(KEYINPUT53), .A3(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT53), .ZN(new_n878));
  AND4_X1   g692(.A1(KEYINPUT52), .A2(new_n695), .A3(new_n867), .A4(new_n870), .ZN(new_n879));
  XNOR2_X1  g693(.A(KEYINPUT114), .B(KEYINPUT52), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n880), .B1(new_n874), .B2(new_n870), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n878), .B1(new_n882), .B2(new_n864), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n877), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(KEYINPUT54), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT54), .ZN(new_n886));
  INV_X1    g700(.A(new_n871), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n875), .B1(new_n887), .B2(new_n880), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n878), .B1(new_n865), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(KEYINPUT52), .B1(new_n874), .B2(new_n870), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n879), .A2(new_n890), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n891), .A2(new_n864), .A3(KEYINPUT53), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n886), .B1(new_n889), .B2(new_n892), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n833), .A2(new_n853), .A3(new_n885), .A4(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(KEYINPUT119), .ZN(new_n895));
  OAI21_X1  g709(.A(KEYINPUT53), .B1(new_n882), .B2(new_n864), .ZN(new_n896));
  AND2_X1   g710(.A1(new_n760), .A2(new_n749), .ZN(new_n897));
  INV_X1    g711(.A(new_n857), .ZN(new_n898));
  INV_X1    g712(.A(new_n858), .ZN(new_n899));
  AND3_X1   g713(.A1(new_n898), .A2(new_n899), .A3(new_n863), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n876), .A2(new_n897), .A3(new_n878), .A4(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(KEYINPUT54), .B1(new_n896), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n902), .B1(KEYINPUT54), .B2(new_n884), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT119), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n903), .A2(new_n904), .A3(new_n833), .A4(new_n853), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n489), .A2(new_n398), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n895), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n683), .A2(new_n678), .A3(new_n603), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n821), .B(KEYINPUT49), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n909), .A2(new_n677), .A3(new_n716), .ZN(new_n910));
  OR4_X1    g724(.A1(new_n484), .A2(new_n908), .A3(new_n910), .A4(new_n679), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n907), .A2(new_n911), .ZN(G75));
  NAND4_X1  g726(.A1(new_n896), .A2(new_n901), .A3(G210), .A4(G902), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT56), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n913), .A2(KEYINPUT120), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n390), .A2(new_n392), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n916), .B(new_n400), .Z(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT55), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  OR2_X1    g733(.A1(new_n915), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n251), .A2(G952), .ZN(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(KEYINPUT120), .B1(new_n913), .B2(new_n914), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n919), .B1(new_n915), .B2(new_n923), .ZN(new_n924));
  AND3_X1   g738(.A1(new_n920), .A2(new_n922), .A3(new_n924), .ZN(G51));
  NAND2_X1  g739(.A1(new_n896), .A2(new_n901), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n926), .A2(new_n341), .A3(new_n768), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n480), .B(KEYINPUT57), .Z(new_n928));
  AND3_X1   g742(.A1(new_n896), .A2(KEYINPUT54), .A3(new_n901), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n928), .B1(new_n929), .B2(new_n902), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n697), .B(KEYINPUT121), .Z(new_n931));
  AOI21_X1  g745(.A(new_n927), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g746(.A(KEYINPUT122), .B1(new_n932), .B2(new_n921), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT122), .ZN(new_n934));
  INV_X1    g748(.A(new_n931), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n896), .A2(KEYINPUT54), .A3(new_n901), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n893), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n935), .B1(new_n937), .B2(new_n928), .ZN(new_n938));
  OAI211_X1 g752(.A(new_n934), .B(new_n922), .C1(new_n938), .C2(new_n927), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n933), .A2(new_n939), .ZN(G54));
  NOR2_X1   g754(.A1(new_n889), .A2(new_n892), .ZN(new_n941));
  NAND2_X1  g755(.A1(KEYINPUT58), .A2(G475), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(KEYINPUT123), .ZN(new_n943));
  OR2_X1    g757(.A1(new_n942), .A2(KEYINPUT123), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n941), .A2(G902), .A3(new_n943), .A4(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n570), .ZN(new_n946));
  AND2_X1   g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n945), .A2(new_n946), .ZN(new_n948));
  NOR3_X1   g762(.A1(new_n947), .A2(new_n948), .A3(new_n921), .ZN(G60));
  NAND2_X1  g763(.A1(G478), .A2(G902), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n950), .B(KEYINPUT59), .Z(new_n951));
  OAI21_X1  g765(.A(new_n601), .B1(new_n903), .B2(new_n951), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n601), .A2(new_n951), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n937), .A2(new_n953), .ZN(new_n954));
  AND3_X1   g768(.A1(new_n952), .A2(new_n922), .A3(new_n954), .ZN(G63));
  NAND2_X1  g769(.A1(G217), .A2(G902), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n956), .B(KEYINPUT60), .Z(new_n957));
  NAND2_X1  g771(.A1(new_n941), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n340), .A2(new_n342), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT124), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n960), .A2(new_n961), .A3(new_n922), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n941), .B(new_n957), .C1(new_n641), .C2(new_n642), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n960), .A2(new_n922), .A3(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT61), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n962), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n921), .B1(new_n958), .B2(new_n959), .ZN(new_n967));
  OAI211_X1 g781(.A(new_n967), .B(new_n963), .C1(new_n961), .C2(KEYINPUT61), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n966), .A2(new_n968), .ZN(G66));
  AOI21_X1  g783(.A(new_n398), .B1(new_n496), .B2(G224), .ZN(new_n970));
  INV_X1    g784(.A(new_n859), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n970), .B1(new_n971), .B2(new_n251), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n916), .B1(G898), .B2(new_n251), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n972), .B(new_n973), .Z(G69));
  AND2_X1   g788(.A1(new_n789), .A2(new_n796), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n779), .A2(new_n869), .A3(new_n745), .ZN(new_n976));
  AND2_X1   g790(.A1(new_n976), .A2(new_n874), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n975), .A2(new_n977), .A3(new_n251), .A4(new_n897), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n978), .B1(new_n662), .B2(new_n251), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n270), .B1(new_n272), .B2(new_n274), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n980), .B(KEYINPUT125), .Z(new_n981));
  XOR2_X1   g795(.A(new_n981), .B(new_n565), .Z(new_n982));
  NAND2_X1  g796(.A1(new_n979), .A2(new_n982), .ZN(new_n983));
  NAND4_X1  g797(.A1(new_n669), .A2(new_n355), .A3(new_n854), .A4(new_n732), .ZN(new_n984));
  AOI21_X1  g798(.A(KEYINPUT62), .B1(new_n685), .B2(new_n874), .ZN(new_n985));
  AND3_X1   g799(.A1(new_n685), .A2(KEYINPUT62), .A3(new_n874), .ZN(new_n986));
  OAI211_X1 g800(.A(new_n975), .B(new_n984), .C1(new_n985), .C2(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(new_n982), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n987), .A2(new_n251), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n983), .A2(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(new_n251), .ZN(new_n991));
  NAND2_X1  g805(.A1(G227), .A2(G900), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n990), .B(new_n993), .ZN(G72));
  NAND4_X1  g808(.A1(new_n975), .A2(new_n977), .A3(new_n897), .A4(new_n859), .ZN(new_n995));
  NAND2_X1  g809(.A1(G472), .A2(G902), .ZN(new_n996));
  XOR2_X1   g810(.A(new_n996), .B(KEYINPUT63), .Z(new_n997));
  XNOR2_X1  g811(.A(new_n997), .B(KEYINPUT126), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n995), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n284), .B1(new_n999), .B2(KEYINPUT127), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT127), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n995), .A2(new_n1001), .A3(new_n998), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n1000), .A2(new_n672), .A3(new_n1002), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n998), .B1(new_n987), .B2(new_n971), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n921), .B1(new_n1004), .B2(new_n673), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n277), .A2(new_n285), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n884), .A2(new_n997), .A3(new_n1006), .ZN(new_n1007));
  AND3_X1   g821(.A1(new_n1003), .A2(new_n1005), .A3(new_n1007), .ZN(G57));
endmodule


