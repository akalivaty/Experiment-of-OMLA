//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 1 1 1 0 1 0 1 0 1 1 1 0 0 1 0 1 1 0 1 1 1 1 0 1 1 1 0 1 1 1 0 1 0 0 1 1 1 0 0 0 1 0 1 0 1 1 0 1 1 1 1 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:35 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n435, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n563, new_n565,
    new_n566, new_n567, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n599, new_n600, new_n601, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n625, new_n626, new_n627, new_n628, new_n629, new_n632,
    new_n634, new_n635, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n853, new_n854, new_n855, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1199, new_n1200, new_n1201;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT65), .B(G132), .Z(new_n435));
  INV_X1    g010(.A(new_n435), .ZN(G219));
  XNOR2_X1  g011(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT66), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G219), .A2(G218), .A3(G221), .A4(G220), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2104), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(KEYINPUT3), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n460), .A2(new_n462), .A3(G125), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT67), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT67), .ZN(new_n465));
  NAND4_X1  g040(.A1(new_n460), .A2(new_n462), .A3(new_n465), .A4(G125), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n464), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  OAI21_X1  g044(.A(KEYINPUT68), .B1(new_n459), .B2(KEYINPUT3), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(new_n460), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n459), .A2(KEYINPUT68), .A3(KEYINPUT3), .ZN(new_n473));
  NAND4_X1  g048(.A1(new_n471), .A2(G137), .A3(new_n472), .A4(new_n473), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n472), .A2(G101), .A3(G2104), .ZN(new_n475));
  AND2_X1   g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AND2_X1   g051(.A1(new_n469), .A2(new_n476), .ZN(G160));
  AND2_X1   g052(.A1(new_n471), .A2(new_n473), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(new_n472), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT69), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n478), .A2(KEYINPUT69), .A3(new_n472), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(G100), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n484), .A2(new_n472), .A3(KEYINPUT71), .ZN(new_n485));
  AOI21_X1  g060(.A(KEYINPUT71), .B1(new_n484), .B2(new_n472), .ZN(new_n486));
  OAI21_X1  g061(.A(G2104), .B1(new_n472), .B2(G112), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  AOI22_X1  g063(.A1(new_n483), .A2(G136), .B1(new_n485), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n478), .A2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT70), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n478), .A2(KEYINPUT70), .A3(G2105), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G124), .ZN(new_n495));
  AND2_X1   g070(.A1(new_n489), .A2(new_n495), .ZN(G162));
  NAND2_X1  g071(.A1(new_n460), .A2(new_n462), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n498), .A2(new_n472), .A3(G138), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n471), .A2(G138), .A3(new_n472), .A4(new_n473), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n500), .B1(new_n501), .B2(KEYINPUT4), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n471), .A2(G126), .A3(G2105), .A4(new_n473), .ZN(new_n503));
  OR2_X1    g078(.A1(G102), .A2(G2105), .ZN(new_n504));
  OAI211_X1 g079(.A(new_n504), .B(G2104), .C1(G114), .C2(new_n472), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n502), .A2(new_n506), .ZN(G164));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(KEYINPUT6), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT6), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G651), .ZN(new_n511));
  AND2_X1   g086(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G50), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT5), .B(G543), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n515), .A2(new_n509), .A3(new_n511), .ZN(new_n516));
  INV_X1    g091(.A(G88), .ZN(new_n517));
  OAI22_X1  g092(.A1(new_n513), .A2(new_n514), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n515), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n519), .A2(new_n508), .ZN(new_n520));
  OR2_X1    g095(.A1(new_n518), .A2(new_n520), .ZN(G303));
  INV_X1    g096(.A(G303), .ZN(G166));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n523), .B(KEYINPUT7), .ZN(new_n524));
  INV_X1    g099(.A(G89), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n524), .B1(new_n516), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(KEYINPUT72), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT72), .ZN(new_n528));
  OAI211_X1 g103(.A(new_n528), .B(new_n524), .C1(new_n516), .C2(new_n525), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n509), .A2(new_n511), .ZN(new_n531));
  INV_X1    g106(.A(G543), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AND2_X1   g108(.A1(G63), .A2(G651), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n533), .A2(G51), .B1(new_n515), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n530), .A2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT73), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n530), .A2(KEYINPUT73), .A3(new_n535), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(new_n539), .ZN(G168));
  INV_X1    g115(.A(G52), .ZN(new_n541));
  INV_X1    g116(.A(G90), .ZN(new_n542));
  OAI22_X1  g117(.A1(new_n513), .A2(new_n541), .B1(new_n516), .B2(new_n542), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n515), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n544), .A2(new_n508), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n543), .A2(new_n545), .ZN(G171));
  NAND2_X1  g121(.A1(G68), .A2(G543), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n532), .A2(KEYINPUT5), .ZN(new_n548));
  INV_X1    g123(.A(KEYINPUT5), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G543), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(G56), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n547), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G651), .ZN(new_n554));
  OR2_X1    g129(.A1(new_n554), .A2(KEYINPUT74), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n554), .A2(KEYINPUT74), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n551), .A2(new_n531), .ZN(new_n557));
  AOI22_X1  g132(.A1(G81), .A2(new_n557), .B1(new_n533), .B2(G43), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n555), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT75), .ZN(G153));
  AND3_X1   g137(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G36), .ZN(G176));
  NAND2_X1  g139(.A1(G1), .A2(G3), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT8), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  XOR2_X1   g142(.A(new_n567), .B(KEYINPUT76), .Z(G188));
  INV_X1    g143(.A(G53), .ZN(new_n569));
  OAI211_X1 g144(.A(KEYINPUT77), .B(KEYINPUT9), .C1(new_n513), .C2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(KEYINPUT77), .A2(KEYINPUT9), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n533), .A2(G53), .A3(new_n571), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n570), .A2(new_n572), .B1(G91), .B2(new_n557), .ZN(new_n573));
  NAND2_X1  g148(.A1(G78), .A2(G543), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT78), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n515), .B(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(G65), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n574), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT79), .ZN(new_n579));
  AND3_X1   g154(.A1(new_n578), .A2(new_n579), .A3(G651), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n579), .B1(new_n578), .B2(G651), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n573), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT80), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI211_X1 g159(.A(KEYINPUT80), .B(new_n573), .C1(new_n580), .C2(new_n581), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(G299));
  INV_X1    g161(.A(G171), .ZN(G301));
  INV_X1    g162(.A(G168), .ZN(G286));
  OAI21_X1  g163(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT81), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n589), .B(new_n590), .ZN(new_n591));
  AOI22_X1  g166(.A1(G87), .A2(new_n557), .B1(new_n533), .B2(G49), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n593), .A2(KEYINPUT82), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT82), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n595), .B1(new_n591), .B2(new_n592), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(G288));
  NAND3_X1  g173(.A1(new_n512), .A2(G86), .A3(new_n515), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n512), .A2(G48), .A3(G543), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n515), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n601));
  OAI211_X1 g176(.A(new_n599), .B(new_n600), .C1(new_n601), .C2(new_n508), .ZN(G305));
  AOI22_X1  g177(.A1(G85), .A2(new_n557), .B1(new_n533), .B2(G47), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n508), .B2(new_n604), .ZN(G290));
  NAND2_X1  g180(.A1(G301), .A2(G868), .ZN(new_n606));
  INV_X1    g181(.A(G66), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n576), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(G79), .A2(G543), .ZN(new_n609));
  XOR2_X1   g184(.A(new_n609), .B(KEYINPUT84), .Z(new_n610));
  OAI21_X1  g185(.A(G651), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n533), .A2(KEYINPUT83), .ZN(new_n612));
  INV_X1    g187(.A(G54), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT83), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n613), .B1(new_n513), .B2(new_n614), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n557), .A2(KEYINPUT10), .A3(G92), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT10), .ZN(new_n617));
  INV_X1    g192(.A(G92), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n516), .B2(new_n618), .ZN(new_n619));
  AOI22_X1  g194(.A1(new_n612), .A2(new_n615), .B1(new_n616), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n611), .A2(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(new_n621), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n606), .B1(new_n622), .B2(G868), .ZN(G284));
  OAI21_X1  g198(.A(new_n606), .B1(new_n622), .B2(G868), .ZN(G321));
  INV_X1    g199(.A(KEYINPUT85), .ZN(new_n625));
  INV_X1    g200(.A(G868), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(G168), .B2(new_n626), .ZN(new_n627));
  NOR2_X1   g202(.A1(G168), .A2(new_n626), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n628), .B1(G299), .B2(new_n626), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n627), .B1(new_n629), .B2(new_n625), .ZN(G297));
  OAI21_X1  g205(.A(new_n627), .B1(new_n629), .B2(new_n625), .ZN(G280));
  INV_X1    g206(.A(G559), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n622), .B1(new_n632), .B2(G860), .ZN(G148));
  NAND2_X1  g208(.A1(new_n559), .A2(new_n626), .ZN(new_n634));
  NOR2_X1   g209(.A1(new_n621), .A2(G559), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n634), .B1(new_n635), .B2(new_n626), .ZN(G323));
  XNOR2_X1  g211(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g212(.A1(new_n494), .A2(G123), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n483), .A2(G135), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n472), .A2(G111), .ZN(new_n640));
  OAI21_X1  g215(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n641));
  OAI211_X1 g216(.A(new_n638), .B(new_n639), .C1(new_n640), .C2(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(KEYINPUT89), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2096), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT86), .B(KEYINPUT12), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT87), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n472), .A2(G2104), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n497), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n646), .B(new_n648), .Z(new_n649));
  XOR2_X1   g224(.A(KEYINPUT88), .B(G2100), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT13), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n649), .B(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n644), .A2(new_n652), .ZN(G156));
  XOR2_X1   g228(.A(KEYINPUT15), .B(G2435), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2438), .ZN(new_n655));
  XOR2_X1   g230(.A(G2427), .B(G2430), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT90), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n655), .A2(new_n657), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n658), .A2(new_n659), .A3(KEYINPUT14), .ZN(new_n660));
  XOR2_X1   g235(.A(KEYINPUT91), .B(KEYINPUT16), .Z(new_n661));
  XNOR2_X1  g236(.A(G2451), .B(G2454), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n660), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2443), .B(G2446), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1341), .B(G1348), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n666), .A2(new_n667), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n668), .A2(G14), .A3(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(KEYINPUT92), .Z(G401));
  XOR2_X1   g246(.A(G2084), .B(G2090), .Z(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G2067), .B(G2678), .Z(new_n674));
  NOR2_X1   g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G2072), .B(G2078), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT18), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n673), .A2(new_n674), .ZN(new_n679));
  AND3_X1   g254(.A1(new_n679), .A2(KEYINPUT17), .A3(new_n676), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n676), .B1(new_n679), .B2(KEYINPUT17), .ZN(new_n681));
  NOR3_X1   g256(.A1(new_n680), .A2(new_n681), .A3(new_n675), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G2096), .B(G2100), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(G227));
  XOR2_X1   g260(.A(G1956), .B(G2474), .Z(new_n686));
  XOR2_X1   g261(.A(G1961), .B(G1966), .Z(new_n687));
  AND2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n686), .A2(new_n687), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1971), .B(G1976), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT19), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n689), .A2(new_n691), .A3(new_n693), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n689), .A2(new_n693), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(KEYINPUT20), .ZN(new_n697));
  OAI221_X1 g272(.A(new_n694), .B1(new_n693), .B2(new_n691), .C1(new_n696), .C2(new_n697), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n698), .B1(new_n697), .B2(new_n696), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT94), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1991), .B(G1996), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT93), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(G1981), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(G1986), .Z(new_n704));
  XNOR2_X1  g279(.A(new_n700), .B(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n706));
  OR2_X1    g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n705), .A2(new_n706), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n707), .A2(new_n708), .ZN(G229));
  INV_X1    g284(.A(KEYINPUT96), .ZN(new_n710));
  AND2_X1   g285(.A1(KEYINPUT95), .A2(G16), .ZN(new_n711));
  NOR2_X1   g286(.A1(KEYINPUT95), .A2(G16), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(G22), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n710), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n713), .A2(new_n714), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(G303), .B2(new_n713), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n715), .B1(new_n717), .B2(new_n710), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(G1971), .ZN(new_n719));
  INV_X1    g294(.A(new_n593), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(G16), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G16), .B2(G23), .ZN(new_n722));
  XOR2_X1   g297(.A(KEYINPUT33), .B(G1976), .Z(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  OAI211_X1 g300(.A(new_n721), .B(new_n723), .C1(G16), .C2(G23), .ZN(new_n726));
  MUX2_X1   g301(.A(G6), .B(G305), .S(G16), .Z(new_n727));
  XOR2_X1   g302(.A(KEYINPUT32), .B(G1981), .Z(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n725), .A2(new_n726), .A3(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT34), .ZN(new_n731));
  OR3_X1    g306(.A1(new_n719), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n731), .B1(new_n719), .B2(new_n730), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(G29), .ZN(new_n735));
  AND2_X1   g310(.A1(new_n735), .A2(G25), .ZN(new_n736));
  OAI21_X1  g311(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n737));
  INV_X1    g312(.A(G107), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n737), .B1(new_n738), .B2(G2105), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(new_n483), .B2(G131), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n494), .A2(G119), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n736), .B1(new_n742), .B2(G29), .ZN(new_n743));
  XOR2_X1   g318(.A(KEYINPUT35), .B(G1991), .Z(new_n744));
  AND2_X1   g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n743), .A2(new_n744), .ZN(new_n746));
  MUX2_X1   g321(.A(G24), .B(G290), .S(new_n713), .Z(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(G1986), .ZN(new_n748));
  NOR3_X1   g323(.A1(new_n745), .A2(new_n746), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n734), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n750), .A2(KEYINPUT97), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT97), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n734), .A2(new_n752), .A3(new_n749), .ZN(new_n753));
  AND3_X1   g328(.A1(new_n751), .A2(KEYINPUT36), .A3(new_n753), .ZN(new_n754));
  AOI21_X1  g329(.A(KEYINPUT36), .B1(new_n751), .B2(new_n753), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g331(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(KEYINPUT99), .Z(new_n758));
  NOR2_X1   g333(.A1(new_n459), .A2(G2105), .ZN(new_n759));
  AOI22_X1  g334(.A1(new_n758), .A2(KEYINPUT26), .B1(G105), .B2(new_n759), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(KEYINPUT26), .B2(new_n758), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(new_n483), .B2(G141), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n494), .A2(G129), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(KEYINPUT100), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n766), .A2(G29), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G29), .B2(G32), .ZN(new_n768));
  XNOR2_X1  g343(.A(KEYINPUT27), .B(G1996), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT101), .Z(new_n770));
  NAND2_X1  g345(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT30), .B(G28), .ZN(new_n772));
  AND2_X1   g347(.A1(new_n772), .A2(new_n735), .ZN(new_n773));
  XOR2_X1   g348(.A(KEYINPUT31), .B(G11), .Z(new_n774));
  NAND2_X1  g349(.A1(G171), .A2(G16), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G5), .B2(G16), .ZN(new_n776));
  INV_X1    g351(.A(G1961), .ZN(new_n777));
  AOI211_X1 g352(.A(new_n773), .B(new_n774), .C1(new_n776), .C2(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n622), .A2(G16), .ZN(new_n779));
  INV_X1    g354(.A(G1348), .ZN(new_n780));
  OR2_X1    g355(.A1(G4), .A2(G16), .ZN(new_n781));
  AND3_X1   g356(.A1(new_n779), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n780), .B1(new_n779), .B2(new_n781), .ZN(new_n783));
  OAI221_X1 g358(.A(new_n778), .B1(new_n777), .B2(new_n776), .C1(new_n782), .C2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n735), .A2(G27), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G164), .B2(new_n735), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(G2078), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n784), .A2(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(new_n770), .ZN(new_n789));
  OAI211_X1 g364(.A(new_n767), .B(new_n789), .C1(G29), .C2(G32), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n643), .A2(G29), .ZN(new_n791));
  NAND4_X1  g366(.A1(new_n771), .A2(new_n788), .A3(new_n790), .A4(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n735), .A2(G35), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G162), .B2(new_n735), .ZN(new_n794));
  XNOR2_X1  g369(.A(KEYINPUT29), .B(G2090), .ZN(new_n795));
  INV_X1    g370(.A(new_n795), .ZN(new_n796));
  OR2_X1    g371(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n794), .A2(new_n796), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n483), .A2(G139), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n759), .A2(G103), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT25), .ZN(new_n801));
  NAND2_X1  g376(.A1(G115), .A2(G2104), .ZN(new_n802));
  INV_X1    g377(.A(G127), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n802), .B1(new_n497), .B2(new_n803), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n801), .B1(G2105), .B2(new_n804), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n799), .A2(G29), .A3(new_n805), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(G29), .B2(G33), .ZN(new_n807));
  INV_X1    g382(.A(G2072), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n809), .A2(KEYINPUT98), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(KEYINPUT98), .ZN(new_n811));
  AOI22_X1  g386(.A1(new_n797), .A2(new_n798), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(G16), .A2(G21), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(G168), .B2(G16), .ZN(new_n814));
  INV_X1    g389(.A(G1966), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  MUX2_X1   g391(.A(G19), .B(new_n559), .S(new_n713), .Z(new_n817));
  INV_X1    g392(.A(G1341), .ZN(new_n818));
  AND2_X1   g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n817), .A2(new_n818), .ZN(new_n820));
  OAI22_X1  g395(.A1(new_n819), .A2(new_n820), .B1(new_n807), .B2(new_n808), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT24), .ZN(new_n822));
  INV_X1    g397(.A(G34), .ZN(new_n823));
  AOI21_X1  g398(.A(G29), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(new_n822), .B2(new_n823), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(G160), .B2(new_n735), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(G2084), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n821), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n812), .A2(new_n816), .A3(new_n828), .ZN(new_n829));
  OAI21_X1  g404(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n830));
  INV_X1    g405(.A(G116), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n830), .B1(new_n831), .B2(G2105), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n832), .B1(new_n483), .B2(G140), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n494), .A2(G128), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(new_n835), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n836), .A2(new_n735), .ZN(new_n837));
  AND2_X1   g412(.A1(new_n735), .A2(G26), .ZN(new_n838));
  OAI21_X1  g413(.A(KEYINPUT28), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n838), .A2(KEYINPUT28), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(G2067), .ZN(new_n842));
  NOR3_X1   g417(.A1(new_n792), .A2(new_n829), .A3(new_n842), .ZN(new_n843));
  OAI21_X1  g418(.A(G20), .B1(new_n711), .B2(new_n712), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(KEYINPUT23), .Z(new_n845));
  AOI21_X1  g420(.A(new_n845), .B1(G299), .B2(G16), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT102), .ZN(new_n847));
  INV_X1    g422(.A(G1956), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n847), .B(new_n848), .ZN(new_n849));
  AND3_X1   g424(.A1(new_n843), .A2(new_n849), .A3(KEYINPUT103), .ZN(new_n850));
  AOI21_X1  g425(.A(KEYINPUT103), .B1(new_n843), .B2(new_n849), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n756), .B1(new_n850), .B2(new_n851), .ZN(G150));
  INV_X1    g427(.A(KEYINPUT104), .ZN(new_n853));
  NAND2_X1  g428(.A1(G150), .A2(new_n853), .ZN(new_n854));
  OAI211_X1 g429(.A(new_n756), .B(KEYINPUT104), .C1(new_n850), .C2(new_n851), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(G311));
  NOR2_X1   g431(.A1(new_n621), .A2(new_n632), .ZN(new_n857));
  XNOR2_X1  g432(.A(KEYINPUT106), .B(KEYINPUT38), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n857), .B(new_n858), .ZN(new_n859));
  AOI22_X1  g434(.A1(new_n515), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n860));
  OR2_X1    g435(.A1(new_n860), .A2(new_n508), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n557), .A2(G93), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n533), .A2(G55), .ZN(new_n863));
  AND3_X1   g438(.A1(new_n862), .A2(KEYINPUT105), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(KEYINPUT105), .B1(new_n862), .B2(new_n863), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n861), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(new_n559), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n859), .B(new_n868), .ZN(new_n869));
  OR2_X1    g444(.A1(new_n869), .A2(KEYINPUT39), .ZN(new_n870));
  OR2_X1    g445(.A1(new_n870), .A2(KEYINPUT107), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(KEYINPUT107), .ZN(new_n872));
  AOI21_X1  g447(.A(G860), .B1(new_n869), .B2(KEYINPUT39), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n871), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  XOR2_X1   g449(.A(new_n874), .B(KEYINPUT108), .Z(new_n875));
  NAND2_X1  g450(.A1(new_n866), .A2(G860), .ZN(new_n876));
  XOR2_X1   g451(.A(KEYINPUT109), .B(KEYINPUT37), .Z(new_n877));
  XNOR2_X1  g452(.A(new_n876), .B(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n875), .A2(new_n878), .ZN(G145));
  XOR2_X1   g454(.A(new_n643), .B(G160), .Z(new_n880));
  INV_X1    g455(.A(G162), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n880), .B(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n766), .A2(new_n799), .A3(new_n805), .ZN(new_n884));
  XOR2_X1   g459(.A(new_n835), .B(G164), .Z(new_n885));
  NAND2_X1  g460(.A1(new_n799), .A2(new_n805), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n764), .A2(new_n886), .ZN(new_n887));
  AND3_X1   g462(.A1(new_n884), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n885), .B1(new_n884), .B2(new_n887), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n494), .A2(G130), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n483), .A2(G142), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n472), .A2(G118), .ZN(new_n893));
  OAI21_X1  g468(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n894));
  OAI211_X1 g469(.A(new_n891), .B(new_n892), .C1(new_n893), .C2(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(new_n742), .ZN(new_n896));
  XOR2_X1   g471(.A(new_n896), .B(new_n649), .Z(new_n897));
  OR2_X1    g472(.A1(new_n890), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n890), .A2(new_n897), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(G37), .B1(new_n883), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n899), .A2(KEYINPUT110), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT110), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n890), .A2(new_n903), .A3(new_n897), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n882), .A2(new_n902), .A3(new_n904), .A4(new_n898), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n901), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(KEYINPUT40), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT40), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n901), .A2(new_n908), .A3(new_n905), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n907), .A2(new_n909), .ZN(G395));
  NAND3_X1  g485(.A1(new_n584), .A2(new_n585), .A3(new_n622), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n622), .B1(new_n584), .B2(new_n585), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT41), .ZN(new_n914));
  NOR3_X1   g489(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(G299), .A2(new_n621), .ZN(new_n916));
  AOI21_X1  g491(.A(KEYINPUT41), .B1(new_n916), .B2(new_n911), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  XOR2_X1   g493(.A(new_n867), .B(new_n635), .Z(new_n919));
  NOR2_X1   g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n916), .A2(new_n911), .ZN(new_n921));
  AND2_X1   g496(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  OR3_X1    g497(.A1(new_n920), .A2(KEYINPUT42), .A3(new_n922), .ZN(new_n923));
  OAI21_X1  g498(.A(KEYINPUT42), .B1(new_n920), .B2(new_n922), .ZN(new_n924));
  XNOR2_X1  g499(.A(G303), .B(G305), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n593), .B(G290), .ZN(new_n927));
  OR2_X1    g502(.A1(new_n927), .A2(KEYINPUT111), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(KEYINPUT111), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n926), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n925), .B1(new_n927), .B2(KEYINPUT111), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n923), .A2(new_n924), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(G868), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n933), .B1(new_n923), .B2(new_n924), .ZN(new_n936));
  AND2_X1   g511(.A1(new_n866), .A2(new_n626), .ZN(new_n937));
  OAI22_X1  g512(.A1(new_n935), .A2(new_n936), .B1(KEYINPUT112), .B2(new_n937), .ZN(new_n938));
  OR2_X1    g513(.A1(new_n935), .A2(new_n936), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n938), .B1(new_n939), .B2(KEYINPUT112), .ZN(G295));
  OAI21_X1  g515(.A(new_n938), .B1(new_n939), .B2(KEYINPUT112), .ZN(G331));
  INV_X1    g516(.A(KEYINPUT43), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT116), .ZN(new_n943));
  INV_X1    g518(.A(new_n539), .ZN(new_n944));
  AOI21_X1  g519(.A(KEYINPUT73), .B1(new_n530), .B2(new_n535), .ZN(new_n945));
  OAI21_X1  g520(.A(G301), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n538), .A2(new_n539), .A3(G171), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n867), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  AND2_X1   g524(.A1(new_n946), .A2(new_n947), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(new_n867), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  AND3_X1   g527(.A1(new_n867), .A2(new_n946), .A3(new_n947), .ZN(new_n953));
  OAI21_X1  g528(.A(KEYINPUT113), .B1(new_n953), .B2(new_n948), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT113), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n951), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n912), .A2(new_n913), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n954), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  AOI22_X1  g533(.A1(new_n918), .A2(new_n952), .B1(new_n958), .B2(KEYINPUT115), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT115), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n954), .A2(new_n956), .A3(new_n960), .A4(new_n957), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n933), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n954), .A2(new_n956), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n918), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n957), .A2(new_n951), .A3(new_n949), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n964), .A2(new_n933), .A3(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(G37), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n943), .B1(new_n962), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n918), .A2(new_n952), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n958), .A2(KEYINPUT115), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n970), .A2(new_n971), .A3(new_n961), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(new_n932), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n973), .A2(KEYINPUT116), .A3(new_n967), .A4(new_n966), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n942), .B1(new_n969), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n964), .A2(new_n965), .ZN(new_n976));
  AND2_X1   g551(.A1(new_n932), .A2(KEYINPUT114), .ZN(new_n977));
  AND2_X1   g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n967), .B1(new_n976), .B2(new_n977), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n980), .A2(KEYINPUT43), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT44), .B1(new_n975), .B2(new_n981), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n973), .A2(new_n942), .A3(new_n967), .A4(new_n966), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n983), .B1(new_n980), .B2(new_n942), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT44), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n982), .A2(new_n986), .ZN(G397));
  INV_X1    g562(.A(KEYINPUT127), .ZN(new_n988));
  INV_X1    g563(.A(G1384), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n989), .B1(new_n502), .B2(new_n506), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(KEYINPUT50), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n469), .A2(new_n476), .A3(G40), .ZN(new_n992));
  INV_X1    g567(.A(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(G2090), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT50), .ZN(new_n995));
  OAI211_X1 g570(.A(new_n995), .B(new_n989), .C1(new_n502), .C2(new_n506), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n991), .A2(new_n993), .A3(new_n994), .A4(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT117), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n992), .B1(KEYINPUT50), .B2(new_n990), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n1000), .A2(KEYINPUT117), .A3(new_n994), .A4(new_n996), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT45), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n990), .A2(new_n1002), .ZN(new_n1003));
  OAI211_X1 g578(.A(KEYINPUT45), .B(new_n989), .C1(new_n502), .C2(new_n506), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1003), .A2(new_n993), .A3(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(G1971), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n999), .A2(new_n1001), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(G303), .A2(G8), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n1009), .B(KEYINPUT55), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1008), .A2(G8), .A3(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(KEYINPUT63), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n992), .B1(new_n1002), .B2(new_n990), .ZN(new_n1014));
  AOI21_X1  g589(.A(G1966), .B1(new_n1014), .B2(new_n1004), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT122), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n991), .A2(new_n993), .A3(new_n996), .ZN(new_n1017));
  OAI22_X1  g592(.A1(new_n1015), .A2(new_n1016), .B1(G2084), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1005), .A2(new_n815), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1019), .A2(KEYINPUT122), .ZN(new_n1020));
  OAI211_X1 g595(.A(G8), .B(G168), .C1(new_n1018), .C2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1013), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT123), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1008), .A2(G8), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(new_n1010), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n599), .A2(new_n600), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n515), .A2(G61), .ZN(new_n1027));
  NAND2_X1  g602(.A1(G73), .A2(G543), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n508), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g604(.A(G1981), .B1(new_n1026), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(KEYINPUT119), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT119), .ZN(new_n1032));
  NAND3_X1  g607(.A1(G305), .A2(new_n1032), .A3(G1981), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1026), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1029), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT118), .ZN(new_n1037));
  INV_X1    g612(.A(G1981), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .A4(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(KEYINPUT118), .B1(G305), .B2(G1981), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1034), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT49), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n990), .A2(new_n992), .ZN(new_n1045));
  INV_X1    g620(.A(G8), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1034), .A2(new_n1041), .A3(KEYINPUT49), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1044), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n720), .A2(G1976), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1047), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(KEYINPUT52), .ZN(new_n1052));
  INV_X1    g627(.A(G1976), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1053), .B1(new_n594), .B2(new_n596), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT52), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1054), .A2(new_n1047), .A3(new_n1055), .A4(new_n1050), .ZN(new_n1056));
  AND3_X1   g631(.A1(new_n1049), .A2(new_n1052), .A3(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1023), .B1(new_n1025), .B2(new_n1057), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1011), .B1(new_n1008), .B2(G8), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1049), .A2(new_n1052), .A3(new_n1056), .ZN(new_n1060));
  NOR3_X1   g635(.A1(new_n1059), .A2(new_n1060), .A3(KEYINPUT123), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1022), .B1(new_n1058), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT124), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n991), .A2(new_n993), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT120), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1000), .A2(KEYINPUT120), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1067), .A2(new_n1068), .A3(new_n994), .A4(new_n996), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1069), .A2(KEYINPUT121), .A3(new_n1007), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(G8), .ZN(new_n1071));
  AOI21_X1  g646(.A(KEYINPUT121), .B1(new_n1069), .B2(new_n1007), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1010), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1021), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1073), .A2(new_n1057), .A3(new_n1074), .A4(new_n1012), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT63), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  OAI211_X1 g652(.A(KEYINPUT124), .B(new_n1022), .C1(new_n1058), .C2(new_n1061), .ZN(new_n1078));
  AND3_X1   g653(.A1(new_n1064), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1049), .A2(new_n1053), .A3(new_n597), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(new_n1041), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1012), .ZN(new_n1082));
  AOI22_X1  g657(.A1(new_n1081), .A2(new_n1047), .B1(new_n1082), .B2(new_n1057), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n996), .B1(new_n1000), .B2(KEYINPUT120), .ZN(new_n1084));
  AND3_X1   g659(.A1(new_n991), .A2(KEYINPUT120), .A3(new_n993), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n848), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT57), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n582), .A2(new_n1087), .ZN(new_n1088));
  OAI211_X1 g663(.A(KEYINPUT57), .B(new_n573), .C1(new_n580), .C2(new_n581), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  XNOR2_X1  g665(.A(KEYINPUT56), .B(G2072), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1014), .A2(new_n1004), .A3(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1086), .A2(new_n1090), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(KEYINPUT61), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT60), .ZN(new_n1095));
  AOI21_X1  g670(.A(G1348), .B1(new_n1000), .B2(new_n996), .ZN(new_n1096));
  NOR3_X1   g671(.A1(new_n990), .A2(new_n992), .A3(G2067), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1095), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NOR4_X1   g673(.A1(new_n1096), .A2(new_n1095), .A3(new_n622), .A4(new_n1097), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1097), .B1(new_n1017), .B2(new_n780), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n621), .B1(new_n1100), .B2(KEYINPUT60), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1098), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(G1996), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1014), .A2(new_n1103), .A3(new_n1004), .ZN(new_n1104));
  XOR2_X1   g679(.A(KEYINPUT58), .B(G1341), .Z(new_n1105));
  OAI21_X1  g680(.A(new_n1105), .B1(new_n990), .B2(new_n992), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(KEYINPUT59), .B1(new_n1107), .B2(new_n560), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT59), .ZN(new_n1109));
  AOI211_X1 g684(.A(new_n1109), .B(new_n559), .C1(new_n1104), .C2(new_n1106), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT61), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1086), .A2(new_n1112), .A3(new_n1090), .A4(new_n1092), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1094), .A2(new_n1102), .A3(new_n1111), .A4(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1090), .B1(new_n1086), .B2(new_n1092), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1100), .A2(new_n621), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1115), .B1(new_n1093), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1114), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1057), .A2(new_n1012), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1072), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1120), .A2(G8), .A3(new_n1070), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1119), .B1(new_n1121), .B2(new_n1010), .ZN(new_n1122));
  OR2_X1    g697(.A1(new_n1005), .A2(G2078), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT53), .ZN(new_n1124));
  OR3_X1    g699(.A1(new_n1123), .A2(KEYINPUT126), .A3(new_n1124), .ZN(new_n1125));
  XOR2_X1   g700(.A(G171), .B(KEYINPUT54), .Z(new_n1126));
  NAND2_X1  g701(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1127));
  AOI22_X1  g702(.A1(new_n1123), .A2(KEYINPUT126), .B1(new_n777), .B2(new_n1017), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .A4(new_n1128), .ZN(new_n1129));
  OR2_X1    g704(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1017), .A2(new_n777), .ZN(new_n1131));
  AND3_X1   g706(.A1(new_n1130), .A2(new_n1127), .A3(new_n1131), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1129), .B1(new_n1132), .B2(new_n1126), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1118), .A2(new_n1122), .A3(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(G286), .A2(G8), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT125), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1136), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1137));
  AND3_X1   g712(.A1(new_n991), .A2(new_n993), .A3(new_n996), .ZN(new_n1138));
  INV_X1    g713(.A(G2084), .ZN(new_n1139));
  AOI22_X1  g714(.A1(new_n1019), .A2(KEYINPUT122), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1140), .A2(KEYINPUT125), .A3(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1137), .A2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1135), .B1(new_n1143), .B2(KEYINPUT51), .ZN(new_n1144));
  NOR3_X1   g719(.A1(new_n1018), .A2(new_n1020), .A3(new_n1136), .ZN(new_n1145));
  AOI21_X1  g720(.A(KEYINPUT125), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1146));
  OAI21_X1  g721(.A(G168), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT51), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1148), .A2(new_n1046), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g725(.A(G8), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(new_n1148), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1144), .B1(new_n1150), .B2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1083), .B1(new_n1134), .B2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n988), .B1(new_n1079), .B2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(G286), .B1(new_n1137), .B2(new_n1142), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1149), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1152), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1148), .B1(new_n1137), .B2(new_n1142), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1158), .B1(new_n1159), .B2(new_n1135), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1160), .A2(new_n1122), .A3(new_n1118), .A4(new_n1133), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1064), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1161), .A2(new_n1162), .A3(KEYINPUT127), .A4(new_n1083), .ZN(new_n1163));
  OR2_X1    g738(.A1(new_n1160), .A2(KEYINPUT62), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1160), .A2(KEYINPUT62), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1125), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1166));
  AND3_X1   g741(.A1(new_n1122), .A2(G171), .A3(new_n1166), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1164), .A2(new_n1165), .A3(new_n1167), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1155), .A2(new_n1163), .A3(new_n1168), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1003), .A2(new_n992), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n766), .A2(new_n1103), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n764), .A2(G1996), .ZN(new_n1172));
  INV_X1    g747(.A(G2067), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n836), .A2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n835), .A2(G2067), .ZN(new_n1175));
  AND2_X1   g750(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1171), .A2(new_n1172), .A3(new_n1176), .ZN(new_n1177));
  XOR2_X1   g752(.A(new_n742), .B(new_n744), .Z(new_n1178));
  OR2_X1    g753(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  XNOR2_X1  g754(.A(G290), .B(G1986), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1170), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1169), .A2(new_n1181), .ZN(new_n1182));
  NOR2_X1   g757(.A1(G290), .A2(G1986), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1170), .A2(new_n1183), .ZN(new_n1184));
  XOR2_X1   g759(.A(new_n1184), .B(KEYINPUT48), .Z(new_n1185));
  AOI21_X1  g760(.A(new_n1185), .B1(new_n1179), .B2(new_n1170), .ZN(new_n1186));
  INV_X1    g761(.A(new_n1176), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1170), .B1(new_n1187), .B2(new_n764), .ZN(new_n1188));
  NOR3_X1   g763(.A1(new_n1003), .A2(G1996), .A3(new_n992), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1189), .A2(KEYINPUT46), .ZN(new_n1190));
  OR2_X1    g765(.A1(new_n1189), .A2(KEYINPUT46), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1188), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  XOR2_X1   g767(.A(new_n1192), .B(KEYINPUT47), .Z(new_n1193));
  NAND3_X1  g768(.A1(new_n740), .A2(new_n744), .A3(new_n741), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1174), .B1(new_n1177), .B2(new_n1194), .ZN(new_n1195));
  AOI211_X1 g770(.A(new_n1186), .B(new_n1193), .C1(new_n1170), .C2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1182), .A2(new_n1196), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g772(.A(G319), .ZN(new_n1199));
  NOR2_X1   g773(.A1(G227), .A2(new_n1199), .ZN(new_n1200));
  AND4_X1   g774(.A1(new_n670), .A2(new_n707), .A3(new_n708), .A4(new_n1200), .ZN(new_n1201));
  NAND3_X1  g775(.A1(new_n906), .A2(new_n984), .A3(new_n1201), .ZN(G225));
  INV_X1    g776(.A(G225), .ZN(G308));
endmodule


