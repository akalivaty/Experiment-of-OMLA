

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596;

  XNOR2_X1 U326 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U327 ( .A(n442), .B(KEYINPUT118), .ZN(n443) );
  AND2_X1 U328 ( .A1(G232GAT), .A2(G233GAT), .ZN(n294) );
  XOR2_X1 U329 ( .A(n373), .B(KEYINPUT73), .Z(n295) );
  INV_X1 U330 ( .A(KEYINPUT111), .ZN(n385) );
  XNOR2_X1 U331 ( .A(n416), .B(n294), .ZN(n356) );
  XNOR2_X1 U332 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U333 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U334 ( .A(n383), .B(n382), .ZN(n388) );
  XOR2_X1 U335 ( .A(KEYINPUT36), .B(n565), .Z(n594) );
  XOR2_X1 U336 ( .A(n361), .B(n360), .Z(n565) );
  XOR2_X1 U337 ( .A(n351), .B(n329), .Z(n580) );
  XNOR2_X1 U338 ( .A(n468), .B(G190GAT), .ZN(n469) );
  XNOR2_X1 U339 ( .A(n470), .B(n469), .ZN(G1351GAT) );
  XOR2_X1 U340 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n297) );
  XNOR2_X1 U341 ( .A(KEYINPUT84), .B(G183GAT), .ZN(n296) );
  XNOR2_X1 U342 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U343 ( .A(KEYINPUT17), .B(n298), .Z(n448) );
  XOR2_X1 U344 ( .A(G211GAT), .B(KEYINPUT21), .Z(n300) );
  XNOR2_X1 U345 ( .A(G197GAT), .B(G218GAT), .ZN(n299) );
  XNOR2_X1 U346 ( .A(n300), .B(n299), .ZN(n431) );
  XNOR2_X1 U347 ( .A(G36GAT), .B(G190GAT), .ZN(n301) );
  XNOR2_X1 U348 ( .A(n301), .B(KEYINPUT77), .ZN(n355) );
  XNOR2_X1 U349 ( .A(n431), .B(n355), .ZN(n311) );
  INV_X1 U350 ( .A(G92GAT), .ZN(n302) );
  NAND2_X1 U351 ( .A1(G64GAT), .A2(n302), .ZN(n305) );
  INV_X1 U352 ( .A(G64GAT), .ZN(n303) );
  NAND2_X1 U353 ( .A1(n303), .A2(G92GAT), .ZN(n304) );
  NAND2_X1 U354 ( .A1(n305), .A2(n304), .ZN(n307) );
  XNOR2_X1 U355 ( .A(G176GAT), .B(G204GAT), .ZN(n306) );
  XNOR2_X1 U356 ( .A(n307), .B(n306), .ZN(n367) );
  XOR2_X1 U357 ( .A(G169GAT), .B(G8GAT), .Z(n317) );
  XOR2_X1 U358 ( .A(n367), .B(n317), .Z(n309) );
  NAND2_X1 U359 ( .A1(G226GAT), .A2(G233GAT), .ZN(n308) );
  XNOR2_X1 U360 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U361 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U362 ( .A(n448), .B(n312), .Z(n531) );
  INV_X1 U363 ( .A(n531), .ZN(n506) );
  XNOR2_X1 U364 ( .A(G43GAT), .B(KEYINPUT7), .ZN(n313) );
  XNOR2_X1 U365 ( .A(n313), .B(G29GAT), .ZN(n314) );
  XOR2_X1 U366 ( .A(n314), .B(KEYINPUT68), .Z(n316) );
  XNOR2_X1 U367 ( .A(KEYINPUT8), .B(KEYINPUT69), .ZN(n315) );
  XNOR2_X1 U368 ( .A(n316), .B(n315), .ZN(n351) );
  XOR2_X1 U369 ( .A(G113GAT), .B(G1GAT), .Z(n402) );
  XOR2_X1 U370 ( .A(n317), .B(n402), .Z(n319) );
  NAND2_X1 U371 ( .A1(G229GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U372 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U373 ( .A(G141GAT), .B(G22GAT), .Z(n437) );
  XOR2_X1 U374 ( .A(n320), .B(n437), .Z(n328) );
  XOR2_X1 U375 ( .A(G197GAT), .B(G15GAT), .Z(n322) );
  XNOR2_X1 U376 ( .A(G36GAT), .B(G50GAT), .ZN(n321) );
  XNOR2_X1 U377 ( .A(n322), .B(n321), .ZN(n326) );
  XOR2_X1 U378 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n324) );
  XNOR2_X1 U379 ( .A(KEYINPUT70), .B(KEYINPUT67), .ZN(n323) );
  XNOR2_X1 U380 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U381 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U382 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U383 ( .A(G155GAT), .B(G211GAT), .Z(n331) );
  XNOR2_X1 U384 ( .A(G183GAT), .B(G71GAT), .ZN(n330) );
  XNOR2_X1 U385 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U386 ( .A(G57GAT), .B(KEYINPUT13), .Z(n379) );
  XOR2_X1 U387 ( .A(n332), .B(n379), .Z(n334) );
  XNOR2_X1 U388 ( .A(G22GAT), .B(G78GAT), .ZN(n333) );
  XNOR2_X1 U389 ( .A(n334), .B(n333), .ZN(n347) );
  XOR2_X1 U390 ( .A(KEYINPUT81), .B(KEYINPUT80), .Z(n336) );
  NAND2_X1 U391 ( .A1(G231GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U392 ( .A(n336), .B(n335), .ZN(n340) );
  XOR2_X1 U393 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n338) );
  XNOR2_X1 U394 ( .A(KEYINPUT15), .B(KEYINPUT78), .ZN(n337) );
  XNOR2_X1 U395 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U396 ( .A(n340), .B(n339), .Z(n345) );
  XOR2_X1 U397 ( .A(G15GAT), .B(G127GAT), .Z(n450) );
  XOR2_X1 U398 ( .A(KEYINPUT79), .B(G64GAT), .Z(n342) );
  XNOR2_X1 U399 ( .A(G8GAT), .B(G1GAT), .ZN(n341) );
  XNOR2_X1 U400 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U401 ( .A(n450), .B(n343), .ZN(n344) );
  XNOR2_X1 U402 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U403 ( .A(n347), .B(n346), .Z(n588) );
  INV_X1 U404 ( .A(n588), .ZN(n574) );
  XOR2_X1 U405 ( .A(KEYINPUT66), .B(KEYINPUT9), .Z(n349) );
  XNOR2_X1 U406 ( .A(G106GAT), .B(G92GAT), .ZN(n348) );
  XNOR2_X1 U407 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U408 ( .A(n351), .B(n350), .ZN(n361) );
  XOR2_X1 U409 ( .A(KEYINPUT75), .B(KEYINPUT10), .Z(n353) );
  XOR2_X1 U410 ( .A(G50GAT), .B(G162GAT), .Z(n436) );
  XOR2_X1 U411 ( .A(G99GAT), .B(G85GAT), .Z(n366) );
  XNOR2_X1 U412 ( .A(n436), .B(n366), .ZN(n352) );
  XNOR2_X1 U413 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U414 ( .A(n354), .B(KEYINPUT11), .Z(n359) );
  XOR2_X1 U415 ( .A(G134GAT), .B(KEYINPUT76), .Z(n416) );
  XNOR2_X1 U416 ( .A(G218GAT), .B(n357), .ZN(n358) );
  XNOR2_X1 U417 ( .A(n359), .B(n358), .ZN(n360) );
  NOR2_X1 U418 ( .A1(n574), .A2(n594), .ZN(n364) );
  XOR2_X1 U419 ( .A(KEYINPUT45), .B(KEYINPUT110), .Z(n362) );
  XNOR2_X1 U420 ( .A(KEYINPUT65), .B(n362), .ZN(n363) );
  XNOR2_X1 U421 ( .A(n364), .B(n363), .ZN(n384) );
  INV_X1 U422 ( .A(n367), .ZN(n365) );
  NAND2_X1 U423 ( .A1(n365), .A2(n366), .ZN(n370) );
  INV_X1 U424 ( .A(n366), .ZN(n368) );
  NAND2_X1 U425 ( .A1(n368), .A2(n367), .ZN(n369) );
  NAND2_X1 U426 ( .A1(n370), .A2(n369), .ZN(n372) );
  NAND2_X1 U427 ( .A1(G230GAT), .A2(G233GAT), .ZN(n371) );
  XNOR2_X1 U428 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U429 ( .A(G78GAT), .B(G148GAT), .Z(n375) );
  XNOR2_X1 U430 ( .A(G106GAT), .B(KEYINPUT71), .ZN(n374) );
  XNOR2_X1 U431 ( .A(n375), .B(n374), .ZN(n434) );
  XNOR2_X1 U432 ( .A(n434), .B(KEYINPUT72), .ZN(n376) );
  XNOR2_X1 U433 ( .A(n295), .B(n376), .ZN(n383) );
  XOR2_X1 U434 ( .A(KEYINPUT74), .B(KEYINPUT32), .Z(n378) );
  XNOR2_X1 U435 ( .A(KEYINPUT31), .B(KEYINPUT33), .ZN(n377) );
  XOR2_X1 U436 ( .A(n378), .B(n377), .Z(n381) );
  XOR2_X1 U437 ( .A(G120GAT), .B(G71GAT), .Z(n453) );
  XNOR2_X1 U438 ( .A(n453), .B(n379), .ZN(n380) );
  NAND2_X1 U439 ( .A1(n384), .A2(n388), .ZN(n386) );
  NOR2_X1 U440 ( .A1(n580), .A2(n387), .ZN(n396) );
  XNOR2_X1 U441 ( .A(n388), .B(KEYINPUT41), .ZN(n560) );
  NAND2_X1 U442 ( .A1(n560), .A2(n580), .ZN(n390) );
  XOR2_X1 U443 ( .A(KEYINPUT108), .B(KEYINPUT46), .Z(n389) );
  XNOR2_X1 U444 ( .A(n390), .B(n389), .ZN(n391) );
  NOR2_X1 U445 ( .A1(n588), .A2(n391), .ZN(n392) );
  XNOR2_X1 U446 ( .A(n392), .B(KEYINPUT109), .ZN(n393) );
  NOR2_X1 U447 ( .A1(n393), .A2(n565), .ZN(n394) );
  XOR2_X1 U448 ( .A(KEYINPUT47), .B(n394), .Z(n395) );
  NOR2_X1 U449 ( .A1(n396), .A2(n395), .ZN(n397) );
  XNOR2_X1 U450 ( .A(n397), .B(KEYINPUT48), .ZN(n540) );
  NOR2_X1 U451 ( .A1(n506), .A2(n540), .ZN(n398) );
  XNOR2_X1 U452 ( .A(n398), .B(KEYINPUT54), .ZN(n423) );
  XOR2_X1 U453 ( .A(G85GAT), .B(G148GAT), .Z(n400) );
  XNOR2_X1 U454 ( .A(G120GAT), .B(G127GAT), .ZN(n399) );
  XNOR2_X1 U455 ( .A(n400), .B(n399), .ZN(n401) );
  XOR2_X1 U456 ( .A(n401), .B(G162GAT), .Z(n404) );
  XNOR2_X1 U457 ( .A(G29GAT), .B(n402), .ZN(n403) );
  XNOR2_X1 U458 ( .A(n404), .B(n403), .ZN(n422) );
  XOR2_X1 U459 ( .A(KEYINPUT90), .B(KEYINPUT1), .Z(n406) );
  XNOR2_X1 U460 ( .A(G141GAT), .B(G57GAT), .ZN(n405) );
  XNOR2_X1 U461 ( .A(n406), .B(n405), .ZN(n410) );
  XOR2_X1 U462 ( .A(KEYINPUT6), .B(KEYINPUT92), .Z(n408) );
  XNOR2_X1 U463 ( .A(KEYINPUT4), .B(KEYINPUT91), .ZN(n407) );
  XNOR2_X1 U464 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U465 ( .A(n410), .B(n409), .Z(n415) );
  XOR2_X1 U466 ( .A(KEYINPUT5), .B(KEYINPUT89), .Z(n412) );
  NAND2_X1 U467 ( .A1(G225GAT), .A2(G233GAT), .ZN(n411) );
  XNOR2_X1 U468 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U469 ( .A(KEYINPUT93), .B(n413), .ZN(n414) );
  XNOR2_X1 U470 ( .A(n415), .B(n414), .ZN(n417) );
  XOR2_X1 U471 ( .A(n417), .B(n416), .Z(n420) );
  XOR2_X1 U472 ( .A(KEYINPUT0), .B(KEYINPUT83), .Z(n449) );
  XNOR2_X1 U473 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n418) );
  XNOR2_X1 U474 ( .A(n418), .B(KEYINPUT2), .ZN(n430) );
  XNOR2_X1 U475 ( .A(n449), .B(n430), .ZN(n419) );
  XNOR2_X1 U476 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U477 ( .A(n422), .B(n421), .ZN(n528) );
  INV_X1 U478 ( .A(n528), .ZN(n503) );
  NAND2_X1 U479 ( .A1(n423), .A2(n503), .ZN(n424) );
  XNOR2_X1 U480 ( .A(n424), .B(KEYINPUT64), .ZN(n578) );
  XOR2_X1 U481 ( .A(G204GAT), .B(KEYINPUT22), .Z(n426) );
  XNOR2_X1 U482 ( .A(KEYINPUT23), .B(KEYINPUT88), .ZN(n425) );
  XNOR2_X1 U483 ( .A(n426), .B(n425), .ZN(n441) );
  XOR2_X1 U484 ( .A(KEYINPUT87), .B(KEYINPUT24), .Z(n428) );
  NAND2_X1 U485 ( .A1(G228GAT), .A2(G233GAT), .ZN(n427) );
  XNOR2_X1 U486 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U487 ( .A(n429), .B(KEYINPUT86), .Z(n433) );
  XNOR2_X1 U488 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U489 ( .A(n433), .B(n432), .ZN(n435) );
  XOR2_X1 U490 ( .A(n435), .B(n434), .Z(n439) );
  XNOR2_X1 U491 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U492 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U493 ( .A(n441), .B(n440), .ZN(n483) );
  NOR2_X1 U494 ( .A1(n578), .A2(n483), .ZN(n444) );
  INV_X1 U495 ( .A(KEYINPUT55), .ZN(n442) );
  XNOR2_X1 U496 ( .A(n444), .B(n443), .ZN(n462) );
  XOR2_X1 U497 ( .A(G99GAT), .B(G113GAT), .Z(n446) );
  XNOR2_X1 U498 ( .A(G169GAT), .B(G43GAT), .ZN(n445) );
  XNOR2_X1 U499 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U500 ( .A(n448), .B(n447), .ZN(n461) );
  XOR2_X1 U501 ( .A(G190GAT), .B(G134GAT), .Z(n452) );
  XNOR2_X1 U502 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U503 ( .A(n452), .B(n451), .ZN(n454) );
  XOR2_X1 U504 ( .A(n454), .B(n453), .Z(n459) );
  XOR2_X1 U505 ( .A(G176GAT), .B(KEYINPUT85), .Z(n456) );
  NAND2_X1 U506 ( .A1(G227GAT), .A2(G233GAT), .ZN(n455) );
  XNOR2_X1 U507 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U508 ( .A(KEYINPUT20), .B(n457), .ZN(n458) );
  XNOR2_X1 U509 ( .A(n459), .B(n458), .ZN(n460) );
  XOR2_X1 U510 ( .A(n461), .B(n460), .Z(n509) );
  INV_X1 U511 ( .A(n509), .ZN(n542) );
  NAND2_X1 U512 ( .A1(n462), .A2(n542), .ZN(n573) );
  XNOR2_X1 U513 ( .A(KEYINPUT102), .B(n560), .ZN(n545) );
  INV_X1 U514 ( .A(n545), .ZN(n463) );
  NOR2_X1 U515 ( .A1(n573), .A2(n463), .ZN(n467) );
  XNOR2_X1 U516 ( .A(KEYINPUT57), .B(KEYINPUT120), .ZN(n465) );
  XNOR2_X1 U517 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n464) );
  XNOR2_X1 U518 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U519 ( .A(n467), .B(n466), .ZN(G1349GAT) );
  INV_X1 U520 ( .A(n565), .ZN(n471) );
  NOR2_X1 U521 ( .A1(n471), .A2(n573), .ZN(n470) );
  XNOR2_X1 U522 ( .A(KEYINPUT121), .B(KEYINPUT58), .ZN(n468) );
  XOR2_X1 U523 ( .A(KEYINPUT98), .B(KEYINPUT34), .Z(n490) );
  NAND2_X1 U524 ( .A1(n580), .A2(n388), .ZN(n501) );
  XOR2_X1 U525 ( .A(KEYINPUT82), .B(KEYINPUT16), .Z(n473) );
  NAND2_X1 U526 ( .A1(n588), .A2(n471), .ZN(n472) );
  XNOR2_X1 U527 ( .A(n473), .B(n472), .ZN(n488) );
  XOR2_X1 U528 ( .A(KEYINPUT25), .B(KEYINPUT96), .Z(n477) );
  NOR2_X1 U529 ( .A1(n509), .A2(n506), .ZN(n474) );
  NOR2_X1 U530 ( .A1(n483), .A2(n474), .ZN(n475) );
  XNOR2_X1 U531 ( .A(n475), .B(KEYINPUT95), .ZN(n476) );
  XNOR2_X1 U532 ( .A(n477), .B(n476), .ZN(n481) );
  NAND2_X1 U533 ( .A1(n483), .A2(n509), .ZN(n478) );
  XNOR2_X1 U534 ( .A(n478), .B(KEYINPUT26), .ZN(n579) );
  XOR2_X1 U535 ( .A(KEYINPUT27), .B(n531), .Z(n484) );
  NOR2_X1 U536 ( .A1(n579), .A2(n484), .ZN(n479) );
  XOR2_X1 U537 ( .A(KEYINPUT94), .B(n479), .Z(n480) );
  NAND2_X1 U538 ( .A1(n481), .A2(n480), .ZN(n482) );
  NAND2_X1 U539 ( .A1(n503), .A2(n482), .ZN(n486) );
  XOR2_X1 U540 ( .A(KEYINPUT28), .B(n483), .Z(n512) );
  INV_X1 U541 ( .A(n512), .ZN(n536) );
  OR2_X1 U542 ( .A1(n503), .A2(n484), .ZN(n556) );
  NOR2_X1 U543 ( .A1(n536), .A2(n556), .ZN(n541) );
  NAND2_X1 U544 ( .A1(n541), .A2(n509), .ZN(n485) );
  NAND2_X1 U545 ( .A1(n486), .A2(n485), .ZN(n487) );
  XOR2_X1 U546 ( .A(KEYINPUT97), .B(n487), .Z(n498) );
  NAND2_X1 U547 ( .A1(n488), .A2(n498), .ZN(n516) );
  NOR2_X1 U548 ( .A1(n501), .A2(n516), .ZN(n496) );
  NAND2_X1 U549 ( .A1(n496), .A2(n528), .ZN(n489) );
  XNOR2_X1 U550 ( .A(n490), .B(n489), .ZN(n491) );
  XOR2_X1 U551 ( .A(G1GAT), .B(n491), .Z(G1324GAT) );
  XOR2_X1 U552 ( .A(G8GAT), .B(KEYINPUT99), .Z(n493) );
  NAND2_X1 U553 ( .A1(n496), .A2(n531), .ZN(n492) );
  XNOR2_X1 U554 ( .A(n493), .B(n492), .ZN(G1325GAT) );
  XOR2_X1 U555 ( .A(G15GAT), .B(KEYINPUT35), .Z(n495) );
  NAND2_X1 U556 ( .A1(n496), .A2(n542), .ZN(n494) );
  XNOR2_X1 U557 ( .A(n495), .B(n494), .ZN(G1326GAT) );
  NAND2_X1 U558 ( .A1(n496), .A2(n536), .ZN(n497) );
  XNOR2_X1 U559 ( .A(n497), .B(G22GAT), .ZN(G1327GAT) );
  XNOR2_X1 U560 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n505) );
  NAND2_X1 U561 ( .A1(n574), .A2(n498), .ZN(n499) );
  NOR2_X1 U562 ( .A1(n499), .A2(n594), .ZN(n500) );
  XNOR2_X1 U563 ( .A(n500), .B(KEYINPUT37), .ZN(n527) );
  NOR2_X1 U564 ( .A1(n527), .A2(n501), .ZN(n502) );
  XOR2_X1 U565 ( .A(KEYINPUT38), .B(n502), .Z(n513) );
  NOR2_X1 U566 ( .A1(n503), .A2(n513), .ZN(n504) );
  XNOR2_X1 U567 ( .A(n505), .B(n504), .ZN(G1328GAT) );
  NOR2_X1 U568 ( .A1(n513), .A2(n506), .ZN(n507) );
  XOR2_X1 U569 ( .A(KEYINPUT100), .B(n507), .Z(n508) );
  XNOR2_X1 U570 ( .A(G36GAT), .B(n508), .ZN(G1329GAT) );
  NOR2_X1 U571 ( .A1(n513), .A2(n509), .ZN(n510) );
  XOR2_X1 U572 ( .A(KEYINPUT40), .B(n510), .Z(n511) );
  XNOR2_X1 U573 ( .A(G43GAT), .B(n511), .ZN(G1330GAT) );
  NOR2_X1 U574 ( .A1(n513), .A2(n512), .ZN(n515) );
  XNOR2_X1 U575 ( .A(G50GAT), .B(KEYINPUT101), .ZN(n514) );
  XNOR2_X1 U576 ( .A(n515), .B(n514), .ZN(G1331GAT) );
  XNOR2_X1 U577 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n518) );
  INV_X1 U578 ( .A(n580), .ZN(n570) );
  NAND2_X1 U579 ( .A1(n545), .A2(n570), .ZN(n526) );
  NOR2_X1 U580 ( .A1(n526), .A2(n516), .ZN(n522) );
  NAND2_X1 U581 ( .A1(n522), .A2(n528), .ZN(n517) );
  XNOR2_X1 U582 ( .A(n518), .B(n517), .ZN(G1332GAT) );
  XOR2_X1 U583 ( .A(G64GAT), .B(KEYINPUT103), .Z(n520) );
  NAND2_X1 U584 ( .A1(n522), .A2(n531), .ZN(n519) );
  XNOR2_X1 U585 ( .A(n520), .B(n519), .ZN(G1333GAT) );
  NAND2_X1 U586 ( .A1(n522), .A2(n542), .ZN(n521) );
  XNOR2_X1 U587 ( .A(n521), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U588 ( .A(KEYINPUT104), .B(KEYINPUT43), .Z(n524) );
  NAND2_X1 U589 ( .A1(n522), .A2(n536), .ZN(n523) );
  XNOR2_X1 U590 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U591 ( .A(G78GAT), .B(n525), .ZN(G1335GAT) );
  XOR2_X1 U592 ( .A(G85GAT), .B(KEYINPUT105), .Z(n530) );
  NOR2_X1 U593 ( .A1(n527), .A2(n526), .ZN(n537) );
  NAND2_X1 U594 ( .A1(n537), .A2(n528), .ZN(n529) );
  XNOR2_X1 U595 ( .A(n530), .B(n529), .ZN(G1336GAT) );
  XNOR2_X1 U596 ( .A(G92GAT), .B(KEYINPUT106), .ZN(n533) );
  NAND2_X1 U597 ( .A1(n531), .A2(n537), .ZN(n532) );
  XNOR2_X1 U598 ( .A(n533), .B(n532), .ZN(G1337GAT) );
  XOR2_X1 U599 ( .A(G99GAT), .B(KEYINPUT107), .Z(n535) );
  NAND2_X1 U600 ( .A1(n537), .A2(n542), .ZN(n534) );
  XNOR2_X1 U601 ( .A(n535), .B(n534), .ZN(G1338GAT) );
  NAND2_X1 U602 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U603 ( .A(n538), .B(KEYINPUT44), .ZN(n539) );
  XNOR2_X1 U604 ( .A(G106GAT), .B(n539), .ZN(G1339GAT) );
  NAND2_X1 U605 ( .A1(n542), .A2(n541), .ZN(n543) );
  NOR2_X1 U606 ( .A1(n540), .A2(n543), .ZN(n553) );
  NAND2_X1 U607 ( .A1(n553), .A2(n580), .ZN(n544) );
  XNOR2_X1 U608 ( .A(n544), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT113), .B(KEYINPUT49), .Z(n547) );
  NAND2_X1 U610 ( .A1(n553), .A2(n545), .ZN(n546) );
  XNOR2_X1 U611 ( .A(n547), .B(n546), .ZN(n549) );
  XOR2_X1 U612 ( .A(G120GAT), .B(KEYINPUT112), .Z(n548) );
  XNOR2_X1 U613 ( .A(n549), .B(n548), .ZN(G1341GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT50), .B(KEYINPUT114), .Z(n551) );
  NAND2_X1 U615 ( .A1(n553), .A2(n588), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n551), .B(n550), .ZN(n552) );
  XOR2_X1 U617 ( .A(G127GAT), .B(n552), .Z(G1342GAT) );
  XOR2_X1 U618 ( .A(G134GAT), .B(KEYINPUT51), .Z(n555) );
  NAND2_X1 U619 ( .A1(n553), .A2(n565), .ZN(n554) );
  XNOR2_X1 U620 ( .A(n555), .B(n554), .ZN(G1343GAT) );
  OR2_X1 U621 ( .A1(n579), .A2(n556), .ZN(n557) );
  NOR2_X1 U622 ( .A1(n540), .A2(n557), .ZN(n566) );
  AND2_X1 U623 ( .A1(n580), .A2(n566), .ZN(n559) );
  XNOR2_X1 U624 ( .A(G141GAT), .B(KEYINPUT115), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n559), .B(n558), .ZN(G1344GAT) );
  XOR2_X1 U626 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n562) );
  NAND2_X1 U627 ( .A1(n566), .A2(n560), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U629 ( .A(G148GAT), .B(n563), .ZN(G1345GAT) );
  NAND2_X1 U630 ( .A1(n566), .A2(n588), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n564), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U632 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n568) );
  NAND2_X1 U633 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U635 ( .A(G162GAT), .B(n569), .ZN(G1347GAT) );
  NOR2_X1 U636 ( .A1(n570), .A2(n573), .ZN(n572) );
  XNOR2_X1 U637 ( .A(G169GAT), .B(KEYINPUT119), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(G1348GAT) );
  NOR2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U640 ( .A(G183GAT), .B(n575), .Z(G1350GAT) );
  XOR2_X1 U641 ( .A(KEYINPUT60), .B(KEYINPUT123), .Z(n577) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(KEYINPUT122), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(n583) );
  NOR2_X1 U644 ( .A1(n578), .A2(n579), .ZN(n589) );
  NAND2_X1 U645 ( .A1(n589), .A2(n580), .ZN(n581) );
  XOR2_X1 U646 ( .A(KEYINPUT59), .B(n581), .Z(n582) );
  XNOR2_X1 U647 ( .A(n583), .B(n582), .ZN(G1352GAT) );
  INV_X1 U648 ( .A(n589), .ZN(n593) );
  NOR2_X1 U649 ( .A1(n593), .A2(n388), .ZN(n587) );
  XOR2_X1 U650 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n585) );
  XNOR2_X1 U651 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n584) );
  XNOR2_X1 U652 ( .A(n585), .B(n584), .ZN(n586) );
  XNOR2_X1 U653 ( .A(n587), .B(n586), .ZN(G1353GAT) );
  NAND2_X1 U654 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U655 ( .A(n590), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U656 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n592) );
  XNOR2_X1 U657 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n591) );
  XNOR2_X1 U658 ( .A(n592), .B(n591), .ZN(n596) );
  NOR2_X1 U659 ( .A1(n594), .A2(n593), .ZN(n595) );
  XOR2_X1 U660 ( .A(n596), .B(n595), .Z(G1355GAT) );
endmodule

