//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 0 1 1 1 1 1 1 0 0 0 0 1 1 0 0 1 0 1 0 1 0 0 1 0 0 0 0 1 0 0 0 1 1 0 0 1 0 0 1 0 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:38 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1299,
    new_n1300;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT0), .Z(new_n209));
  AOI22_X1  g0009(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n210));
  INV_X1    g0010(.A(G87), .ZN(new_n211));
  INV_X1    g0011(.A(G250), .ZN(new_n212));
  OAI21_X1  g0012(.A(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  AOI21_X1  g0013(.A(new_n213), .B1(G116), .B2(G270), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G58), .A2(G232), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G107), .A2(G264), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G50), .A2(G226), .ZN(new_n217));
  NAND4_X1  g0017(.A1(new_n214), .A2(new_n215), .A3(new_n216), .A4(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(G68), .ZN(new_n219));
  INV_X1    g0019(.A(G238), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n206), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT1), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  INV_X1    g0024(.A(G20), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g0026(.A(new_n201), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(G50), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  AOI211_X1 g0029(.A(new_n209), .B(new_n223), .C1(new_n226), .C2(new_n229), .ZN(G361));
  XOR2_X1   g0030(.A(KEYINPUT64), .B(KEYINPUT2), .Z(new_n231));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G226), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G250), .B(G257), .Z(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n235), .B(new_n238), .Z(G358));
  XOR2_X1   g0039(.A(G68), .B(G77), .Z(new_n240));
  XOR2_X1   g0040(.A(G50), .B(G58), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G351));
  NOR2_X1   g0046(.A1(G41), .A2(G45), .ZN(new_n247));
  INV_X1    g0047(.A(KEYINPUT65), .ZN(new_n248));
  INV_X1    g0048(.A(G274), .ZN(new_n249));
  NOR4_X1   g0049(.A1(new_n247), .A2(new_n248), .A3(new_n249), .A4(G1), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n249), .A2(G1), .ZN(new_n251));
  INV_X1    g0051(.A(G41), .ZN(new_n252));
  INV_X1    g0052(.A(G45), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  AOI21_X1  g0054(.A(KEYINPUT65), .B1(new_n251), .B2(new_n254), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n250), .A2(new_n255), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n224), .B1(G33), .B2(G41), .ZN(new_n257));
  AND2_X1   g0057(.A1(KEYINPUT66), .A2(G1), .ZN(new_n258));
  NOR2_X1   g0058(.A1(KEYINPUT66), .A2(G1), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n254), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT67), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  OAI211_X1 g0062(.A(new_n254), .B(KEYINPUT67), .C1(new_n258), .C2(new_n259), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n257), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n256), .B1(new_n264), .B2(G226), .ZN(new_n265));
  INV_X1    g0065(.A(G33), .ZN(new_n266));
  OAI211_X1 g0066(.A(G1), .B(G13), .C1(new_n266), .C2(new_n252), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT3), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(new_n266), .ZN(new_n269));
  NAND2_X1  g0069(.A1(KEYINPUT3), .A2(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NOR2_X1   g0071(.A1(G222), .A2(G1698), .ZN(new_n272));
  INV_X1    g0072(.A(G1698), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n273), .A2(G223), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n271), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n275), .B1(G77), .B2(new_n271), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n265), .B1(new_n267), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G200), .ZN(new_n278));
  INV_X1    g0078(.A(G190), .ZN(new_n279));
  OR2_X1    g0079(.A1(KEYINPUT68), .A2(G58), .ZN(new_n280));
  NAND2_X1  g0080(.A1(KEYINPUT68), .A2(G58), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n280), .A2(KEYINPUT8), .A3(new_n281), .ZN(new_n282));
  OR2_X1    g0082(.A1(KEYINPUT8), .A2(G58), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n266), .A2(G20), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G150), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n225), .A2(new_n266), .ZN(new_n288));
  OAI22_X1  g0088(.A1(new_n284), .A2(new_n286), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n289), .B1(G20), .B2(new_n203), .ZN(new_n290));
  NAND3_X1  g0090(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(new_n224), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  OAI211_X1 g0093(.A(G13), .B(G20), .C1(new_n258), .C2(new_n259), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n202), .ZN(new_n295));
  XNOR2_X1  g0095(.A(KEYINPUT66), .B(G1), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n292), .B1(new_n296), .B2(G20), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n295), .B1(new_n297), .B2(new_n202), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT69), .ZN(new_n299));
  AND2_X1   g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n298), .A2(new_n299), .ZN(new_n301));
  OAI22_X1  g0101(.A1(new_n290), .A2(new_n293), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  AND2_X1   g0102(.A1(new_n302), .A2(KEYINPUT9), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n302), .A2(KEYINPUT9), .ZN(new_n304));
  OAI221_X1 g0104(.A(new_n278), .B1(new_n279), .B2(new_n277), .C1(new_n303), .C2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT10), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT73), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n306), .B1(new_n278), .B2(new_n307), .ZN(new_n308));
  XNOR2_X1  g0108(.A(new_n305), .B(new_n308), .ZN(new_n309));
  XOR2_X1   g0109(.A(KEYINPUT70), .B(G179), .Z(new_n310));
  OR2_X1    g0110(.A1(new_n277), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G169), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n277), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n311), .A2(new_n302), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n309), .A2(new_n314), .ZN(new_n315));
  XOR2_X1   g0115(.A(KEYINPUT8), .B(G58), .Z(new_n316));
  NOR2_X1   g0116(.A1(G20), .A2(G33), .ZN(new_n317));
  AOI22_X1  g0117(.A1(new_n316), .A2(new_n317), .B1(G20), .B2(G77), .ZN(new_n318));
  XNOR2_X1  g0118(.A(KEYINPUT15), .B(G87), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(KEYINPUT71), .ZN(new_n320));
  OR2_X1    g0120(.A1(KEYINPUT15), .A2(G87), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT71), .ZN(new_n322));
  NAND2_X1  g0122(.A1(KEYINPUT15), .A2(G87), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n321), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n320), .A2(new_n324), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n318), .B1(new_n325), .B2(new_n286), .ZN(new_n326));
  INV_X1    g0126(.A(G77), .ZN(new_n327));
  INV_X1    g0127(.A(new_n294), .ZN(new_n328));
  AOI22_X1  g0128(.A1(new_n326), .A2(new_n292), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n297), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n329), .B1(new_n327), .B2(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n271), .A2(G232), .A3(new_n273), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n271), .A2(G238), .A3(G1698), .ZN(new_n333));
  INV_X1    g0133(.A(G107), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n332), .B(new_n333), .C1(new_n334), .C2(new_n271), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n256), .B1(new_n335), .B2(new_n257), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n264), .A2(G244), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n331), .B1(G200), .B2(new_n338), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n339), .B1(new_n279), .B2(new_n338), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n338), .A2(new_n312), .ZN(new_n341));
  INV_X1    g0141(.A(new_n310), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n336), .A2(new_n342), .A3(new_n337), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n341), .A2(new_n331), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n340), .A2(new_n344), .ZN(new_n345));
  XNOR2_X1  g0145(.A(new_n345), .B(KEYINPUT72), .ZN(new_n346));
  INV_X1    g0146(.A(new_n263), .ZN(new_n347));
  AOI21_X1  g0147(.A(KEYINPUT67), .B1(new_n296), .B2(new_n254), .ZN(new_n348));
  OAI211_X1 g0148(.A(G232), .B(new_n267), .C1(new_n347), .C2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n256), .ZN(new_n350));
  INV_X1    g0150(.A(G223), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n273), .ZN(new_n352));
  INV_X1    g0152(.A(G226), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(G1698), .ZN(new_n354));
  AND2_X1   g0154(.A1(KEYINPUT3), .A2(G33), .ZN(new_n355));
  NOR2_X1   g0155(.A1(KEYINPUT3), .A2(G33), .ZN(new_n356));
  OAI211_X1 g0156(.A(new_n352), .B(new_n354), .C1(new_n355), .C2(new_n356), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n266), .A2(new_n211), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n267), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n349), .A2(new_n350), .A3(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(G200), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n349), .A2(new_n350), .ZN(new_n365));
  XNOR2_X1  g0165(.A(KEYINPUT81), .B(G190), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n360), .A2(KEYINPUT80), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT80), .ZN(new_n369));
  AOI211_X1 g0169(.A(new_n369), .B(new_n267), .C1(new_n357), .C2(new_n359), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n367), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n364), .B1(new_n365), .B2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT16), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT78), .ZN(new_n374));
  INV_X1    g0174(.A(G159), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n374), .B1(new_n288), .B2(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n317), .A2(KEYINPUT78), .A3(G159), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  AND2_X1   g0178(.A1(KEYINPUT68), .A2(G58), .ZN(new_n379));
  NOR2_X1   g0179(.A1(KEYINPUT68), .A2(G58), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n201), .B1(new_n381), .B2(G68), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n378), .B1(new_n382), .B2(new_n225), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n269), .A2(new_n225), .A3(new_n270), .ZN(new_n384));
  XNOR2_X1  g0184(.A(KEYINPUT77), .B(KEYINPUT7), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n269), .A2(KEYINPUT7), .A3(new_n225), .A4(new_n270), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n219), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n373), .B1(new_n383), .B2(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n280), .A2(G68), .A3(new_n281), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(new_n227), .ZN(new_n391));
  AOI22_X1  g0191(.A1(new_n391), .A2(G20), .B1(new_n376), .B2(new_n377), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n355), .A2(new_n356), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n393), .A2(new_n385), .A3(new_n225), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n384), .A2(KEYINPUT7), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n394), .A2(new_n395), .A3(G68), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n392), .A2(new_n396), .A3(KEYINPUT16), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n389), .A2(new_n292), .A3(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(G20), .B1(new_n258), .B2(new_n259), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n282), .A2(new_n399), .A3(new_n283), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT79), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n328), .A2(new_n292), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n282), .A2(new_n399), .A3(KEYINPUT79), .A4(new_n283), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n402), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n328), .A2(new_n284), .ZN(new_n406));
  AND2_X1   g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n372), .A2(KEYINPUT17), .A3(new_n398), .A4(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT17), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n398), .A2(new_n407), .ZN(new_n410));
  AOI22_X1  g0210(.A1(new_n269), .A2(new_n270), .B1(new_n351), .B2(new_n273), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n358), .B1(new_n411), .B2(new_n354), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n369), .B1(new_n412), .B2(new_n267), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n360), .A2(KEYINPUT80), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n366), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n256), .B1(new_n264), .B2(G232), .ZN(new_n416));
  AOI22_X1  g0216(.A1(new_n415), .A2(new_n416), .B1(new_n362), .B2(new_n363), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n409), .B1(new_n410), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n408), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n310), .B1(new_n413), .B2(new_n414), .ZN(new_n421));
  AOI22_X1  g0221(.A1(new_n421), .A2(new_n416), .B1(new_n362), .B2(new_n312), .ZN(new_n422));
  AOI21_X1  g0222(.A(KEYINPUT18), .B1(new_n410), .B2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n410), .A2(new_n422), .A3(KEYINPUT18), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n420), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT74), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n256), .A2(new_n428), .ZN(new_n429));
  OAI21_X1  g0229(.A(KEYINPUT74), .B1(new_n250), .B2(new_n255), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n271), .B1(G232), .B2(new_n273), .ZN(new_n432));
  NOR2_X1   g0232(.A1(G226), .A2(G1698), .ZN(new_n433));
  INV_X1    g0233(.A(G97), .ZN(new_n434));
  OAI22_X1  g0234(.A1(new_n432), .A2(new_n433), .B1(new_n266), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(new_n257), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n264), .A2(G238), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n431), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT13), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n431), .A2(new_n436), .A3(new_n437), .A4(KEYINPUT13), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n440), .A2(G169), .A3(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT76), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n442), .B1(new_n443), .B2(KEYINPUT14), .ZN(new_n444));
  AND2_X1   g0244(.A1(KEYINPUT75), .A2(KEYINPUT13), .ZN(new_n445));
  OR2_X1    g0245(.A1(new_n438), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n438), .A2(new_n445), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n446), .A2(G179), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n443), .A2(KEYINPUT14), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n443), .A2(KEYINPUT14), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n440), .A2(G169), .A3(new_n450), .A4(new_n441), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n444), .A2(new_n448), .A3(new_n449), .A4(new_n451), .ZN(new_n452));
  AOI22_X1  g0252(.A1(new_n285), .A2(G77), .B1(G20), .B2(new_n219), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n317), .A2(G50), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n293), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  XOR2_X1   g0255(.A(new_n455), .B(KEYINPUT11), .Z(new_n456));
  OAI21_X1  g0256(.A(new_n456), .B1(new_n219), .B2(new_n330), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n294), .A2(G68), .ZN(new_n458));
  XNOR2_X1  g0258(.A(new_n458), .B(KEYINPUT12), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n452), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n446), .A2(G190), .A3(new_n447), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n440), .A2(G200), .A3(new_n441), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n463), .A2(new_n460), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  NOR4_X1   g0266(.A1(new_n315), .A2(new_n346), .A3(new_n427), .A4(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(new_n225), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(KEYINPUT88), .ZN(new_n470));
  NOR2_X1   g0270(.A1(G97), .A2(G107), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(new_n211), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT88), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n468), .A2(new_n473), .A3(new_n225), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n470), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g0275(.A(G20), .B1(new_n269), .B2(new_n270), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(G68), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT19), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n478), .B1(new_n286), .B2(new_n434), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n475), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(new_n292), .ZN(new_n481));
  AND2_X1   g0281(.A1(new_n320), .A2(new_n324), .ZN(new_n482));
  OAI21_X1  g0282(.A(G33), .B1(new_n258), .B2(new_n259), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n403), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n325), .A2(new_n328), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n481), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(KEYINPUT89), .ZN(new_n487));
  AOI22_X1  g0287(.A1(new_n480), .A2(new_n292), .B1(new_n328), .B2(new_n325), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT89), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n488), .A2(new_n489), .A3(new_n484), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT66), .ZN(new_n492));
  INV_X1    g0292(.A(G1), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(KEYINPUT66), .A2(G1), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n253), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n496), .A2(new_n257), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n220), .A2(new_n273), .ZN(new_n498));
  INV_X1    g0298(.A(G244), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(G1698), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n498), .B(new_n500), .C1(new_n355), .C2(new_n356), .ZN(new_n501));
  NAND2_X1  g0301(.A1(G33), .A2(G116), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI22_X1  g0303(.A1(G250), .A2(new_n497), .B1(new_n503), .B2(new_n257), .ZN(new_n504));
  OAI211_X1 g0304(.A(G45), .B(G274), .C1(new_n258), .C2(new_n259), .ZN(new_n505));
  OAI21_X1  g0305(.A(KEYINPUT87), .B1(new_n505), .B2(new_n257), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT87), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n496), .A2(new_n507), .A3(G274), .A4(new_n267), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(G169), .B1(new_n504), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n497), .A2(G250), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n503), .A2(new_n257), .ZN(new_n512));
  AND3_X1   g0312(.A1(new_n509), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n510), .B1(new_n513), .B2(new_n342), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT90), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n509), .A2(new_n511), .A3(new_n512), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n515), .B1(new_n516), .B2(new_n279), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n504), .A2(KEYINPUT90), .A3(G190), .A4(new_n509), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n403), .A2(G87), .A3(new_n483), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n481), .A2(new_n520), .A3(new_n485), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n363), .B1(new_n504), .B2(new_n509), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n491), .A2(new_n514), .B1(new_n519), .B2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT85), .ZN(new_n525));
  OAI21_X1  g0325(.A(G45), .B1(new_n258), .B2(new_n259), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n252), .A2(KEYINPUT5), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT5), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(G41), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  OAI211_X1 g0330(.A(G257), .B(new_n267), .C1(new_n526), .C2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  XNOR2_X1  g0332(.A(KEYINPUT5), .B(G41), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n496), .A2(G274), .A3(new_n267), .A4(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(G33), .A2(G283), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  OAI211_X1 g0337(.A(G244), .B(new_n273), .C1(new_n355), .C2(new_n356), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT4), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n271), .A2(KEYINPUT4), .A3(G244), .A4(new_n273), .ZN(new_n541));
  OAI211_X1 g0341(.A(G250), .B(G1698), .C1(new_n355), .C2(new_n356), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(KEYINPUT84), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT84), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n271), .A2(new_n544), .A3(G250), .A4(G1698), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n540), .A2(new_n541), .A3(new_n543), .A4(new_n545), .ZN(new_n546));
  AOI211_X1 g0346(.A(new_n532), .B(new_n535), .C1(new_n546), .C2(new_n257), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n525), .B1(new_n547), .B2(new_n363), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT6), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n434), .A2(new_n334), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n549), .B1(new_n550), .B2(new_n471), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT82), .ZN(new_n552));
  NAND2_X1  g0352(.A1(KEYINPUT6), .A2(G97), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n552), .B1(new_n553), .B2(G107), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n334), .A2(KEYINPUT82), .A3(KEYINPUT6), .A4(G97), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n551), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n556), .A2(G20), .B1(G77), .B2(new_n317), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n386), .A2(new_n387), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(G107), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n293), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n294), .A2(G97), .ZN(new_n561));
  XNOR2_X1  g0361(.A(new_n561), .B(KEYINPUT83), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  AND3_X1   g0363(.A1(new_n403), .A2(G97), .A3(new_n483), .ZN(new_n564));
  NOR3_X1   g0364(.A1(new_n560), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n546), .A2(new_n257), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n566), .A2(new_n531), .A3(new_n534), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n567), .A2(KEYINPUT85), .A3(G200), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n547), .A2(G190), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n548), .A2(new_n565), .A3(new_n568), .A4(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(KEYINPUT86), .B1(new_n567), .B2(new_n310), .ZN(new_n571));
  INV_X1    g0371(.A(new_n564), .ZN(new_n572));
  AND2_X1   g0372(.A1(new_n557), .A2(new_n559), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n572), .B(new_n562), .C1(new_n573), .C2(new_n293), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n567), .A2(new_n312), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n535), .B1(new_n546), .B2(new_n257), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT86), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n576), .A2(new_n577), .A3(new_n342), .A4(new_n531), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n571), .A2(new_n574), .A3(new_n575), .A4(new_n578), .ZN(new_n579));
  AND3_X1   g0379(.A1(new_n524), .A2(new_n570), .A3(new_n579), .ZN(new_n580));
  OAI211_X1 g0380(.A(G257), .B(G1698), .C1(new_n355), .C2(new_n356), .ZN(new_n581));
  OAI211_X1 g0381(.A(G250), .B(new_n273), .C1(new_n355), .C2(new_n356), .ZN(new_n582));
  INV_X1    g0382(.A(G294), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n581), .B(new_n582), .C1(new_n266), .C2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n257), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n257), .B1(new_n496), .B2(new_n533), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(G264), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n585), .A2(new_n534), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n363), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n589), .B1(G190), .B2(new_n588), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n403), .A2(G107), .A3(new_n483), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n294), .A2(G107), .ZN(new_n592));
  XNOR2_X1  g0392(.A(new_n592), .B(KEYINPUT25), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n285), .A2(G116), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n225), .A2(G107), .ZN(new_n595));
  XNOR2_X1  g0395(.A(new_n595), .B(KEYINPUT23), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT22), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n597), .B1(new_n476), .B2(G87), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n225), .B(G87), .C1(new_n355), .C2(new_n356), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n599), .A2(KEYINPUT22), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n594), .B(new_n596), .C1(new_n598), .C2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT24), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g0403(.A(new_n599), .B(KEYINPUT22), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n604), .A2(KEYINPUT24), .A3(new_n594), .A4(new_n596), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n603), .A2(new_n605), .A3(new_n292), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n590), .A2(new_n591), .A3(new_n593), .A4(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n606), .A2(new_n591), .A3(new_n593), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n588), .A2(G179), .ZN(new_n609));
  AOI22_X1  g0409(.A1(new_n584), .A2(new_n257), .B1(new_n586), .B2(G264), .ZN(new_n610));
  AOI21_X1  g0410(.A(G169), .B1(new_n610), .B2(new_n534), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n608), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n607), .A2(new_n613), .ZN(new_n614));
  OR2_X1    g0414(.A1(KEYINPUT91), .A2(G303), .ZN(new_n615));
  NAND2_X1  g0415(.A1(KEYINPUT91), .A2(G303), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n615), .A2(new_n269), .A3(new_n270), .A4(new_n616), .ZN(new_n617));
  OAI211_X1 g0417(.A(G257), .B(new_n273), .C1(new_n355), .C2(new_n356), .ZN(new_n618));
  OAI211_X1 g0418(.A(G264), .B(G1698), .C1(new_n355), .C2(new_n356), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n617), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n257), .ZN(new_n621));
  OAI211_X1 g0421(.A(G270), .B(new_n267), .C1(new_n526), .C2(new_n530), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n621), .A2(new_n534), .A3(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(G116), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n328), .A2(new_n624), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n294), .A2(new_n293), .A3(new_n483), .A4(G116), .ZN(new_n626));
  AOI22_X1  g0426(.A1(new_n291), .A2(new_n224), .B1(G20), .B2(new_n624), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n536), .B(new_n225), .C1(G33), .C2(new_n434), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n627), .A2(KEYINPUT20), .A3(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(KEYINPUT20), .B1(new_n627), .B2(new_n628), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n625), .B(new_n626), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n623), .A2(G169), .A3(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT92), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT21), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n623), .A2(KEYINPUT92), .A3(new_n631), .A4(G169), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n623), .A2(KEYINPUT21), .A3(G169), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n621), .A2(G179), .A3(new_n534), .A4(new_n622), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n631), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n623), .A2(G200), .ZN(new_n642));
  INV_X1    g0442(.A(new_n631), .ZN(new_n643));
  OAI211_X1 g0443(.A(new_n642), .B(new_n643), .C1(new_n623), .C2(new_n367), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n637), .A2(new_n641), .A3(new_n644), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n614), .A2(new_n645), .ZN(new_n646));
  AND3_X1   g0446(.A1(new_n467), .A2(new_n580), .A3(new_n646), .ZN(G372));
  INV_X1    g0447(.A(new_n314), .ZN(new_n648));
  AND3_X1   g0448(.A1(new_n410), .A2(new_n422), .A3(KEYINPUT18), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n649), .A2(new_n423), .ZN(new_n650));
  INV_X1    g0450(.A(new_n465), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n651), .B1(new_n462), .B2(new_n344), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n650), .B1(new_n652), .B2(new_n420), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT96), .ZN(new_n654));
  OR2_X1    g0454(.A1(new_n305), .A2(new_n308), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n305), .A2(new_n308), .ZN(new_n656));
  AOI22_X1  g0456(.A1(new_n653), .A2(new_n654), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n652), .A2(new_n420), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(new_n426), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(KEYINPUT96), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n648), .B1(new_n657), .B2(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n613), .A2(new_n641), .A3(new_n637), .ZN(new_n662));
  XNOR2_X1  g0462(.A(new_n510), .B(KEYINPUT93), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n513), .A2(new_n342), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n663), .A2(new_n491), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n523), .A2(KEYINPUT94), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT94), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n667), .B1(new_n521), .B2(new_n522), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n666), .A2(new_n519), .A3(new_n668), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n662), .A2(new_n607), .A3(new_n665), .A4(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n570), .A2(new_n579), .ZN(new_n671));
  OR2_X1    g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n665), .A2(new_n669), .ZN(new_n673));
  NOR3_X1   g0473(.A1(new_n673), .A2(KEYINPUT26), .A3(new_n579), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n491), .A2(new_n514), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n519), .A2(new_n523), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(KEYINPUT26), .B1(new_n678), .B2(new_n579), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT95), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n665), .A2(new_n680), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n663), .A2(KEYINPUT95), .A3(new_n491), .A4(new_n664), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n672), .A2(new_n675), .A3(new_n679), .A4(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n467), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n661), .A2(new_n685), .ZN(G369));
  INV_X1    g0486(.A(G13), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n687), .A2(G20), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n296), .A2(new_n688), .ZN(new_n689));
  OR2_X1    g0489(.A1(new_n689), .A2(KEYINPUT27), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(KEYINPUT27), .ZN(new_n691));
  AND3_X1   g0491(.A1(new_n690), .A2(G213), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g0492(.A(KEYINPUT97), .B(G343), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n613), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n608), .A2(new_n695), .ZN(new_n697));
  XOR2_X1   g0497(.A(new_n697), .B(KEYINPUT98), .Z(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(new_n607), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n696), .B1(new_n699), .B2(new_n613), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n695), .B1(new_n637), .B2(new_n641), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n637), .A2(new_n641), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n694), .A2(new_n643), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n705), .B1(new_n645), .B2(new_n704), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n702), .B1(new_n706), .B2(G330), .ZN(new_n707));
  OAI22_X1  g0507(.A1(new_n701), .A2(new_n707), .B1(new_n613), .B2(new_n695), .ZN(G399));
  INV_X1    g0508(.A(new_n207), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(G41), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(G1), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n471), .A2(new_n211), .A3(new_n624), .ZN(new_n713));
  OAI22_X1  g0513(.A1(new_n712), .A2(new_n713), .B1(new_n228), .B2(new_n711), .ZN(new_n714));
  XNOR2_X1  g0514(.A(new_n714), .B(KEYINPUT28), .ZN(new_n715));
  OAI21_X1  g0515(.A(KEYINPUT26), .B1(new_n673), .B2(new_n579), .ZN(new_n716));
  INV_X1    g0516(.A(new_n579), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(new_n524), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n716), .B1(KEYINPUT26), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n683), .B1(new_n670), .B2(new_n671), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n694), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(KEYINPUT29), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n684), .A2(new_n694), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n722), .B1(new_n723), .B2(KEYINPUT29), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n580), .A2(new_n646), .A3(new_n694), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n513), .A2(new_n310), .ZN(new_n727));
  AND2_X1   g0527(.A1(new_n588), .A2(new_n623), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n727), .A2(new_n728), .A3(new_n567), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT30), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n585), .A2(new_n587), .ZN(new_n731));
  NOR3_X1   g0531(.A1(new_n639), .A2(new_n516), .A3(new_n731), .ZN(new_n732));
  AOI211_X1 g0532(.A(KEYINPUT99), .B(new_n730), .C1(new_n732), .C2(new_n547), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n639), .A2(new_n516), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n547), .A2(new_n734), .A3(new_n610), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT99), .ZN(new_n736));
  AOI21_X1  g0536(.A(KEYINPUT30), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n729), .B1(new_n733), .B2(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n738), .A2(KEYINPUT31), .A3(new_n695), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT100), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n727), .A2(new_n728), .A3(new_n740), .A4(new_n567), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  AND3_X1   g0542(.A1(new_n621), .A2(new_n534), .A3(new_n622), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n513), .A2(new_n743), .A3(G179), .A4(new_n610), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n736), .B1(new_n744), .B2(new_n567), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(new_n730), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n735), .A2(new_n736), .A3(KEYINPUT30), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n742), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n729), .A2(KEYINPUT100), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n694), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  OAI211_X1 g0550(.A(new_n726), .B(new_n739), .C1(new_n750), .C2(KEYINPUT31), .ZN(new_n751));
  AND3_X1   g0551(.A1(new_n751), .A2(KEYINPUT101), .A3(G330), .ZN(new_n752));
  AOI21_X1  g0552(.A(KEYINPUT101), .B1(new_n751), .B2(G330), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n725), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n715), .B1(new_n756), .B2(G1), .ZN(G364));
  OR2_X1    g0557(.A1(new_n706), .A2(G330), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n706), .A2(G330), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n712), .B1(G45), .B2(new_n688), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n758), .A2(new_n759), .A3(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n342), .A2(new_n225), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(G200), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n367), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n764), .A2(G190), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  OAI22_X1  g0568(.A1(new_n202), .A2(new_n766), .B1(new_n768), .B2(new_n219), .ZN(new_n769));
  INV_X1    g0569(.A(KEYINPUT32), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n225), .A2(G179), .ZN(new_n771));
  NOR2_X1   g0571(.A1(G190), .A2(G200), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(new_n375), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n769), .B1(new_n770), .B2(new_n774), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n771), .A2(new_n279), .A3(G200), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G107), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n778), .B1(new_n770), .B2(new_n774), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n771), .A2(G190), .A3(G200), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n763), .A2(new_n772), .ZN(new_n781));
  OAI221_X1 g0581(.A(new_n271), .B1(new_n211), .B2(new_n780), .C1(new_n781), .C2(new_n327), .ZN(new_n782));
  NOR3_X1   g0582(.A1(new_n279), .A2(G179), .A3(G200), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(new_n225), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  AOI211_X1 g0585(.A(new_n779), .B(new_n782), .C1(G97), .C2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n381), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n763), .A2(new_n363), .A3(new_n366), .ZN(new_n788));
  OAI211_X1 g0588(.A(new_n775), .B(new_n786), .C1(new_n787), .C2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(G322), .ZN(new_n790));
  OAI221_X1 g0590(.A(new_n393), .B1(new_n583), .B2(new_n784), .C1(new_n788), .C2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n773), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n791), .B1(G329), .B2(new_n792), .ZN(new_n793));
  XOR2_X1   g0593(.A(KEYINPUT104), .B(G326), .Z(new_n794));
  NAND2_X1  g0594(.A1(new_n765), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(G283), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n795), .B1(new_n796), .B2(new_n776), .ZN(new_n797));
  INV_X1    g0597(.A(new_n780), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n797), .B1(G303), .B2(new_n798), .ZN(new_n799));
  XOR2_X1   g0599(.A(KEYINPUT33), .B(G317), .Z(new_n800));
  OAI211_X1 g0600(.A(new_n793), .B(new_n799), .C1(new_n768), .C2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(G311), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n781), .A2(new_n802), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n789), .B1(new_n801), .B2(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n224), .B1(G20), .B2(new_n312), .ZN(new_n805));
  NOR2_X1   g0605(.A1(G13), .A2(G33), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n807), .A2(G20), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(new_n805), .ZN(new_n809));
  XOR2_X1   g0609(.A(new_n809), .B(KEYINPUT103), .Z(new_n810));
  NOR2_X1   g0610(.A1(new_n709), .A2(new_n393), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(G355), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n242), .A2(G45), .ZN(new_n813));
  XOR2_X1   g0613(.A(new_n813), .B(KEYINPUT102), .Z(new_n814));
  NOR2_X1   g0614(.A1(new_n709), .A2(new_n271), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n815), .B1(G45), .B2(new_n228), .ZN(new_n816));
  OAI221_X1 g0616(.A(new_n812), .B1(G116), .B2(new_n207), .C1(new_n814), .C2(new_n816), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n804), .A2(new_n805), .B1(new_n810), .B2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n808), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n818), .B1(new_n706), .B2(new_n819), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n762), .B1(new_n820), .B2(new_n761), .ZN(G396));
  NAND2_X1  g0621(.A1(new_n331), .A2(new_n695), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n340), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(new_n344), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n344), .A2(new_n695), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  NOR3_X1   g0628(.A1(new_n752), .A2(new_n753), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n751), .A2(G330), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT101), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n751), .A2(KEYINPUT101), .A3(G330), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n827), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n829), .A2(new_n834), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n835), .B(new_n723), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(new_n761), .ZN(new_n837));
  INV_X1    g0637(.A(new_n781), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n767), .A2(G150), .B1(new_n838), .B2(G159), .ZN(new_n839));
  INV_X1    g0639(.A(G137), .ZN(new_n840));
  INV_X1    g0640(.A(G143), .ZN(new_n841));
  OAI221_X1 g0641(.A(new_n839), .B1(new_n840), .B2(new_n766), .C1(new_n841), .C2(new_n788), .ZN(new_n842));
  XNOR2_X1  g0642(.A(KEYINPUT106), .B(KEYINPUT34), .ZN(new_n843));
  XNOR2_X1  g0643(.A(new_n842), .B(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(G132), .ZN(new_n845));
  OAI22_X1  g0645(.A1(new_n784), .A2(new_n787), .B1(new_n845), .B2(new_n773), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n271), .B1(new_n776), .B2(new_n219), .C1(new_n202), .C2(new_n780), .ZN(new_n847));
  NOR3_X1   g0647(.A1(new_n844), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n767), .A2(G283), .B1(new_n838), .B2(G116), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT105), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n765), .A2(G303), .ZN(new_n852));
  AOI22_X1  g0652(.A1(new_n785), .A2(G97), .B1(new_n798), .B2(G107), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n271), .B1(new_n777), .B2(G87), .ZN(new_n855));
  OAI221_X1 g0655(.A(new_n855), .B1(new_n583), .B2(new_n788), .C1(new_n849), .C2(new_n850), .ZN(new_n856));
  AOI211_X1 g0656(.A(new_n854), .B(new_n856), .C1(G311), .C2(new_n792), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n805), .B1(new_n848), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n827), .A2(new_n806), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n805), .A2(new_n806), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(new_n327), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n858), .A2(new_n760), .A3(new_n859), .A4(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n837), .A2(new_n862), .ZN(G384));
  OAI211_X1 g0663(.A(new_n749), .B(new_n741), .C1(new_n733), .C2(new_n737), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(new_n695), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT31), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n864), .A2(KEYINPUT31), .A3(new_n695), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n867), .A2(new_n726), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n461), .A2(new_n695), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n462), .A2(new_n465), .A3(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n452), .A2(new_n461), .A3(new_n695), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n869), .A2(new_n828), .A3(new_n873), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n371), .A2(new_n365), .ZN(new_n875));
  AOI21_X1  g0675(.A(G200), .B1(new_n416), .B2(new_n361), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n398), .B(new_n407), .C1(new_n875), .C2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n410), .A2(new_n422), .ZN(new_n878));
  AND2_X1   g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT107), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT37), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n410), .A2(new_n692), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n879), .A2(new_n880), .A3(new_n881), .A4(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n877), .A2(new_n878), .A3(new_n882), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(KEYINPUT37), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n877), .A2(new_n878), .A3(new_n882), .A4(new_n881), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(KEYINPUT107), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n883), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  OAI211_X1 g0688(.A(new_n410), .B(new_n692), .C1(new_n650), .C2(new_n419), .ZN(new_n889));
  AOI21_X1  g0689(.A(KEYINPUT38), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n397), .A2(new_n292), .ZN(new_n891));
  AOI21_X1  g0691(.A(KEYINPUT16), .B1(new_n392), .B2(new_n396), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n407), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n692), .B(new_n893), .C1(new_n650), .C2(new_n419), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n893), .B1(new_n422), .B2(new_n692), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n895), .A2(new_n877), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n886), .B1(new_n896), .B2(new_n881), .ZN(new_n897));
  AND3_X1   g0697(.A1(new_n894), .A2(KEYINPUT38), .A3(new_n897), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n890), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(KEYINPUT40), .B1(new_n874), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n894), .A2(new_n897), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT38), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n894), .A2(KEYINPUT38), .A3(new_n897), .ZN(new_n904));
  AOI21_X1  g0704(.A(KEYINPUT40), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n524), .A2(new_n570), .A3(new_n579), .ZN(new_n906));
  NOR4_X1   g0706(.A1(new_n906), .A2(new_n614), .A3(new_n645), .A4(new_n695), .ZN(new_n907));
  AOI21_X1  g0707(.A(KEYINPUT31), .B1(new_n864), .B2(new_n695), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n827), .B1(new_n909), .B2(new_n868), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n905), .A2(new_n910), .A3(new_n873), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n900), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(G330), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n467), .A2(G330), .A3(new_n869), .ZN(new_n914));
  AND2_X1   g0714(.A1(new_n467), .A2(new_n869), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n913), .A2(new_n914), .B1(new_n912), .B2(new_n915), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n462), .A2(new_n695), .ZN(new_n917));
  NOR3_X1   g0717(.A1(new_n890), .A2(new_n898), .A3(KEYINPUT39), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT39), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n919), .B1(new_n903), .B2(new_n904), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n917), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n679), .B(new_n683), .C1(new_n670), .C2(new_n671), .ZN(new_n922));
  OAI211_X1 g0722(.A(new_n694), .B(new_n824), .C1(new_n922), .C2(new_n674), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n826), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n903), .A2(new_n904), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n924), .A2(new_n873), .A3(new_n925), .ZN(new_n926));
  OR2_X1    g0726(.A1(new_n426), .A2(new_n692), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n921), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n916), .B(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n724), .A2(new_n467), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n661), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n929), .B(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n296), .B2(new_n688), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n624), .B1(new_n556), .B2(KEYINPUT35), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n934), .B(new_n226), .C1(KEYINPUT35), .C2(new_n556), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(KEYINPUT36), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n229), .A2(G77), .A3(new_n390), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(G50), .B2(new_n219), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n687), .ZN(new_n939));
  OAI211_X1 g0739(.A(new_n933), .B(new_n936), .C1(new_n296), .C2(new_n939), .ZN(G367));
  NAND2_X1  g0740(.A1(new_n777), .A2(G97), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT109), .ZN(new_n942));
  OAI22_X1  g0742(.A1(new_n781), .A2(new_n796), .B1(new_n334), .B2(new_n784), .ZN(new_n943));
  INV_X1    g0743(.A(new_n788), .ZN(new_n944));
  AND2_X1   g0744(.A1(new_n615), .A2(new_n616), .ZN(new_n945));
  AOI22_X1  g0745(.A1(G311), .A2(new_n765), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  OAI221_X1 g0746(.A(new_n941), .B1(new_n942), .B2(new_n943), .C1(new_n946), .C2(KEYINPUT110), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(KEYINPUT110), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n943), .A2(new_n942), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n798), .A2(G116), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n950), .B(KEYINPUT46), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n271), .B1(new_n767), .B2(G294), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n948), .A2(new_n949), .A3(new_n951), .A4(new_n952), .ZN(new_n953));
  AOI211_X1 g0753(.A(new_n947), .B(new_n953), .C1(G317), .C2(new_n792), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n944), .A2(G150), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n785), .A2(G68), .ZN(new_n956));
  OAI221_X1 g0756(.A(new_n956), .B1(new_n202), .B2(new_n781), .C1(new_n766), .C2(new_n841), .ZN(new_n957));
  OAI22_X1  g0757(.A1(new_n787), .A2(new_n780), .B1(new_n840), .B2(new_n773), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n271), .B1(new_n958), .B2(KEYINPUT111), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(KEYINPUT111), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n777), .A2(G77), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n960), .B(new_n961), .C1(new_n768), .C2(new_n375), .ZN(new_n962));
  NOR3_X1   g0762(.A1(new_n957), .A2(new_n959), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n954), .B1(new_n955), .B2(new_n963), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n964), .B(KEYINPUT47), .Z(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n805), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n694), .B1(new_n520), .B2(new_n488), .ZN(new_n967));
  OR2_X1    g0767(.A1(new_n673), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n681), .A2(new_n682), .A3(new_n967), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n968), .A2(new_n808), .A3(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n815), .ZN(new_n971));
  OAI221_X1 g0771(.A(new_n810), .B1(new_n207), .B2(new_n325), .C1(new_n238), .C2(new_n971), .ZN(new_n972));
  NAND4_X1  g0772(.A1(new_n966), .A2(new_n760), .A3(new_n970), .A4(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n700), .B(new_n707), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n755), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n696), .B1(new_n700), .B2(new_n702), .ZN(new_n978));
  INV_X1    g0778(.A(new_n671), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n565), .B2(new_n694), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n717), .A2(new_n695), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n978), .A2(new_n982), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n983), .B(KEYINPUT45), .Z(new_n984));
  NOR2_X1   g0784(.A1(new_n978), .A2(new_n982), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(KEYINPUT44), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n701), .A2(new_n759), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n977), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(new_n756), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n710), .B(KEYINPUT41), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n493), .B1(new_n688), .B2(G45), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n700), .A2(new_n979), .A3(new_n702), .ZN(new_n995));
  XOR2_X1   g0795(.A(KEYINPUT108), .B(KEYINPUT42), .Z(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n579), .B1(new_n980), .B2(new_n613), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n999), .A2(new_n694), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n995), .A2(new_n997), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n998), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n968), .A2(new_n969), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(KEYINPUT43), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n1003), .A2(KEYINPUT43), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NOR3_X1   g0807(.A1(new_n1002), .A2(KEYINPUT43), .A3(new_n1003), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n988), .A2(new_n982), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1009), .B(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n974), .B1(new_n994), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(G387));
  AOI22_X1  g0813(.A1(new_n767), .A2(G311), .B1(new_n838), .B2(new_n945), .ZN(new_n1014));
  INV_X1    g0814(.A(G317), .ZN(new_n1015));
  XOR2_X1   g0815(.A(KEYINPUT114), .B(G322), .Z(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n1014), .B1(new_n1015), .B2(new_n788), .C1(new_n766), .C2(new_n1017), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n1018), .B(KEYINPUT48), .Z(new_n1019));
  OAI22_X1  g0819(.A1(new_n784), .A2(new_n796), .B1(new_n780), .B2(new_n583), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT113), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  AND2_X1   g0822(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1023));
  NOR3_X1   g0823(.A1(new_n1019), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n393), .B1(new_n1024), .B2(KEYINPUT49), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1024), .A2(KEYINPUT49), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1026), .B1(new_n624), .B2(new_n776), .ZN(new_n1027));
  AOI211_X1 g0827(.A(new_n1025), .B(new_n1027), .C1(new_n792), .C2(new_n794), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n765), .A2(G159), .B1(new_n482), .B2(new_n785), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1029), .B1(new_n202), .B2(new_n788), .C1(new_n284), .C2(new_n768), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n941), .B1(new_n327), .B2(new_n780), .C1(new_n287), .C2(new_n773), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n781), .A2(new_n219), .ZN(new_n1032));
  NOR4_X1   g0832(.A1(new_n1030), .A2(new_n393), .A3(new_n1031), .A4(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n805), .B1(new_n1028), .B2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n971), .B1(new_n235), .B2(G45), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1035), .B1(new_n713), .B2(new_n811), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n316), .A2(new_n202), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT50), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n253), .B1(new_n219), .B2(new_n327), .ZN(new_n1039));
  NOR3_X1   g0839(.A1(new_n1038), .A2(new_n713), .A3(new_n1039), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n1036), .A2(new_n1040), .B1(G107), .B2(new_n207), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n761), .B1(new_n1041), .B2(new_n810), .ZN(new_n1042));
  XOR2_X1   g0842(.A(new_n1042), .B(KEYINPUT112), .Z(new_n1043));
  OAI211_X1 g0843(.A(new_n1034), .B(new_n1043), .C1(new_n700), .C2(new_n819), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n710), .B1(new_n756), .B2(new_n975), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1044), .B1(new_n993), .B2(new_n976), .C1(new_n977), .C2(new_n1045), .ZN(G393));
  XOR2_X1   g0846(.A(new_n987), .B(new_n988), .Z(new_n1047));
  OAI211_X1 g0847(.A(new_n710), .B(new_n989), .C1(new_n1047), .C2(new_n977), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n778), .B1(new_n796), .B2(new_n780), .C1(new_n773), .C2(new_n1017), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n766), .A2(new_n1015), .B1(new_n802), .B2(new_n788), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT52), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n271), .B1(new_n838), .B2(G294), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n1051), .B(new_n1052), .C1(new_n624), .C2(new_n784), .ZN(new_n1053));
  AOI211_X1 g0853(.A(new_n1049), .B(new_n1053), .C1(new_n945), .C2(new_n767), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT116), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n271), .B1(new_n773), .B2(new_n841), .C1(new_n219), .C2(new_n780), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(G150), .A2(new_n765), .B1(new_n944), .B2(G159), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(KEYINPUT115), .B(KEYINPUT51), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1057), .B(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n785), .A2(G77), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n767), .A2(G50), .B1(G87), .B2(new_n777), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n1056), .B(new_n1062), .C1(new_n316), .C2(new_n838), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n805), .B1(new_n1055), .B2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n980), .A2(new_n808), .A3(new_n981), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n810), .B1(new_n434), .B2(new_n207), .C1(new_n245), .C2(new_n971), .ZN(new_n1066));
  AND4_X1   g0866(.A1(new_n760), .A2(new_n1064), .A3(new_n1065), .A4(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n993), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1067), .B1(new_n1047), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1048), .A2(new_n1069), .ZN(G390));
  INV_X1    g0870(.A(G330), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n874), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n882), .B1(new_n420), .B2(new_n426), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n886), .B(new_n880), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1074), .B1(new_n1075), .B2(new_n885), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n919), .B(new_n904), .C1(new_n1076), .C2(KEYINPUT38), .ZN(new_n1077));
  AOI21_X1  g0877(.A(KEYINPUT38), .B1(new_n894), .B2(new_n897), .ZN(new_n1078));
  OAI21_X1  g0878(.A(KEYINPUT39), .B1(new_n898), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n924), .A2(new_n873), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n917), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1080), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1082), .B1(new_n890), .B2(new_n898), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n694), .B(new_n824), .C1(new_n719), .C2(new_n720), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n826), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1084), .B1(new_n1086), .B2(new_n873), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1073), .B1(new_n1083), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n873), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(new_n923), .B2(new_n826), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1079), .B(new_n1077), .C1(new_n1090), .C2(new_n917), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1087), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n828), .B(new_n873), .C1(new_n752), .C2(new_n753), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1088), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n1068), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1077), .A2(new_n806), .A3(new_n1079), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n271), .B1(new_n838), .B2(G97), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n1098), .B1(new_n211), .B2(new_n780), .C1(new_n766), .C2(new_n796), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n776), .A2(new_n219), .B1(new_n773), .B2(new_n583), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n944), .A2(G116), .B1(KEYINPUT118), .B2(new_n1100), .ZN(new_n1101));
  OAI221_X1 g0901(.A(new_n1101), .B1(KEYINPUT118), .B2(new_n1100), .C1(new_n334), .C2(new_n768), .ZN(new_n1102));
  AOI211_X1 g0902(.A(new_n1099), .B(new_n1102), .C1(G77), .C2(new_n785), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n780), .A2(new_n287), .ZN(new_n1104));
  XOR2_X1   g0904(.A(KEYINPUT117), .B(KEYINPUT53), .Z(new_n1105));
  XNOR2_X1  g0905(.A(new_n1104), .B(new_n1105), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n785), .A2(G159), .B1(new_n777), .B2(G50), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n1106), .B(new_n1107), .C1(new_n768), .C2(new_n840), .ZN(new_n1108));
  XOR2_X1   g0908(.A(KEYINPUT54), .B(G143), .Z(new_n1109));
  AOI21_X1  g0909(.A(new_n393), .B1(new_n838), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(G128), .ZN(new_n1111));
  OAI221_X1 g0911(.A(new_n1110), .B1(new_n845), .B2(new_n788), .C1(new_n766), .C2(new_n1111), .ZN(new_n1112));
  AOI211_X1 g0912(.A(new_n1108), .B(new_n1112), .C1(G125), .C2(new_n792), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n805), .B1(new_n1103), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n284), .A2(new_n860), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n1097), .A2(new_n760), .A3(new_n1114), .A4(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n910), .A2(G330), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(new_n1089), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1086), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1094), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n828), .B1(new_n752), .B2(new_n753), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1072), .B1(new_n1121), .B2(new_n1089), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n924), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1120), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n930), .A2(new_n661), .A3(new_n914), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  NOR3_X1   g0926(.A1(new_n1083), .A2(new_n1087), .A3(new_n1094), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1072), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n1124), .B(new_n1126), .C1(new_n1127), .C2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(new_n710), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1132));
  AND2_X1   g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1096), .B(new_n1116), .C1(new_n1130), .C2(new_n1133), .ZN(G378));
  XNOR2_X1  g0934(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT121), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n315), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n302), .A2(new_n692), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n648), .B1(new_n655), .B2(new_n656), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(KEYINPUT121), .ZN(new_n1141));
  AND3_X1   g0941(.A1(new_n1138), .A2(new_n1139), .A3(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1139), .B1(new_n1138), .B2(new_n1141), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1136), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1139), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1141), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n1140), .A2(KEYINPUT121), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1145), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1138), .A2(new_n1139), .A3(new_n1141), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1148), .A2(new_n1135), .A3(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1144), .A2(new_n1150), .A3(new_n806), .ZN(new_n1151));
  OAI221_X1 g0951(.A(new_n956), .B1(new_n327), .B2(new_n780), .C1(new_n781), .C2(new_n325), .ZN(new_n1152));
  OAI221_X1 g0952(.A(new_n393), .B1(new_n773), .B2(new_n796), .C1(new_n787), .C2(new_n776), .ZN(new_n1153));
  NOR3_X1   g0953(.A1(new_n1152), .A2(G41), .A3(new_n1153), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(G116), .A2(new_n765), .B1(new_n944), .B2(G107), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1154), .B(new_n1155), .C1(new_n434), .C2(new_n768), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT58), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT119), .ZN(new_n1158));
  AOI21_X1  g0958(.A(G50), .B1(new_n270), .B2(new_n252), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n1156), .A2(new_n1157), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n798), .A2(new_n1109), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1161), .B1(new_n768), .B2(new_n845), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n765), .A2(G125), .ZN(new_n1163));
  OAI221_X1 g0963(.A(new_n1163), .B1(new_n1111), .B2(new_n788), .C1(new_n840), .C2(new_n781), .ZN(new_n1164));
  AOI211_X1 g0964(.A(new_n1162), .B(new_n1164), .C1(G150), .C2(new_n785), .ZN(new_n1165));
  XOR2_X1   g0965(.A(new_n1165), .B(KEYINPUT59), .Z(new_n1166));
  AOI21_X1  g0966(.A(G41), .B1(new_n777), .B2(G159), .ZN(new_n1167));
  OR2_X1    g0967(.A1(KEYINPUT120), .A2(G124), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(KEYINPUT120), .A2(G124), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n792), .A2(new_n1168), .A3(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1167), .A2(new_n266), .A3(new_n1170), .ZN(new_n1171));
  OAI221_X1 g0971(.A(new_n1160), .B1(new_n1157), .B2(new_n1156), .C1(new_n1166), .C2(new_n1171), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1159), .A2(new_n1158), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n805), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n860), .A2(new_n202), .ZN(new_n1175));
  AND4_X1   g0975(.A1(new_n760), .A2(new_n1151), .A3(new_n1174), .A4(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1144), .A2(new_n1150), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1071), .B1(new_n900), .B2(new_n911), .ZN(new_n1178));
  AND2_X1   g0978(.A1(new_n928), .A2(new_n1178), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n928), .A2(new_n1178), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1177), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  AND2_X1   g0981(.A1(new_n926), .A2(new_n927), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n913), .A2(new_n921), .A3(new_n1182), .ZN(new_n1183));
  AND2_X1   g0983(.A1(new_n1144), .A2(new_n1150), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n928), .A2(new_n1178), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1183), .A2(new_n1184), .A3(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1181), .A2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1176), .B1(new_n1187), .B2(new_n1068), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n1129), .A2(new_n1126), .B1(new_n1181), .B2(new_n1186), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n710), .B1(new_n1189), .B2(KEYINPUT57), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1073), .B1(new_n834), .B2(new_n873), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n873), .B1(new_n910), .B2(G330), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(new_n834), .B2(new_n873), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n924), .A2(new_n1191), .B1(new_n1193), .B2(new_n1119), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1126), .B1(new_n1132), .B2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1195), .A2(new_n1187), .A3(KEYINPUT57), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1188), .B1(new_n1190), .B2(new_n1197), .ZN(G375));
  OAI211_X1 g0998(.A(new_n1125), .B(new_n1120), .C1(new_n1123), .C2(new_n1122), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1131), .A2(new_n991), .A3(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1089), .A2(new_n806), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n767), .A2(new_n1109), .B1(new_n838), .B2(G150), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n1202), .B1(new_n845), .B2(new_n766), .C1(new_n787), .C2(new_n776), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n944), .A2(G137), .B1(G128), .B2(new_n792), .ZN(new_n1204));
  OAI221_X1 g1004(.A(new_n1204), .B1(new_n202), .B2(new_n784), .C1(new_n375), .C2(new_n780), .ZN(new_n1205));
  NOR3_X1   g1005(.A1(new_n1203), .A2(new_n1205), .A3(new_n393), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n838), .A2(G107), .B1(new_n482), .B2(new_n785), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1207), .B1(new_n624), .B2(new_n768), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n271), .B1(new_n944), .B2(G283), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n798), .A2(G97), .B1(new_n792), .B2(G303), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1209), .A2(new_n961), .A3(new_n1210), .ZN(new_n1211));
  AOI211_X1 g1011(.A(new_n1208), .B(new_n1211), .C1(G294), .C2(new_n765), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n805), .B1(new_n1206), .B2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n860), .A2(new_n219), .ZN(new_n1214));
  AND4_X1   g1014(.A1(new_n760), .A2(new_n1201), .A3(new_n1213), .A4(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(new_n1124), .B2(new_n1068), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1200), .A2(new_n1216), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(new_n1217), .B(KEYINPUT122), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(G381));
  INV_X1    g1019(.A(G375), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1130), .A2(new_n1133), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1096), .A2(new_n1116), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1220), .A2(new_n1223), .ZN(new_n1224));
  NOR3_X1   g1024(.A1(new_n1224), .A2(G396), .A3(G393), .ZN(new_n1225));
  NOR3_X1   g1025(.A1(G387), .A2(G381), .A3(G390), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1225), .A2(new_n837), .A3(new_n862), .A4(new_n1226), .ZN(G407));
  OAI211_X1 g1027(.A(G407), .B(G213), .C1(new_n693), .C2(new_n1224), .ZN(G409));
  INV_X1    g1028(.A(KEYINPUT123), .ZN(new_n1229));
  INV_X1    g1029(.A(G213), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n693), .A2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1195), .A2(new_n1187), .A3(new_n991), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1188), .A2(new_n1233), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1232), .B1(new_n1234), .B2(G378), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(G378), .B2(G375), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT60), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1199), .A2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1191), .A2(new_n924), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1239), .A2(KEYINPUT60), .A3(new_n1125), .A4(new_n1120), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1238), .A2(new_n710), .A3(new_n1131), .A4(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(new_n1216), .ZN(new_n1242));
  INV_X1    g1042(.A(G384), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(G384), .A2(new_n1241), .A3(new_n1216), .ZN(new_n1245));
  AND2_X1   g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1229), .B1(new_n1236), .B2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT57), .ZN(new_n1248));
  NOR3_X1   g1048(.A1(new_n1179), .A2(new_n1180), .A3(new_n1177), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1184), .B1(new_n1183), .B2(new_n1185), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1125), .B1(new_n1095), .B2(new_n1124), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1248), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1253), .A2(new_n710), .A3(new_n1196), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1223), .B1(new_n1254), .B2(new_n1188), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1256));
  NOR4_X1   g1056(.A1(new_n1255), .A2(new_n1235), .A3(KEYINPUT123), .A4(new_n1256), .ZN(new_n1257));
  NOR3_X1   g1057(.A1(new_n1247), .A2(new_n1257), .A3(KEYINPUT62), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(G375), .A2(G378), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1235), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1259), .A2(new_n1260), .A3(new_n1246), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(KEYINPUT62), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT61), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1231), .A2(G2897), .ZN(new_n1264));
  XOR2_X1   g1064(.A(new_n1264), .B(KEYINPUT124), .Z(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1246), .A2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1256), .A2(new_n1265), .ZN(new_n1268));
  OAI211_X1 g1068(.A(new_n1267), .B(new_n1268), .C1(new_n1255), .C2(new_n1235), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1262), .A2(new_n1263), .A3(new_n1269), .ZN(new_n1270));
  OAI21_X1  g1070(.A(KEYINPUT127), .B1(new_n1258), .B2(new_n1270), .ZN(new_n1271));
  XNOR2_X1  g1071(.A(G393), .B(G396), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT125), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1273), .B1(new_n1048), .B2(new_n1069), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1272), .B1(G387), .B2(new_n1274), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1012), .B1(G390), .B2(KEYINPUT125), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1275), .B1(new_n1274), .B2(new_n1276), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(G387), .A2(KEYINPUT126), .A3(new_n1069), .A4(new_n1048), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT126), .ZN(new_n1279));
  OAI21_X1  g1079(.A(G390), .B1(new_n1012), .B2(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1278), .A2(new_n1272), .A3(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1277), .A2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1261), .A2(KEYINPUT123), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT62), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1236), .A2(new_n1229), .A3(new_n1246), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1284), .A2(new_n1285), .A3(new_n1286), .ZN(new_n1287));
  AND2_X1   g1087(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1236), .ZN(new_n1289));
  AOI21_X1  g1089(.A(KEYINPUT61), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT127), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1287), .A2(new_n1290), .A3(new_n1291), .A4(new_n1262), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1271), .A2(new_n1283), .A3(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT63), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1294), .B1(new_n1247), .B2(new_n1257), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1236), .A2(KEYINPUT63), .A3(new_n1246), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1282), .A2(new_n1295), .A3(new_n1290), .A4(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1293), .A2(new_n1297), .ZN(G405));
  NAND2_X1  g1098(.A1(new_n1224), .A2(new_n1259), .ZN(new_n1299));
  XNOR2_X1  g1099(.A(new_n1299), .B(new_n1246), .ZN(new_n1300));
  XNOR2_X1  g1100(.A(new_n1300), .B(new_n1282), .ZN(G402));
endmodule


