

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U558 ( .A1(G651), .A2(G543), .ZN(n801) );
  OR2_X1 U559 ( .A1(n704), .A2(n703), .ZN(n705) );
  AND2_X1 U560 ( .A1(n624), .A2(n623), .ZN(n626) );
  NOR2_X1 U561 ( .A1(n524), .A2(n745), .ZN(n521) );
  XNOR2_X1 U562 ( .A(KEYINPUT40), .B(KEYINPUT107), .ZN(n522) );
  XOR2_X1 U563 ( .A(n656), .B(n655), .Z(n523) );
  AND2_X1 U564 ( .A1(n985), .A2(n767), .ZN(n524) );
  OR2_X1 U565 ( .A1(n717), .A2(n716), .ZN(n525) );
  AND2_X1 U566 ( .A1(n714), .A2(n713), .ZN(n526) );
  INV_X1 U567 ( .A(KEYINPUT29), .ZN(n655) );
  INV_X1 U568 ( .A(n975), .ZN(n703) );
  OR2_X1 U569 ( .A1(n706), .A2(n705), .ZN(n714) );
  XNOR2_X1 U570 ( .A(n612), .B(KEYINPUT14), .ZN(n613) );
  XNOR2_X1 U571 ( .A(n614), .B(n613), .ZN(n624) );
  XOR2_X1 U572 ( .A(KEYINPUT17), .B(n527), .Z(n886) );
  XNOR2_X1 U573 ( .A(n626), .B(n625), .ZN(n981) );
  NOR2_X1 U574 ( .A1(G2104), .A2(G2105), .ZN(n527) );
  NAND2_X1 U575 ( .A1(G138), .A2(n886), .ZN(n529) );
  INV_X1 U576 ( .A(G2105), .ZN(n530) );
  AND2_X1 U577 ( .A1(n530), .A2(G2104), .ZN(n887) );
  NAND2_X1 U578 ( .A1(G102), .A2(n887), .ZN(n528) );
  NAND2_X1 U579 ( .A1(n529), .A2(n528), .ZN(n534) );
  NOR2_X1 U580 ( .A1(G2104), .A2(n530), .ZN(n890) );
  NAND2_X1 U581 ( .A1(G126), .A2(n890), .ZN(n532) );
  AND2_X1 U582 ( .A1(G2104), .A2(G2105), .ZN(n891) );
  NAND2_X1 U583 ( .A1(G114), .A2(n891), .ZN(n531) );
  NAND2_X1 U584 ( .A1(n532), .A2(n531), .ZN(n533) );
  NOR2_X1 U585 ( .A1(n534), .A2(n533), .ZN(G164) );
  NAND2_X1 U586 ( .A1(n886), .A2(G137), .ZN(n537) );
  NAND2_X1 U587 ( .A1(G101), .A2(n887), .ZN(n535) );
  XOR2_X1 U588 ( .A(KEYINPUT23), .B(n535), .Z(n536) );
  NAND2_X1 U589 ( .A1(n537), .A2(n536), .ZN(n541) );
  NAND2_X1 U590 ( .A1(G125), .A2(n890), .ZN(n539) );
  NAND2_X1 U591 ( .A1(G113), .A2(n891), .ZN(n538) );
  NAND2_X1 U592 ( .A1(n539), .A2(n538), .ZN(n540) );
  NOR2_X1 U593 ( .A1(n541), .A2(n540), .ZN(G160) );
  XOR2_X1 U594 ( .A(G543), .B(KEYINPUT0), .Z(n582) );
  NOR2_X1 U595 ( .A1(G651), .A2(n582), .ZN(n797) );
  NAND2_X1 U596 ( .A1(n797), .A2(G52), .ZN(n544) );
  XNOR2_X1 U597 ( .A(G651), .B(KEYINPUT65), .ZN(n546) );
  NOR2_X1 U598 ( .A1(G543), .A2(n546), .ZN(n542) );
  XOR2_X2 U599 ( .A(KEYINPUT1), .B(n542), .Z(n798) );
  NAND2_X1 U600 ( .A1(G64), .A2(n798), .ZN(n543) );
  NAND2_X1 U601 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U602 ( .A(KEYINPUT66), .B(n545), .ZN(n551) );
  NAND2_X1 U603 ( .A1(G90), .A2(n801), .ZN(n548) );
  NOR2_X2 U604 ( .A1(n582), .A2(n546), .ZN(n805) );
  NAND2_X1 U605 ( .A1(G77), .A2(n805), .ZN(n547) );
  NAND2_X1 U606 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U607 ( .A(KEYINPUT9), .B(n549), .Z(n550) );
  NOR2_X1 U608 ( .A1(n551), .A2(n550), .ZN(G171) );
  NAND2_X1 U609 ( .A1(n801), .A2(G91), .ZN(n552) );
  XOR2_X1 U610 ( .A(KEYINPUT67), .B(n552), .Z(n554) );
  NAND2_X1 U611 ( .A1(G78), .A2(n805), .ZN(n553) );
  NAND2_X1 U612 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U613 ( .A(KEYINPUT68), .B(n555), .Z(n559) );
  NAND2_X1 U614 ( .A1(n798), .A2(G65), .ZN(n557) );
  NAND2_X1 U615 ( .A1(n797), .A2(G53), .ZN(n556) );
  AND2_X1 U616 ( .A1(n557), .A2(n556), .ZN(n558) );
  NAND2_X1 U617 ( .A1(n559), .A2(n558), .ZN(G299) );
  NAND2_X1 U618 ( .A1(n801), .A2(G89), .ZN(n560) );
  XNOR2_X1 U619 ( .A(n560), .B(KEYINPUT4), .ZN(n562) );
  NAND2_X1 U620 ( .A1(G76), .A2(n805), .ZN(n561) );
  NAND2_X1 U621 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U622 ( .A(KEYINPUT5), .B(n563), .ZN(n569) );
  NAND2_X1 U623 ( .A1(n797), .A2(G51), .ZN(n565) );
  NAND2_X1 U624 ( .A1(G63), .A2(n798), .ZN(n564) );
  NAND2_X1 U625 ( .A1(n565), .A2(n564), .ZN(n567) );
  XOR2_X1 U626 ( .A(KEYINPUT76), .B(KEYINPUT6), .Z(n566) );
  XNOR2_X1 U627 ( .A(n567), .B(n566), .ZN(n568) );
  NAND2_X1 U628 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U629 ( .A(KEYINPUT7), .B(n570), .ZN(G168) );
  NAND2_X1 U630 ( .A1(G88), .A2(n801), .ZN(n572) );
  NAND2_X1 U631 ( .A1(G50), .A2(n797), .ZN(n571) );
  NAND2_X1 U632 ( .A1(n572), .A2(n571), .ZN(n575) );
  NAND2_X1 U633 ( .A1(G75), .A2(n805), .ZN(n573) );
  XNOR2_X1 U634 ( .A(KEYINPUT83), .B(n573), .ZN(n574) );
  NOR2_X1 U635 ( .A1(n575), .A2(n574), .ZN(n577) );
  NAND2_X1 U636 ( .A1(G62), .A2(n798), .ZN(n576) );
  NAND2_X1 U637 ( .A1(n577), .A2(n576), .ZN(G303) );
  XOR2_X1 U638 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U639 ( .A1(G49), .A2(n797), .ZN(n579) );
  NAND2_X1 U640 ( .A1(G74), .A2(G651), .ZN(n578) );
  NAND2_X1 U641 ( .A1(n579), .A2(n578), .ZN(n580) );
  NOR2_X1 U642 ( .A1(n798), .A2(n580), .ZN(n581) );
  XNOR2_X1 U643 ( .A(n581), .B(KEYINPUT80), .ZN(n584) );
  NAND2_X1 U644 ( .A1(G87), .A2(n582), .ZN(n583) );
  NAND2_X1 U645 ( .A1(n584), .A2(n583), .ZN(G288) );
  NAND2_X1 U646 ( .A1(G48), .A2(n797), .ZN(n585) );
  XNOR2_X1 U647 ( .A(n585), .B(KEYINPUT82), .ZN(n593) );
  NAND2_X1 U648 ( .A1(n805), .A2(G73), .ZN(n586) );
  XNOR2_X1 U649 ( .A(n586), .B(KEYINPUT2), .ZN(n588) );
  NAND2_X1 U650 ( .A1(G61), .A2(n798), .ZN(n587) );
  NAND2_X1 U651 ( .A1(n588), .A2(n587), .ZN(n591) );
  NAND2_X1 U652 ( .A1(G86), .A2(n801), .ZN(n589) );
  XNOR2_X1 U653 ( .A(KEYINPUT81), .B(n589), .ZN(n590) );
  NOR2_X1 U654 ( .A1(n591), .A2(n590), .ZN(n592) );
  NAND2_X1 U655 ( .A1(n593), .A2(n592), .ZN(G305) );
  INV_X1 U656 ( .A(G303), .ZN(G166) );
  NAND2_X1 U657 ( .A1(n797), .A2(G47), .ZN(n595) );
  NAND2_X1 U658 ( .A1(G60), .A2(n798), .ZN(n594) );
  NAND2_X1 U659 ( .A1(n595), .A2(n594), .ZN(n598) );
  NAND2_X1 U660 ( .A1(n801), .A2(G85), .ZN(n596) );
  XOR2_X1 U661 ( .A(KEYINPUT64), .B(n596), .Z(n597) );
  NOR2_X1 U662 ( .A1(n598), .A2(n597), .ZN(n600) );
  NAND2_X1 U663 ( .A1(G72), .A2(n805), .ZN(n599) );
  NAND2_X1 U664 ( .A1(n600), .A2(n599), .ZN(G290) );
  NOR2_X1 U665 ( .A1(G164), .A2(G1384), .ZN(n719) );
  NAND2_X1 U666 ( .A1(G160), .A2(G40), .ZN(n718) );
  INV_X1 U667 ( .A(n718), .ZN(n601) );
  NAND2_X2 U668 ( .A1(n719), .A2(n601), .ZN(n674) );
  NAND2_X1 U669 ( .A1(G8), .A2(n674), .ZN(n717) );
  INV_X1 U670 ( .A(G1961), .ZN(n1000) );
  NAND2_X1 U671 ( .A1(n674), .A2(n1000), .ZN(n603) );
  INV_X1 U672 ( .A(n674), .ZN(n639) );
  XNOR2_X1 U673 ( .A(G2078), .B(KEYINPUT25), .ZN(n961) );
  NAND2_X1 U674 ( .A1(n639), .A2(n961), .ZN(n602) );
  NAND2_X1 U675 ( .A1(n603), .A2(n602), .ZN(n661) );
  NAND2_X1 U676 ( .A1(n661), .A2(G171), .ZN(n683) );
  NAND2_X1 U677 ( .A1(G66), .A2(n798), .ZN(n610) );
  NAND2_X1 U678 ( .A1(G92), .A2(n801), .ZN(n605) );
  NAND2_X1 U679 ( .A1(G54), .A2(n797), .ZN(n604) );
  NAND2_X1 U680 ( .A1(n605), .A2(n604), .ZN(n608) );
  NAND2_X1 U681 ( .A1(G79), .A2(n805), .ZN(n606) );
  XNOR2_X1 U682 ( .A(KEYINPUT75), .B(n606), .ZN(n607) );
  NOR2_X1 U683 ( .A1(n608), .A2(n607), .ZN(n609) );
  NAND2_X1 U684 ( .A1(n610), .A2(n609), .ZN(n611) );
  XOR2_X1 U685 ( .A(KEYINPUT15), .B(n611), .Z(n978) );
  NAND2_X1 U686 ( .A1(n798), .A2(G56), .ZN(n614) );
  INV_X1 U687 ( .A(KEYINPUT71), .ZN(n612) );
  AND2_X1 U688 ( .A1(G43), .A2(n797), .ZN(n622) );
  NAND2_X1 U689 ( .A1(G68), .A2(n805), .ZN(n618) );
  NAND2_X1 U690 ( .A1(G81), .A2(n801), .ZN(n615) );
  XNOR2_X1 U691 ( .A(n615), .B(KEYINPUT12), .ZN(n616) );
  XNOR2_X1 U692 ( .A(n616), .B(KEYINPUT72), .ZN(n617) );
  NAND2_X1 U693 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U694 ( .A(n619), .B(KEYINPUT73), .ZN(n620) );
  XNOR2_X1 U695 ( .A(KEYINPUT13), .B(n620), .ZN(n621) );
  NOR2_X1 U696 ( .A1(n622), .A2(n621), .ZN(n623) );
  INV_X1 U697 ( .A(KEYINPUT74), .ZN(n625) );
  NAND2_X1 U698 ( .A1(G1341), .A2(n674), .ZN(n627) );
  XOR2_X1 U699 ( .A(KEYINPUT96), .B(n627), .Z(n628) );
  NOR2_X1 U700 ( .A1(n981), .A2(n628), .ZN(n631) );
  NAND2_X1 U701 ( .A1(G1996), .A2(n639), .ZN(n629) );
  XNOR2_X1 U702 ( .A(KEYINPUT26), .B(n629), .ZN(n630) );
  NAND2_X1 U703 ( .A1(n631), .A2(n630), .ZN(n638) );
  NOR2_X1 U704 ( .A1(n978), .A2(n638), .ZN(n632) );
  XNOR2_X1 U705 ( .A(n632), .B(KEYINPUT97), .ZN(n636) );
  NOR2_X1 U706 ( .A1(G2067), .A2(n674), .ZN(n634) );
  NOR2_X1 U707 ( .A1(n639), .A2(G1348), .ZN(n633) );
  NOR2_X1 U708 ( .A1(n634), .A2(n633), .ZN(n635) );
  NAND2_X1 U709 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U710 ( .A(n637), .B(KEYINPUT98), .ZN(n648) );
  NAND2_X1 U711 ( .A1(n638), .A2(n978), .ZN(n646) );
  INV_X1 U712 ( .A(G299), .ZN(n809) );
  NAND2_X1 U713 ( .A1(n639), .A2(G2072), .ZN(n640) );
  XNOR2_X1 U714 ( .A(KEYINPUT27), .B(n640), .ZN(n643) );
  NAND2_X1 U715 ( .A1(G1956), .A2(n674), .ZN(n641) );
  XOR2_X1 U716 ( .A(KEYINPUT94), .B(n641), .Z(n642) );
  NOR2_X1 U717 ( .A1(n643), .A2(n642), .ZN(n650) );
  NOR2_X1 U718 ( .A1(n809), .A2(n650), .ZN(n645) );
  XNOR2_X1 U719 ( .A(KEYINPUT28), .B(KEYINPUT95), .ZN(n644) );
  XNOR2_X1 U720 ( .A(n645), .B(n644), .ZN(n649) );
  AND2_X1 U721 ( .A1(n646), .A2(n649), .ZN(n647) );
  NAND2_X1 U722 ( .A1(n648), .A2(n647), .ZN(n654) );
  INV_X1 U723 ( .A(n649), .ZN(n652) );
  NAND2_X1 U724 ( .A1(n809), .A2(n650), .ZN(n651) );
  OR2_X1 U725 ( .A1(n652), .A2(n651), .ZN(n653) );
  NAND2_X1 U726 ( .A1(n654), .A2(n653), .ZN(n656) );
  NAND2_X1 U727 ( .A1(n683), .A2(n523), .ZN(n665) );
  NOR2_X1 U728 ( .A1(G1966), .A2(n717), .ZN(n671) );
  NOR2_X1 U729 ( .A1(n674), .A2(G2084), .ZN(n657) );
  XNOR2_X1 U730 ( .A(n657), .B(KEYINPUT93), .ZN(n668) );
  NAND2_X1 U731 ( .A1(G8), .A2(n668), .ZN(n658) );
  NOR2_X1 U732 ( .A1(n671), .A2(n658), .ZN(n659) );
  XOR2_X1 U733 ( .A(KEYINPUT30), .B(n659), .Z(n660) );
  NOR2_X1 U734 ( .A1(G168), .A2(n660), .ZN(n663) );
  NOR2_X1 U735 ( .A1(G171), .A2(n661), .ZN(n662) );
  NOR2_X1 U736 ( .A1(n663), .A2(n662), .ZN(n664) );
  XOR2_X1 U737 ( .A(KEYINPUT31), .B(n664), .Z(n687) );
  NAND2_X1 U738 ( .A1(n665), .A2(n687), .ZN(n667) );
  INV_X1 U739 ( .A(KEYINPUT99), .ZN(n666) );
  XNOR2_X1 U740 ( .A(n667), .B(n666), .ZN(n673) );
  INV_X1 U741 ( .A(n668), .ZN(n669) );
  AND2_X1 U742 ( .A1(G8), .A2(n669), .ZN(n670) );
  NOR2_X1 U743 ( .A1(n671), .A2(n670), .ZN(n672) );
  NAND2_X1 U744 ( .A1(n673), .A2(n672), .ZN(n694) );
  INV_X1 U745 ( .A(G8), .ZN(n680) );
  NOR2_X1 U746 ( .A1(G1971), .A2(n717), .ZN(n676) );
  NOR2_X1 U747 ( .A1(G2090), .A2(n674), .ZN(n675) );
  NOR2_X1 U748 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U749 ( .A(n677), .B(KEYINPUT100), .ZN(n678) );
  NAND2_X1 U750 ( .A1(n678), .A2(G303), .ZN(n679) );
  OR2_X1 U751 ( .A1(n680), .A2(n679), .ZN(n686) );
  INV_X1 U752 ( .A(n686), .ZN(n682) );
  AND2_X1 U753 ( .A1(G286), .A2(G8), .ZN(n681) );
  OR2_X1 U754 ( .A1(n682), .A2(n681), .ZN(n685) );
  AND2_X1 U755 ( .A1(n683), .A2(n685), .ZN(n684) );
  NAND2_X1 U756 ( .A1(n523), .A2(n684), .ZN(n691) );
  INV_X1 U757 ( .A(n685), .ZN(n689) );
  AND2_X1 U758 ( .A1(n687), .A2(n686), .ZN(n688) );
  OR2_X1 U759 ( .A1(n689), .A2(n688), .ZN(n690) );
  AND2_X1 U760 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U761 ( .A(n692), .B(KEYINPUT32), .ZN(n693) );
  NAND2_X1 U762 ( .A1(n694), .A2(n693), .ZN(n709) );
  NOR2_X1 U763 ( .A1(G1976), .A2(G288), .ZN(n988) );
  NOR2_X1 U764 ( .A1(G1971), .A2(G303), .ZN(n695) );
  XOR2_X1 U765 ( .A(n695), .B(KEYINPUT101), .Z(n696) );
  NOR2_X1 U766 ( .A1(n988), .A2(n696), .ZN(n697) );
  XNOR2_X1 U767 ( .A(n697), .B(KEYINPUT102), .ZN(n698) );
  NAND2_X1 U768 ( .A1(n709), .A2(n698), .ZN(n699) );
  NAND2_X1 U769 ( .A1(G1976), .A2(G288), .ZN(n991) );
  NAND2_X1 U770 ( .A1(n699), .A2(n991), .ZN(n700) );
  NOR2_X1 U771 ( .A1(n717), .A2(n700), .ZN(n701) );
  NOR2_X1 U772 ( .A1(n701), .A2(KEYINPUT33), .ZN(n706) );
  NAND2_X1 U773 ( .A1(n988), .A2(KEYINPUT33), .ZN(n702) );
  NOR2_X1 U774 ( .A1(n702), .A2(n717), .ZN(n704) );
  XOR2_X1 U775 ( .A(G1981), .B(G305), .Z(n975) );
  NAND2_X1 U776 ( .A1(G8), .A2(G166), .ZN(n707) );
  NOR2_X1 U777 ( .A1(G2090), .A2(n707), .ZN(n708) );
  XNOR2_X1 U778 ( .A(n708), .B(KEYINPUT103), .ZN(n710) );
  NAND2_X1 U779 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U780 ( .A(n711), .B(KEYINPUT104), .ZN(n712) );
  NAND2_X1 U781 ( .A1(n712), .A2(n717), .ZN(n713) );
  NOR2_X1 U782 ( .A1(G1981), .A2(G305), .ZN(n715) );
  XOR2_X1 U783 ( .A(n715), .B(KEYINPUT24), .Z(n716) );
  NAND2_X1 U784 ( .A1(n526), .A2(n525), .ZN(n742) );
  XNOR2_X1 U785 ( .A(G1986), .B(G290), .ZN(n985) );
  NOR2_X1 U786 ( .A1(n719), .A2(n718), .ZN(n720) );
  XOR2_X1 U787 ( .A(KEYINPUT85), .B(n720), .Z(n767) );
  NAND2_X1 U788 ( .A1(n891), .A2(G117), .ZN(n721) );
  XNOR2_X1 U789 ( .A(n721), .B(KEYINPUT90), .ZN(n723) );
  NAND2_X1 U790 ( .A1(G129), .A2(n890), .ZN(n722) );
  NAND2_X1 U791 ( .A1(n723), .A2(n722), .ZN(n727) );
  NAND2_X1 U792 ( .A1(G105), .A2(n887), .ZN(n724) );
  XNOR2_X1 U793 ( .A(n724), .B(KEYINPUT38), .ZN(n725) );
  XNOR2_X1 U794 ( .A(n725), .B(KEYINPUT91), .ZN(n726) );
  NOR2_X1 U795 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U796 ( .A(n728), .B(KEYINPUT92), .ZN(n730) );
  NAND2_X1 U797 ( .A1(G141), .A2(n886), .ZN(n729) );
  NAND2_X1 U798 ( .A1(n730), .A2(n729), .ZN(n879) );
  NAND2_X1 U799 ( .A1(n879), .A2(G1996), .ZN(n740) );
  NAND2_X1 U800 ( .A1(G107), .A2(n891), .ZN(n731) );
  XOR2_X1 U801 ( .A(KEYINPUT88), .B(n731), .Z(n736) );
  NAND2_X1 U802 ( .A1(G131), .A2(n886), .ZN(n733) );
  NAND2_X1 U803 ( .A1(G95), .A2(n887), .ZN(n732) );
  NAND2_X1 U804 ( .A1(n733), .A2(n732), .ZN(n734) );
  XOR2_X1 U805 ( .A(KEYINPUT89), .B(n734), .Z(n735) );
  NOR2_X1 U806 ( .A1(n736), .A2(n735), .ZN(n738) );
  NAND2_X1 U807 ( .A1(n890), .A2(G119), .ZN(n737) );
  NAND2_X1 U808 ( .A1(n738), .A2(n737), .ZN(n897) );
  NAND2_X1 U809 ( .A1(n897), .A2(G1991), .ZN(n739) );
  AND2_X1 U810 ( .A1(n740), .A2(n739), .ZN(n935) );
  INV_X1 U811 ( .A(n767), .ZN(n741) );
  NOR2_X1 U812 ( .A1(n935), .A2(n741), .ZN(n745) );
  NAND2_X1 U813 ( .A1(n742), .A2(n521), .ZN(n765) );
  XOR2_X1 U814 ( .A(KEYINPUT105), .B(KEYINPUT39), .Z(n749) );
  NOR2_X1 U815 ( .A1(G1996), .A2(n879), .ZN(n942) );
  NOR2_X1 U816 ( .A1(G1986), .A2(G290), .ZN(n743) );
  NOR2_X1 U817 ( .A1(G1991), .A2(n897), .ZN(n930) );
  NOR2_X1 U818 ( .A1(n743), .A2(n930), .ZN(n744) );
  NOR2_X1 U819 ( .A1(n745), .A2(n744), .ZN(n746) );
  NOR2_X1 U820 ( .A1(n942), .A2(n746), .ZN(n747) );
  XNOR2_X1 U821 ( .A(n747), .B(KEYINPUT106), .ZN(n748) );
  XNOR2_X1 U822 ( .A(n749), .B(n748), .ZN(n750) );
  NAND2_X1 U823 ( .A1(n750), .A2(n767), .ZN(n763) );
  XOR2_X1 U824 ( .A(G2067), .B(KEYINPUT37), .Z(n766) );
  XNOR2_X1 U825 ( .A(KEYINPUT34), .B(KEYINPUT86), .ZN(n754) );
  NAND2_X1 U826 ( .A1(G140), .A2(n886), .ZN(n752) );
  NAND2_X1 U827 ( .A1(G104), .A2(n887), .ZN(n751) );
  NAND2_X1 U828 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U829 ( .A(n754), .B(n753), .ZN(n760) );
  NAND2_X1 U830 ( .A1(n890), .A2(G128), .ZN(n755) );
  XOR2_X1 U831 ( .A(KEYINPUT87), .B(n755), .Z(n757) );
  NAND2_X1 U832 ( .A1(n891), .A2(G116), .ZN(n756) );
  NAND2_X1 U833 ( .A1(n757), .A2(n756), .ZN(n758) );
  XOR2_X1 U834 ( .A(KEYINPUT35), .B(n758), .Z(n759) );
  NOR2_X1 U835 ( .A1(n760), .A2(n759), .ZN(n761) );
  XOR2_X1 U836 ( .A(KEYINPUT36), .B(n761), .Z(n900) );
  NOR2_X1 U837 ( .A1(n766), .A2(n900), .ZN(n947) );
  NAND2_X1 U838 ( .A1(n947), .A2(n767), .ZN(n762) );
  AND2_X1 U839 ( .A1(n763), .A2(n762), .ZN(n764) );
  NAND2_X1 U840 ( .A1(n765), .A2(n764), .ZN(n769) );
  AND2_X1 U841 ( .A1(n766), .A2(n900), .ZN(n933) );
  NAND2_X1 U842 ( .A1(n933), .A2(n767), .ZN(n768) );
  NAND2_X1 U843 ( .A1(n769), .A2(n768), .ZN(n770) );
  XNOR2_X1 U844 ( .A(n770), .B(n522), .ZN(G329) );
  AND2_X1 U845 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U846 ( .A(G57), .ZN(G237) );
  INV_X1 U847 ( .A(G132), .ZN(G219) );
  NAND2_X1 U848 ( .A1(G7), .A2(G661), .ZN(n771) );
  XNOR2_X1 U849 ( .A(n771), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U850 ( .A(KEYINPUT11), .B(KEYINPUT70), .Z(n773) );
  INV_X1 U851 ( .A(G223), .ZN(n835) );
  NAND2_X1 U852 ( .A1(G567), .A2(n835), .ZN(n772) );
  XNOR2_X1 U853 ( .A(n773), .B(n772), .ZN(G234) );
  INV_X1 U854 ( .A(G860), .ZN(n779) );
  OR2_X1 U855 ( .A1(n779), .A2(n981), .ZN(G153) );
  INV_X1 U856 ( .A(G171), .ZN(G301) );
  NAND2_X1 U857 ( .A1(G868), .A2(G301), .ZN(n775) );
  INV_X1 U858 ( .A(G868), .ZN(n819) );
  NAND2_X1 U859 ( .A1(n978), .A2(n819), .ZN(n774) );
  NAND2_X1 U860 ( .A1(n775), .A2(n774), .ZN(G284) );
  NAND2_X1 U861 ( .A1(n809), .A2(n819), .ZN(n776) );
  XNOR2_X1 U862 ( .A(n776), .B(KEYINPUT77), .ZN(n778) );
  NOR2_X1 U863 ( .A1(n819), .A2(G286), .ZN(n777) );
  NOR2_X1 U864 ( .A1(n778), .A2(n777), .ZN(G297) );
  NAND2_X1 U865 ( .A1(n779), .A2(G559), .ZN(n780) );
  INV_X1 U866 ( .A(n978), .ZN(n795) );
  NAND2_X1 U867 ( .A1(n780), .A2(n795), .ZN(n781) );
  XNOR2_X1 U868 ( .A(n781), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U869 ( .A1(n981), .A2(G868), .ZN(n784) );
  NAND2_X1 U870 ( .A1(G868), .A2(n795), .ZN(n782) );
  NOR2_X1 U871 ( .A1(G559), .A2(n782), .ZN(n783) );
  NOR2_X1 U872 ( .A1(n784), .A2(n783), .ZN(G282) );
  NAND2_X1 U873 ( .A1(G123), .A2(n890), .ZN(n785) );
  XNOR2_X1 U874 ( .A(n785), .B(KEYINPUT78), .ZN(n786) );
  XNOR2_X1 U875 ( .A(n786), .B(KEYINPUT18), .ZN(n788) );
  NAND2_X1 U876 ( .A1(G111), .A2(n891), .ZN(n787) );
  NAND2_X1 U877 ( .A1(n788), .A2(n787), .ZN(n792) );
  NAND2_X1 U878 ( .A1(G135), .A2(n886), .ZN(n790) );
  NAND2_X1 U879 ( .A1(G99), .A2(n887), .ZN(n789) );
  NAND2_X1 U880 ( .A1(n790), .A2(n789), .ZN(n791) );
  NOR2_X1 U881 ( .A1(n792), .A2(n791), .ZN(n929) );
  XNOR2_X1 U882 ( .A(n929), .B(G2096), .ZN(n794) );
  INV_X1 U883 ( .A(G2100), .ZN(n793) );
  NAND2_X1 U884 ( .A1(n794), .A2(n793), .ZN(G156) );
  NAND2_X1 U885 ( .A1(n795), .A2(G559), .ZN(n817) );
  XNOR2_X1 U886 ( .A(n981), .B(n817), .ZN(n796) );
  NOR2_X1 U887 ( .A1(G860), .A2(n796), .ZN(n808) );
  NAND2_X1 U888 ( .A1(n797), .A2(G55), .ZN(n800) );
  NAND2_X1 U889 ( .A1(G67), .A2(n798), .ZN(n799) );
  NAND2_X1 U890 ( .A1(n800), .A2(n799), .ZN(n804) );
  NAND2_X1 U891 ( .A1(G93), .A2(n801), .ZN(n802) );
  XNOR2_X1 U892 ( .A(KEYINPUT79), .B(n802), .ZN(n803) );
  NOR2_X1 U893 ( .A1(n804), .A2(n803), .ZN(n807) );
  NAND2_X1 U894 ( .A1(G80), .A2(n805), .ZN(n806) );
  NAND2_X1 U895 ( .A1(n807), .A2(n806), .ZN(n820) );
  XOR2_X1 U896 ( .A(n808), .B(n820), .Z(G145) );
  XNOR2_X1 U897 ( .A(G305), .B(G288), .ZN(n815) );
  XNOR2_X1 U898 ( .A(KEYINPUT84), .B(KEYINPUT19), .ZN(n811) );
  XNOR2_X1 U899 ( .A(G290), .B(n809), .ZN(n810) );
  XNOR2_X1 U900 ( .A(n811), .B(n810), .ZN(n812) );
  XNOR2_X1 U901 ( .A(G166), .B(n812), .ZN(n813) );
  XNOR2_X1 U902 ( .A(n813), .B(n820), .ZN(n814) );
  XNOR2_X1 U903 ( .A(n815), .B(n814), .ZN(n816) );
  XNOR2_X1 U904 ( .A(n981), .B(n816), .ZN(n904) );
  XOR2_X1 U905 ( .A(n904), .B(n817), .Z(n818) );
  NAND2_X1 U906 ( .A1(G868), .A2(n818), .ZN(n822) );
  NAND2_X1 U907 ( .A1(n820), .A2(n819), .ZN(n821) );
  NAND2_X1 U908 ( .A1(n822), .A2(n821), .ZN(G295) );
  NAND2_X1 U909 ( .A1(G2084), .A2(G2078), .ZN(n823) );
  XOR2_X1 U910 ( .A(KEYINPUT20), .B(n823), .Z(n824) );
  NAND2_X1 U911 ( .A1(G2090), .A2(n824), .ZN(n825) );
  XNOR2_X1 U912 ( .A(KEYINPUT21), .B(n825), .ZN(n826) );
  NAND2_X1 U913 ( .A1(n826), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U914 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U915 ( .A(KEYINPUT69), .B(G82), .ZN(G220) );
  NOR2_X1 U916 ( .A1(G219), .A2(G220), .ZN(n827) );
  XOR2_X1 U917 ( .A(KEYINPUT22), .B(n827), .Z(n828) );
  NOR2_X1 U918 ( .A1(G218), .A2(n828), .ZN(n829) );
  NAND2_X1 U919 ( .A1(G96), .A2(n829), .ZN(n922) );
  NAND2_X1 U920 ( .A1(n922), .A2(G2106), .ZN(n833) );
  NAND2_X1 U921 ( .A1(G120), .A2(G108), .ZN(n830) );
  NOR2_X1 U922 ( .A1(G237), .A2(n830), .ZN(n831) );
  NAND2_X1 U923 ( .A1(G69), .A2(n831), .ZN(n923) );
  NAND2_X1 U924 ( .A1(n923), .A2(G567), .ZN(n832) );
  NAND2_X1 U925 ( .A1(n833), .A2(n832), .ZN(n841) );
  NAND2_X1 U926 ( .A1(G483), .A2(G661), .ZN(n834) );
  NOR2_X1 U927 ( .A1(n841), .A2(n834), .ZN(n840) );
  NAND2_X1 U928 ( .A1(n840), .A2(G36), .ZN(G176) );
  NAND2_X1 U929 ( .A1(G2106), .A2(n835), .ZN(G217) );
  NAND2_X1 U930 ( .A1(G15), .A2(G2), .ZN(n836) );
  XNOR2_X1 U931 ( .A(KEYINPUT109), .B(n836), .ZN(n837) );
  NAND2_X1 U932 ( .A1(n837), .A2(G661), .ZN(n838) );
  XNOR2_X1 U933 ( .A(KEYINPUT110), .B(n838), .ZN(G259) );
  NAND2_X1 U934 ( .A1(G3), .A2(G1), .ZN(n839) );
  NAND2_X1 U935 ( .A1(n840), .A2(n839), .ZN(G188) );
  INV_X1 U936 ( .A(n841), .ZN(G319) );
  XOR2_X1 U937 ( .A(KEYINPUT42), .B(G2090), .Z(n843) );
  XNOR2_X1 U938 ( .A(G2078), .B(G2072), .ZN(n842) );
  XNOR2_X1 U939 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U940 ( .A(n844), .B(G2100), .Z(n846) );
  XNOR2_X1 U941 ( .A(G2084), .B(G2067), .ZN(n845) );
  XNOR2_X1 U942 ( .A(n846), .B(n845), .ZN(n850) );
  XOR2_X1 U943 ( .A(G2096), .B(KEYINPUT43), .Z(n848) );
  XNOR2_X1 U944 ( .A(KEYINPUT111), .B(G2678), .ZN(n847) );
  XNOR2_X1 U945 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U946 ( .A(n850), .B(n849), .Z(G227) );
  XOR2_X1 U947 ( .A(G1976), .B(G1981), .Z(n852) );
  XNOR2_X1 U948 ( .A(G1966), .B(G1971), .ZN(n851) );
  XNOR2_X1 U949 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U950 ( .A(n853), .B(KEYINPUT41), .Z(n855) );
  XNOR2_X1 U951 ( .A(G1961), .B(G1956), .ZN(n854) );
  XNOR2_X1 U952 ( .A(n855), .B(n854), .ZN(n859) );
  XOR2_X1 U953 ( .A(G2474), .B(G1986), .Z(n857) );
  XNOR2_X1 U954 ( .A(G1996), .B(G1991), .ZN(n856) );
  XNOR2_X1 U955 ( .A(n857), .B(n856), .ZN(n858) );
  XNOR2_X1 U956 ( .A(n859), .B(n858), .ZN(G229) );
  NAND2_X1 U957 ( .A1(G124), .A2(n890), .ZN(n860) );
  XNOR2_X1 U958 ( .A(n860), .B(KEYINPUT44), .ZN(n863) );
  NAND2_X1 U959 ( .A1(G100), .A2(n887), .ZN(n861) );
  XNOR2_X1 U960 ( .A(n861), .B(KEYINPUT112), .ZN(n862) );
  NAND2_X1 U961 ( .A1(n863), .A2(n862), .ZN(n867) );
  NAND2_X1 U962 ( .A1(G136), .A2(n886), .ZN(n865) );
  NAND2_X1 U963 ( .A1(G112), .A2(n891), .ZN(n864) );
  NAND2_X1 U964 ( .A1(n865), .A2(n864), .ZN(n866) );
  NOR2_X1 U965 ( .A1(n867), .A2(n866), .ZN(G162) );
  XOR2_X1 U966 ( .A(KEYINPUT48), .B(KEYINPUT115), .Z(n869) );
  XNOR2_X1 U967 ( .A(n929), .B(KEYINPUT46), .ZN(n868) );
  XNOR2_X1 U968 ( .A(n869), .B(n868), .ZN(n882) );
  NAND2_X1 U969 ( .A1(n890), .A2(G130), .ZN(n870) );
  XOR2_X1 U970 ( .A(KEYINPUT113), .B(n870), .Z(n872) );
  NAND2_X1 U971 ( .A1(n891), .A2(G118), .ZN(n871) );
  NAND2_X1 U972 ( .A1(n872), .A2(n871), .ZN(n873) );
  XNOR2_X1 U973 ( .A(KEYINPUT114), .B(n873), .ZN(n878) );
  NAND2_X1 U974 ( .A1(G142), .A2(n886), .ZN(n875) );
  NAND2_X1 U975 ( .A1(G106), .A2(n887), .ZN(n874) );
  NAND2_X1 U976 ( .A1(n875), .A2(n874), .ZN(n876) );
  XOR2_X1 U977 ( .A(n876), .B(KEYINPUT45), .Z(n877) );
  NOR2_X1 U978 ( .A1(n878), .A2(n877), .ZN(n880) );
  XNOR2_X1 U979 ( .A(n880), .B(n879), .ZN(n881) );
  XOR2_X1 U980 ( .A(n882), .B(n881), .Z(n884) );
  XNOR2_X1 U981 ( .A(G160), .B(G164), .ZN(n883) );
  XNOR2_X1 U982 ( .A(n884), .B(n883), .ZN(n885) );
  XNOR2_X1 U983 ( .A(G162), .B(n885), .ZN(n899) );
  NAND2_X1 U984 ( .A1(G139), .A2(n886), .ZN(n889) );
  NAND2_X1 U985 ( .A1(G103), .A2(n887), .ZN(n888) );
  NAND2_X1 U986 ( .A1(n889), .A2(n888), .ZN(n896) );
  NAND2_X1 U987 ( .A1(G127), .A2(n890), .ZN(n893) );
  NAND2_X1 U988 ( .A1(G115), .A2(n891), .ZN(n892) );
  NAND2_X1 U989 ( .A1(n893), .A2(n892), .ZN(n894) );
  XOR2_X1 U990 ( .A(KEYINPUT47), .B(n894), .Z(n895) );
  NOR2_X1 U991 ( .A1(n896), .A2(n895), .ZN(n925) );
  XNOR2_X1 U992 ( .A(n897), .B(n925), .ZN(n898) );
  XNOR2_X1 U993 ( .A(n899), .B(n898), .ZN(n901) );
  XNOR2_X1 U994 ( .A(n901), .B(n900), .ZN(n902) );
  NOR2_X1 U995 ( .A1(G37), .A2(n902), .ZN(G395) );
  XNOR2_X1 U996 ( .A(G286), .B(G301), .ZN(n903) );
  XNOR2_X1 U997 ( .A(n903), .B(n978), .ZN(n905) );
  XNOR2_X1 U998 ( .A(n905), .B(n904), .ZN(n906) );
  NOR2_X1 U999 ( .A1(G37), .A2(n906), .ZN(G397) );
  XOR2_X1 U1000 ( .A(KEYINPUT108), .B(G2446), .Z(n908) );
  XNOR2_X1 U1001 ( .A(G2443), .B(G2454), .ZN(n907) );
  XNOR2_X1 U1002 ( .A(n908), .B(n907), .ZN(n909) );
  XOR2_X1 U1003 ( .A(n909), .B(G2451), .Z(n911) );
  XNOR2_X1 U1004 ( .A(G1341), .B(G1348), .ZN(n910) );
  XNOR2_X1 U1005 ( .A(n911), .B(n910), .ZN(n915) );
  XOR2_X1 U1006 ( .A(G2435), .B(G2427), .Z(n913) );
  XNOR2_X1 U1007 ( .A(G2430), .B(G2438), .ZN(n912) );
  XNOR2_X1 U1008 ( .A(n913), .B(n912), .ZN(n914) );
  XOR2_X1 U1009 ( .A(n915), .B(n914), .Z(n916) );
  NAND2_X1 U1010 ( .A1(G14), .A2(n916), .ZN(n924) );
  NAND2_X1 U1011 ( .A1(G319), .A2(n924), .ZN(n919) );
  NOR2_X1 U1012 ( .A1(G227), .A2(G229), .ZN(n917) );
  XNOR2_X1 U1013 ( .A(KEYINPUT49), .B(n917), .ZN(n918) );
  NOR2_X1 U1014 ( .A1(n919), .A2(n918), .ZN(n921) );
  NOR2_X1 U1015 ( .A1(G395), .A2(G397), .ZN(n920) );
  NAND2_X1 U1016 ( .A1(n921), .A2(n920), .ZN(G225) );
  XOR2_X1 U1017 ( .A(KEYINPUT116), .B(G225), .Z(G308) );
  XNOR2_X1 U1018 ( .A(G108), .B(KEYINPUT117), .ZN(G238) );
  INV_X1 U1020 ( .A(G120), .ZN(G236) );
  INV_X1 U1021 ( .A(G96), .ZN(G221) );
  NOR2_X1 U1022 ( .A1(n923), .A2(n922), .ZN(G325) );
  INV_X1 U1023 ( .A(G325), .ZN(G261) );
  INV_X1 U1024 ( .A(G69), .ZN(G235) );
  INV_X1 U1025 ( .A(n924), .ZN(G401) );
  INV_X1 U1026 ( .A(KEYINPUT55), .ZN(n951) );
  XNOR2_X1 U1027 ( .A(KEYINPUT120), .B(KEYINPUT52), .ZN(n949) );
  XOR2_X1 U1028 ( .A(G2072), .B(n925), .Z(n927) );
  XOR2_X1 U1029 ( .A(G164), .B(G2078), .Z(n926) );
  NOR2_X1 U1030 ( .A1(n927), .A2(n926), .ZN(n928) );
  XOR2_X1 U1031 ( .A(KEYINPUT50), .B(n928), .Z(n940) );
  NOR2_X1 U1032 ( .A1(n930), .A2(n929), .ZN(n931) );
  XOR2_X1 U1033 ( .A(KEYINPUT118), .B(n931), .Z(n932) );
  NOR2_X1 U1034 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1035 ( .A1(n935), .A2(n934), .ZN(n937) );
  XOR2_X1 U1036 ( .A(G160), .B(G2084), .Z(n936) );
  NOR2_X1 U1037 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1038 ( .A(KEYINPUT119), .B(n938), .ZN(n939) );
  NOR2_X1 U1039 ( .A1(n940), .A2(n939), .ZN(n945) );
  XOR2_X1 U1040 ( .A(G2090), .B(G162), .Z(n941) );
  NOR2_X1 U1041 ( .A1(n942), .A2(n941), .ZN(n943) );
  XOR2_X1 U1042 ( .A(KEYINPUT51), .B(n943), .Z(n944) );
  NAND2_X1 U1043 ( .A1(n945), .A2(n944), .ZN(n946) );
  NOR2_X1 U1044 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1045 ( .A(n949), .B(n948), .ZN(n950) );
  NAND2_X1 U1046 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1047 ( .A1(n952), .A2(G29), .ZN(n1031) );
  XOR2_X1 U1048 ( .A(KEYINPUT55), .B(KEYINPUT122), .Z(n971) );
  XNOR2_X1 U1049 ( .A(G2090), .B(G35), .ZN(n966) );
  XNOR2_X1 U1050 ( .A(G1996), .B(G32), .ZN(n954) );
  XNOR2_X1 U1051 ( .A(G26), .B(G2067), .ZN(n953) );
  NOR2_X1 U1052 ( .A1(n954), .A2(n953), .ZN(n960) );
  XOR2_X1 U1053 ( .A(G2072), .B(G33), .Z(n955) );
  NAND2_X1 U1054 ( .A1(n955), .A2(G28), .ZN(n958) );
  XOR2_X1 U1055 ( .A(G25), .B(G1991), .Z(n956) );
  XNOR2_X1 U1056 ( .A(KEYINPUT121), .B(n956), .ZN(n957) );
  NOR2_X1 U1057 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1058 ( .A1(n960), .A2(n959), .ZN(n963) );
  XOR2_X1 U1059 ( .A(G27), .B(n961), .Z(n962) );
  NOR2_X1 U1060 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1061 ( .A(KEYINPUT53), .B(n964), .ZN(n965) );
  NOR2_X1 U1062 ( .A1(n966), .A2(n965), .ZN(n969) );
  XOR2_X1 U1063 ( .A(G2084), .B(G34), .Z(n967) );
  XNOR2_X1 U1064 ( .A(KEYINPUT54), .B(n967), .ZN(n968) );
  NAND2_X1 U1065 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1066 ( .A(n971), .B(n970), .ZN(n973) );
  INV_X1 U1067 ( .A(G29), .ZN(n972) );
  NAND2_X1 U1068 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1069 ( .A1(G11), .A2(n974), .ZN(n1029) );
  XNOR2_X1 U1070 ( .A(G16), .B(KEYINPUT56), .ZN(n999) );
  XNOR2_X1 U1071 ( .A(G1966), .B(G168), .ZN(n976) );
  NAND2_X1 U1072 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1073 ( .A(n977), .B(KEYINPUT57), .ZN(n997) );
  XNOR2_X1 U1074 ( .A(G299), .B(G1956), .ZN(n980) );
  XNOR2_X1 U1075 ( .A(n978), .B(G1348), .ZN(n979) );
  NOR2_X1 U1076 ( .A1(n980), .A2(n979), .ZN(n987) );
  XOR2_X1 U1077 ( .A(n981), .B(G1341), .Z(n983) );
  XNOR2_X1 U1078 ( .A(G171), .B(G1961), .ZN(n982) );
  NAND2_X1 U1079 ( .A1(n983), .A2(n982), .ZN(n984) );
  NOR2_X1 U1080 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1081 ( .A1(n987), .A2(n986), .ZN(n995) );
  XOR2_X1 U1082 ( .A(n988), .B(KEYINPUT123), .Z(n990) );
  XOR2_X1 U1083 ( .A(G166), .B(G1971), .Z(n989) );
  NOR2_X1 U1084 ( .A1(n990), .A2(n989), .ZN(n992) );
  NAND2_X1 U1085 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1086 ( .A(KEYINPUT124), .B(n993), .ZN(n994) );
  NOR2_X1 U1087 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1088 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1089 ( .A1(n999), .A2(n998), .ZN(n1027) );
  INV_X1 U1090 ( .A(G16), .ZN(n1025) );
  XNOR2_X1 U1091 ( .A(G5), .B(n1000), .ZN(n1015) );
  XNOR2_X1 U1092 ( .A(G1956), .B(G20), .ZN(n1005) );
  XNOR2_X1 U1093 ( .A(G1341), .B(G19), .ZN(n1002) );
  XNOR2_X1 U1094 ( .A(G1981), .B(G6), .ZN(n1001) );
  NOR2_X1 U1095 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1096 ( .A(KEYINPUT125), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1097 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1098 ( .A(KEYINPUT126), .B(n1006), .ZN(n1009) );
  XNOR2_X1 U1099 ( .A(G1348), .B(KEYINPUT59), .ZN(n1007) );
  XNOR2_X1 U1100 ( .A(n1007), .B(G4), .ZN(n1008) );
  NAND2_X1 U1101 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1102 ( .A(n1010), .B(KEYINPUT60), .ZN(n1011) );
  XOR2_X1 U1103 ( .A(KEYINPUT127), .B(n1011), .Z(n1013) );
  XNOR2_X1 U1104 ( .A(G1966), .B(G21), .ZN(n1012) );
  NOR2_X1 U1105 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1106 ( .A1(n1015), .A2(n1014), .ZN(n1022) );
  XNOR2_X1 U1107 ( .A(G1971), .B(G22), .ZN(n1017) );
  XNOR2_X1 U1108 ( .A(G23), .B(G1976), .ZN(n1016) );
  NOR2_X1 U1109 ( .A1(n1017), .A2(n1016), .ZN(n1019) );
  XOR2_X1 U1110 ( .A(G1986), .B(G24), .Z(n1018) );
  NAND2_X1 U1111 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1112 ( .A(KEYINPUT58), .B(n1020), .ZN(n1021) );
  NOR2_X1 U1113 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1114 ( .A(KEYINPUT61), .B(n1023), .ZN(n1024) );
  NAND2_X1 U1115 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1116 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NOR2_X1 U1117 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NAND2_X1 U1118 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XOR2_X1 U1119 ( .A(KEYINPUT62), .B(n1032), .Z(G311) );
  INV_X1 U1120 ( .A(G311), .ZN(G150) );
endmodule

