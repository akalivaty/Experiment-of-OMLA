//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 1 0 1 0 1 0 0 0 1 1 0 1 0 0 0 0 1 0 0 1 0 1 0 1 0 1 1 0 0 0 1 1 1 1 1 1 1 0 1 1 0 1 0 0 1 0 1 0 1 0 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:22 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n807, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n828, new_n829, new_n830, new_n831,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031;
  INV_X1    g000(.A(KEYINPUT89), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT9), .B(G234), .ZN(new_n188));
  OAI21_X1  g002(.A(G221), .B1(new_n188), .B2(G902), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G104), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(G107), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT85), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT3), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT3), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT85), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n192), .B1(new_n194), .B2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n191), .A2(G107), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n195), .A2(KEYINPUT85), .ZN(new_n199));
  INV_X1    g013(.A(G107), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G104), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n198), .B1(new_n199), .B2(new_n201), .ZN(new_n202));
  OAI21_X1  g016(.A(G101), .B1(new_n197), .B2(new_n202), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n200), .A2(G104), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n204), .B1(new_n192), .B2(new_n194), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n193), .A2(KEYINPUT3), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n201), .B1(new_n199), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G101), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n205), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n203), .A2(new_n209), .A3(KEYINPUT4), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT64), .ZN(new_n211));
  OR2_X1    g025(.A1(KEYINPUT0), .A2(G128), .ZN(new_n212));
  NAND2_X1  g026(.A1(KEYINPUT0), .A2(G128), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g028(.A(G143), .B(G146), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n211), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G146), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G143), .ZN(new_n218));
  INV_X1    g032(.A(G143), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G146), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n221), .A2(KEYINPUT64), .A3(new_n213), .A4(new_n212), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT65), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n223), .B1(new_n219), .B2(G146), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n217), .A2(KEYINPUT65), .A3(G143), .ZN(new_n225));
  INV_X1    g039(.A(new_n213), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n224), .A2(new_n225), .A3(new_n220), .A4(new_n226), .ZN(new_n227));
  AND3_X1   g041(.A1(new_n216), .A2(new_n222), .A3(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT4), .ZN(new_n229));
  OAI211_X1 g043(.A(new_n229), .B(G101), .C1(new_n197), .C2(new_n202), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n210), .A2(new_n228), .A3(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n224), .A2(new_n225), .A3(new_n220), .ZN(new_n232));
  OAI21_X1  g046(.A(KEYINPUT1), .B1(new_n219), .B2(G146), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G128), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(G128), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n236), .A2(KEYINPUT1), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n224), .A2(new_n225), .A3(new_n237), .A4(new_n220), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n235), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n201), .A2(new_n198), .A3(KEYINPUT86), .ZN(new_n240));
  OR3_X1    g054(.A1(new_n191), .A2(KEYINPUT86), .A3(G107), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n240), .A2(new_n241), .A3(G101), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n239), .A2(new_n209), .A3(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT10), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n234), .A2(new_n221), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(new_n238), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n247), .A2(new_n209), .A3(KEYINPUT10), .A4(new_n242), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT11), .ZN(new_n249));
  INV_X1    g063(.A(G134), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n249), .B1(new_n250), .B2(G137), .ZN(new_n251));
  INV_X1    g065(.A(G137), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n252), .A2(KEYINPUT11), .A3(G134), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n250), .A2(G137), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n251), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G131), .ZN(new_n256));
  AOI21_X1  g070(.A(G131), .B1(new_n250), .B2(G137), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n251), .A2(new_n257), .A3(new_n253), .ZN(new_n258));
  AND3_X1   g072(.A1(new_n256), .A2(KEYINPUT87), .A3(new_n258), .ZN(new_n259));
  AOI21_X1  g073(.A(KEYINPUT87), .B1(new_n256), .B2(new_n258), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n231), .A2(new_n245), .A3(new_n248), .A4(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n209), .A2(new_n242), .ZN(new_n263));
  AND4_X1   g077(.A1(new_n224), .A2(new_n225), .A3(new_n237), .A4(new_n220), .ZN(new_n264));
  AOI22_X1  g078(.A1(new_n233), .A2(G128), .B1(new_n218), .B2(new_n220), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(new_n243), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n256), .A2(new_n258), .ZN(new_n269));
  AOI21_X1  g083(.A(KEYINPUT12), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT12), .ZN(new_n271));
  AND2_X1   g085(.A1(new_n251), .A2(new_n253), .ZN(new_n272));
  AOI22_X1  g086(.A1(new_n272), .A2(new_n257), .B1(new_n255), .B2(G131), .ZN(new_n273));
  AOI211_X1 g087(.A(new_n271), .B(new_n273), .C1(new_n267), .C2(new_n243), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n262), .B1(new_n270), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G953), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(G227), .ZN(new_n277));
  XNOR2_X1  g091(.A(new_n277), .B(KEYINPUT84), .ZN(new_n278));
  XNOR2_X1  g092(.A(G110), .B(G140), .ZN(new_n279));
  XOR2_X1   g093(.A(new_n278), .B(new_n279), .Z(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  AND2_X1   g095(.A1(new_n262), .A2(new_n280), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n231), .A2(new_n245), .A3(new_n248), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(new_n269), .ZN(new_n284));
  AOI22_X1  g098(.A1(new_n275), .A2(new_n281), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(G469), .B1(new_n285), .B2(G902), .ZN(new_n286));
  INV_X1    g100(.A(G902), .ZN(new_n287));
  XOR2_X1   g101(.A(KEYINPUT88), .B(G469), .Z(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n270), .A2(new_n274), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n262), .A2(new_n280), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n280), .B1(new_n284), .B2(new_n262), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n287), .B(new_n289), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  AOI211_X1 g108(.A(new_n187), .B(new_n190), .C1(new_n286), .C2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n275), .A2(new_n281), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n282), .A2(new_n284), .ZN(new_n297));
  AOI21_X1  g111(.A(G902), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(G469), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n294), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(KEYINPUT89), .B1(new_n300), .B2(new_n189), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n295), .A2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(G237), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n303), .A2(new_n276), .A3(G214), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT92), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(G143), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  XNOR2_X1  g121(.A(KEYINPUT92), .B(G143), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n307), .B1(new_n308), .B2(new_n304), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n309), .A2(KEYINPUT17), .A3(G131), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(G131), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT17), .ZN(new_n312));
  INV_X1    g126(.A(new_n304), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n219), .A2(KEYINPUT92), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n306), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(G131), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n316), .A2(new_n317), .A3(new_n307), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n311), .A2(new_n312), .A3(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT16), .ZN(new_n320));
  INV_X1    g134(.A(G140), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n320), .A2(new_n321), .A3(G125), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(G125), .ZN(new_n323));
  INV_X1    g137(.A(G125), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G140), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  OAI211_X1 g140(.A(G146), .B(new_n322), .C1(new_n326), .C2(new_n320), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(KEYINPUT78), .ZN(new_n328));
  NOR3_X1   g142(.A1(new_n324), .A2(KEYINPUT16), .A3(G140), .ZN(new_n329));
  XNOR2_X1  g143(.A(G125), .B(G140), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n329), .B1(new_n330), .B2(KEYINPUT16), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n331), .A2(G146), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n328), .A2(new_n332), .ZN(new_n333));
  NOR3_X1   g147(.A1(new_n331), .A2(KEYINPUT78), .A3(G146), .ZN(new_n334));
  OAI211_X1 g148(.A(new_n310), .B(new_n319), .C1(new_n333), .C2(new_n334), .ZN(new_n335));
  XNOR2_X1  g149(.A(G113), .B(G122), .ZN(new_n336));
  XNOR2_X1  g150(.A(new_n336), .B(new_n191), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT94), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n307), .B(new_n338), .C1(new_n304), .C2(new_n308), .ZN(new_n339));
  NAND2_X1  g153(.A1(KEYINPUT18), .A2(G131), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n340), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n316), .A2(new_n338), .A3(new_n342), .A4(new_n307), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT95), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT80), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n326), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n330), .A2(KEYINPUT80), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n347), .A2(new_n348), .A3(new_n217), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n326), .A2(KEYINPUT93), .A3(G146), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT93), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n351), .B1(new_n330), .B2(new_n217), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n349), .A2(new_n350), .A3(new_n352), .ZN(new_n353));
  AND3_X1   g167(.A1(new_n344), .A2(new_n345), .A3(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n345), .B1(new_n344), .B2(new_n353), .ZN(new_n355));
  OAI211_X1 g169(.A(new_n335), .B(new_n337), .C1(new_n354), .C2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n311), .A2(new_n318), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT19), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n347), .A2(new_n348), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n326), .A2(KEYINPUT19), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n359), .A2(new_n217), .A3(new_n360), .ZN(new_n361));
  AND3_X1   g175(.A1(new_n357), .A2(new_n361), .A3(new_n327), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n344), .A2(new_n353), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(KEYINPUT95), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n344), .A2(new_n345), .A3(new_n353), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n362), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n356), .B1(new_n366), .B2(new_n337), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT20), .ZN(new_n368));
  NOR2_X1   g182(.A1(G475), .A2(G902), .ZN(new_n369));
  AND3_X1   g183(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT96), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n367), .A2(new_n371), .ZN(new_n372));
  OAI211_X1 g186(.A(new_n356), .B(KEYINPUT96), .C1(new_n366), .C2(new_n337), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n372), .A2(new_n369), .A3(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n370), .B1(new_n374), .B2(KEYINPUT20), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n335), .B1(new_n354), .B2(new_n355), .ZN(new_n376));
  INV_X1    g190(.A(new_n337), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(G902), .B1(new_n378), .B2(new_n356), .ZN(new_n379));
  INV_X1    g193(.A(G475), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n375), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n276), .A2(G952), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n383), .B1(G234), .B2(G237), .ZN(new_n384));
  INV_X1    g198(.A(G234), .ZN(new_n385));
  OAI211_X1 g199(.A(G902), .B(G953), .C1(new_n385), .C2(new_n303), .ZN(new_n386));
  XOR2_X1   g200(.A(new_n386), .B(KEYINPUT100), .Z(new_n387));
  XNOR2_X1  g201(.A(KEYINPUT21), .B(G898), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n384), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(G217), .ZN(new_n391));
  NOR3_X1   g205(.A1(new_n188), .A2(new_n391), .A3(G953), .ZN(new_n392));
  XNOR2_X1  g206(.A(new_n392), .B(KEYINPUT99), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(G122), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G116), .ZN(new_n396));
  INV_X1    g210(.A(G116), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(G122), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(G107), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n396), .A2(new_n398), .A3(new_n200), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n219), .A2(G128), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n236), .A2(G143), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n403), .A2(new_n404), .A3(new_n250), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT13), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n407), .B1(new_n236), .B2(G143), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n219), .A2(KEYINPUT13), .A3(G128), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n408), .A2(new_n404), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(G134), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT97), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n410), .A2(KEYINPUT97), .A3(G134), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n406), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n405), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n250), .B1(new_n403), .B2(new_n404), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n401), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT14), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n419), .A2(new_n397), .A3(G122), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n419), .B1(new_n397), .B2(G122), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(KEYINPUT98), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n421), .A2(KEYINPUT98), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n396), .B(new_n420), .C1(new_n423), .C2(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n418), .B1(new_n425), .B2(G107), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n394), .B1(new_n415), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n413), .A2(new_n414), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n428), .A2(new_n405), .A3(new_n402), .ZN(new_n429));
  OR2_X1    g243(.A1(new_n416), .A2(new_n417), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n420), .A2(new_n396), .ZN(new_n431));
  INV_X1    g245(.A(new_n424), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n431), .B1(new_n432), .B2(new_n422), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n401), .B(new_n430), .C1(new_n433), .C2(new_n200), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n429), .A2(new_n434), .A3(new_n393), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n427), .A2(new_n435), .A3(new_n287), .ZN(new_n436));
  INV_X1    g250(.A(G478), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n437), .A2(KEYINPUT15), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n436), .B(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n382), .A2(new_n390), .A3(new_n440), .ZN(new_n441));
  OAI21_X1  g255(.A(G214), .B1(G237), .B2(G902), .ZN(new_n442));
  AND3_X1   g256(.A1(KEYINPUT68), .A2(KEYINPUT2), .A3(G113), .ZN(new_n443));
  AOI21_X1  g257(.A(KEYINPUT68), .B1(KEYINPUT2), .B2(G113), .ZN(new_n444));
  OR2_X1    g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT70), .ZN(new_n446));
  OR2_X1    g260(.A1(KEYINPUT2), .A2(G113), .ZN(new_n447));
  XNOR2_X1  g261(.A(G116), .B(G119), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n445), .A2(new_n446), .A3(new_n447), .A4(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n447), .B1(new_n443), .B2(new_n444), .ZN(new_n450));
  XOR2_X1   g264(.A(G116), .B(G119), .Z(new_n451));
  OAI21_X1  g265(.A(KEYINPUT70), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n448), .A2(KEYINPUT5), .ZN(new_n453));
  NOR3_X1   g267(.A1(new_n397), .A2(KEYINPUT5), .A3(G119), .ZN(new_n454));
  INV_X1    g268(.A(G113), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  AOI22_X1  g270(.A1(new_n449), .A2(new_n452), .B1(new_n453), .B2(new_n456), .ZN(new_n457));
  NOR3_X1   g271(.A1(new_n197), .A2(new_n202), .A3(G101), .ZN(new_n458));
  AND3_X1   g272(.A1(new_n240), .A2(G101), .A3(new_n241), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n457), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n210), .A2(new_n230), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n445), .A2(KEYINPUT69), .A3(new_n447), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT69), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n448), .B1(new_n450), .B2(new_n464), .ZN(new_n465));
  AOI22_X1  g279(.A1(new_n449), .A2(new_n452), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n461), .B1(new_n462), .B2(new_n466), .ZN(new_n467));
  XNOR2_X1  g281(.A(G110), .B(G122), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  OAI211_X1 g284(.A(new_n461), .B(new_n468), .C1(new_n462), .C2(new_n466), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n470), .A2(KEYINPUT6), .A3(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT6), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n467), .A2(new_n473), .A3(new_n469), .ZN(new_n474));
  NOR3_X1   g288(.A1(new_n264), .A2(new_n265), .A3(G125), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n216), .A2(new_n222), .A3(new_n227), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n475), .B1(G125), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n276), .A2(G224), .ZN(new_n478));
  XNOR2_X1  g292(.A(new_n477), .B(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n472), .A2(new_n474), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n478), .A2(KEYINPUT7), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n477), .A2(new_n482), .ZN(new_n483));
  AND2_X1   g297(.A1(new_n471), .A2(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(KEYINPUT91), .B1(new_n477), .B2(new_n482), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n266), .A2(new_n324), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n486), .B1(new_n228), .B2(new_n324), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT91), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n487), .A2(new_n488), .A3(new_n481), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n449), .A2(new_n452), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n453), .A2(KEYINPUT90), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n453), .A2(KEYINPUT90), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(new_n456), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n490), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(new_n460), .ZN(new_n495));
  XOR2_X1   g309(.A(new_n468), .B(KEYINPUT8), .Z(new_n496));
  AOI21_X1  g310(.A(new_n496), .B1(new_n457), .B2(new_n263), .ZN(new_n497));
  AOI22_X1  g311(.A1(new_n485), .A2(new_n489), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(G902), .B1(new_n484), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(G210), .B1(G237), .B2(G902), .ZN(new_n500));
  AND3_X1   g314(.A1(new_n480), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n500), .B1(new_n480), .B2(new_n499), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n442), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NOR3_X1   g317(.A1(new_n302), .A2(new_n441), .A3(new_n503), .ZN(new_n504));
  XNOR2_X1  g318(.A(KEYINPUT26), .B(G101), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n303), .A2(new_n276), .A3(G210), .ZN(new_n506));
  OR2_X1    g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n505), .A2(new_n506), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g323(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n507), .A2(new_n510), .A3(new_n508), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  XOR2_X1   g328(.A(KEYINPUT73), .B(KEYINPUT28), .Z(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n269), .A2(new_n227), .A3(new_n216), .A4(new_n222), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT66), .ZN(new_n518));
  AND3_X1   g332(.A1(new_n251), .A2(new_n257), .A3(new_n253), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n252), .A2(G134), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n317), .B1(new_n520), .B2(new_n254), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n518), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n521), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n523), .A2(KEYINPUT66), .A3(new_n258), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n522), .A2(new_n247), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n517), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n463), .A2(new_n465), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n490), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n247), .A2(new_n258), .A3(new_n523), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n466), .A2(new_n517), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n516), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n523), .A2(new_n258), .ZN(new_n534));
  OAI22_X1  g348(.A1(new_n476), .A2(new_n273), .B1(new_n266), .B2(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n528), .B1(new_n535), .B2(KEYINPUT74), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT74), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n517), .A2(new_n537), .A3(new_n530), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT28), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n514), .B1(new_n533), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT31), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n517), .A2(KEYINPUT30), .A3(new_n530), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(new_n528), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT30), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n526), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT67), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n526), .A2(KEYINPUT67), .A3(new_n546), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n545), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  OAI211_X1 g365(.A(KEYINPUT72), .B(new_n514), .C1(new_n535), .C2(new_n528), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(KEYINPUT72), .B1(new_n531), .B2(new_n514), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n543), .B1(new_n551), .B2(new_n555), .ZN(new_n556));
  AND2_X1   g370(.A1(new_n544), .A2(new_n528), .ZN(new_n557));
  AOI21_X1  g371(.A(KEYINPUT67), .B1(new_n526), .B2(new_n546), .ZN(new_n558));
  AOI211_X1 g372(.A(new_n548), .B(KEYINPUT30), .C1(new_n517), .C2(new_n525), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n514), .B1(new_n535), .B2(new_n528), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT72), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(new_n552), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n560), .A2(KEYINPUT31), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n542), .B1(new_n556), .B2(new_n565), .ZN(new_n566));
  NOR2_X1   g380(.A1(G472), .A2(G902), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NOR3_X1   g382(.A1(new_n566), .A2(KEYINPUT32), .A3(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT32), .ZN(new_n570));
  INV_X1    g384(.A(new_n514), .ZN(new_n571));
  AOI21_X1  g385(.A(KEYINPUT28), .B1(new_n536), .B2(new_n538), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n571), .B1(new_n532), .B2(new_n572), .ZN(new_n573));
  AND3_X1   g387(.A1(new_n560), .A2(KEYINPUT31), .A3(new_n564), .ZN(new_n574));
  AOI21_X1  g388(.A(KEYINPUT31), .B1(new_n560), .B2(new_n564), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n570), .B1(new_n576), .B2(new_n567), .ZN(new_n577));
  INV_X1    g391(.A(G472), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n535), .B(new_n466), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n541), .B1(new_n579), .B2(new_n540), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n514), .A2(KEYINPUT29), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n287), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n533), .A2(new_n541), .A3(new_n514), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n514), .B1(new_n560), .B2(new_n531), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n583), .B1(new_n584), .B2(KEYINPUT75), .ZN(new_n585));
  NOR3_X1   g399(.A1(new_n532), .A2(new_n572), .A3(new_n571), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT75), .ZN(new_n587));
  AOI21_X1  g401(.A(KEYINPUT29), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n582), .B1(new_n585), .B2(new_n588), .ZN(new_n589));
  OAI22_X1  g403(.A1(new_n569), .A2(new_n577), .B1(new_n578), .B2(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(KEYINPUT22), .B(G137), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n276), .A2(G221), .A3(G234), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n591), .B(new_n592), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n322), .B1(new_n326), .B2(new_n320), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(new_n217), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n595), .A2(KEYINPUT78), .A3(new_n327), .ZN(new_n596));
  OR3_X1    g410(.A1(new_n331), .A2(KEYINPUT78), .A3(G146), .ZN(new_n597));
  INV_X1    g411(.A(G119), .ZN(new_n598));
  OAI21_X1  g412(.A(KEYINPUT77), .B1(new_n598), .B2(G128), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT77), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n600), .A2(new_n236), .A3(G119), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n598), .A2(G128), .ZN(new_n602));
  AND3_X1   g416(.A1(new_n599), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  XOR2_X1   g417(.A(KEYINPUT24), .B(G110), .Z(new_n604));
  NAND3_X1  g418(.A1(new_n236), .A2(KEYINPUT23), .A3(G119), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n598), .A2(G128), .ZN(new_n606));
  OAI211_X1 g420(.A(new_n602), .B(new_n605), .C1(new_n606), .C2(KEYINPUT23), .ZN(new_n607));
  AOI22_X1  g421(.A1(new_n603), .A2(new_n604), .B1(new_n607), .B2(G110), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n596), .A2(new_n597), .A3(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(KEYINPUT79), .B(G110), .ZN(new_n610));
  OAI22_X1  g424(.A1(new_n603), .A2(new_n604), .B1(new_n607), .B2(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n611), .A2(new_n349), .A3(new_n327), .ZN(new_n612));
  AND3_X1   g426(.A1(new_n609), .A2(KEYINPUT81), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(KEYINPUT81), .B1(new_n609), .B2(new_n612), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n593), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT25), .ZN(new_n616));
  INV_X1    g430(.A(new_n593), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n609), .A2(new_n612), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT81), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n615), .A2(new_n616), .A3(new_n287), .A4(new_n620), .ZN(new_n621));
  OAI21_X1  g435(.A(G217), .B1(new_n385), .B2(G902), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(KEYINPUT76), .ZN(new_n623));
  AND2_X1   g437(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  XOR2_X1   g438(.A(KEYINPUT82), .B(KEYINPUT25), .Z(new_n625));
  NAND2_X1  g439(.A1(new_n615), .A2(new_n620), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n625), .B1(new_n626), .B2(G902), .ZN(new_n627));
  INV_X1    g441(.A(new_n626), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n622), .A2(new_n287), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  AOI22_X1  g444(.A1(new_n624), .A2(new_n627), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n590), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n632), .A2(KEYINPUT83), .ZN(new_n633));
  INV_X1    g447(.A(new_n631), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n585), .A2(new_n588), .ZN(new_n635));
  INV_X1    g449(.A(new_n582), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(G472), .ZN(new_n638));
  OAI21_X1  g452(.A(KEYINPUT32), .B1(new_n566), .B2(new_n568), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n576), .A2(new_n570), .A3(new_n567), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n634), .B1(new_n638), .B2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT83), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n504), .B1(new_n633), .B2(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(G101), .ZN(G3));
  AND3_X1   g460(.A1(new_n239), .A2(new_n209), .A3(new_n242), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n247), .B1(new_n209), .B2(new_n242), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n269), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n271), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n268), .A2(KEYINPUT12), .A3(new_n269), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n280), .B1(new_n652), .B2(new_n262), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n458), .A2(new_n244), .A3(new_n459), .ZN(new_n654));
  AOI22_X1  g468(.A1(new_n654), .A2(new_n247), .B1(new_n243), .B2(new_n244), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n273), .B1(new_n655), .B2(new_n231), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n291), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n287), .B1(new_n653), .B2(new_n657), .ZN(new_n658));
  AND4_X1   g472(.A1(new_n231), .A2(new_n245), .A3(new_n248), .A4(new_n261), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n281), .B1(new_n656), .B2(new_n659), .ZN(new_n660));
  OAI211_X1 g474(.A(new_n262), .B(new_n280), .C1(new_n270), .C2(new_n274), .ZN(new_n661));
  AOI21_X1  g475(.A(G902), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  AOI22_X1  g476(.A1(new_n658), .A2(G469), .B1(new_n662), .B2(new_n289), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n187), .B1(new_n663), .B2(new_n190), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n300), .A2(KEYINPUT89), .A3(new_n189), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n578), .B1(new_n576), .B2(new_n287), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n667), .B1(new_n567), .B2(new_n576), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n666), .A2(new_n668), .A3(new_n631), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(KEYINPUT101), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT101), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n666), .A2(new_n668), .A3(new_n671), .A4(new_n631), .ZN(new_n672));
  AND2_X1   g486(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  AND2_X1   g487(.A1(new_n427), .A2(new_n435), .ZN(new_n674));
  AND3_X1   g488(.A1(new_n674), .A2(KEYINPUT102), .A3(KEYINPUT33), .ZN(new_n675));
  AOI21_X1  g489(.A(KEYINPUT33), .B1(new_n674), .B2(KEYINPUT102), .ZN(new_n676));
  OAI211_X1 g490(.A(G478), .B(new_n287), .C1(new_n675), .C2(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n436), .A2(new_n437), .ZN(new_n678));
  AND2_X1   g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n374), .A2(KEYINPUT20), .ZN(new_n680));
  INV_X1    g494(.A(new_n370), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n381), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n679), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  OAI211_X1 g498(.A(new_n390), .B(new_n442), .C1(new_n501), .C2(new_n502), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  AOI21_X1  g500(.A(KEYINPUT103), .B1(new_n684), .B2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT103), .ZN(new_n688));
  NOR4_X1   g502(.A1(new_n382), .A2(new_n685), .A3(new_n679), .A4(new_n688), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n673), .B1(new_n687), .B2(new_n689), .ZN(new_n690));
  XOR2_X1   g504(.A(KEYINPUT34), .B(G104), .Z(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(G6));
  NAND4_X1  g506(.A1(new_n372), .A2(new_n368), .A3(new_n369), .A4(new_n373), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n680), .A2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n436), .B(new_n438), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n696), .B1(new_n379), .B2(new_n380), .ZN(new_n697));
  NOR3_X1   g511(.A1(new_n695), .A2(new_n685), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n673), .A2(new_n698), .ZN(new_n699));
  XOR2_X1   g513(.A(KEYINPUT35), .B(G107), .Z(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(G9));
  NOR2_X1   g515(.A1(new_n617), .A2(KEYINPUT36), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(KEYINPUT104), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(new_n618), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n630), .ZN(new_n705));
  INV_X1    g519(.A(new_n627), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n621), .A2(new_n623), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n705), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  AND2_X1   g522(.A1(new_n668), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n504), .A2(new_n709), .ZN(new_n710));
  XOR2_X1   g524(.A(KEYINPUT37), .B(G110), .Z(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(KEYINPUT105), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n710), .B(new_n712), .ZN(G12));
  AOI22_X1  g527(.A1(new_n624), .A2(new_n627), .B1(new_n630), .B2(new_n704), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n503), .A2(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(G900), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n384), .B1(new_n387), .B2(new_n716), .ZN(new_n717));
  AOI211_X1 g531(.A(new_n717), .B(new_n697), .C1(new_n680), .C2(new_n693), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n666), .A2(new_n590), .A3(new_n715), .A4(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G128), .ZN(G30));
  XOR2_X1   g534(.A(new_n717), .B(KEYINPUT39), .Z(new_n721));
  NAND2_X1  g535(.A1(new_n666), .A2(new_n721), .ZN(new_n722));
  OR2_X1    g536(.A1(new_n722), .A2(KEYINPUT40), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n440), .B1(new_n682), .B2(new_n683), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n724), .A2(new_n442), .A3(new_n714), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n551), .A2(new_n555), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n579), .A2(new_n514), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  OAI21_X1  g542(.A(G472), .B1(new_n728), .B2(G902), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n729), .B1(new_n569), .B2(new_n577), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n501), .A2(new_n502), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(KEYINPUT38), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n725), .A2(new_n731), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n722), .A2(KEYINPUT40), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n723), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G143), .ZN(G45));
  NAND2_X1  g551(.A1(new_n677), .A2(new_n678), .ZN(new_n738));
  INV_X1    g552(.A(new_n717), .ZN(new_n739));
  OAI211_X1 g553(.A(new_n738), .B(new_n739), .C1(new_n375), .C2(new_n381), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n741), .A2(new_n666), .A3(new_n590), .A4(new_n715), .ZN(new_n742));
  XNOR2_X1  g556(.A(KEYINPUT106), .B(G146), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n742), .B(new_n743), .ZN(G48));
  OAI21_X1  g558(.A(new_n287), .B1(new_n292), .B2(new_n293), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(KEYINPUT107), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT107), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n662), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n746), .A2(G469), .A3(new_n748), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n190), .B1(new_n662), .B2(new_n289), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n749), .A2(new_n631), .A3(new_n750), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n751), .B1(new_n638), .B2(new_n641), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n752), .B1(new_n687), .B2(new_n689), .ZN(new_n753));
  XNOR2_X1  g567(.A(KEYINPUT41), .B(G113), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n753), .B(new_n754), .ZN(G15));
  NAND2_X1  g569(.A1(new_n752), .A2(new_n698), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G116), .ZN(G18));
  NOR2_X1   g571(.A1(new_n441), .A2(new_n714), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT108), .ZN(new_n759));
  OAI21_X1  g573(.A(G469), .B1(new_n662), .B2(new_n747), .ZN(new_n760));
  AOI211_X1 g574(.A(KEYINPUT107), .B(G902), .C1(new_n660), .C2(new_n661), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n750), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n759), .B1(new_n762), .B2(new_n503), .ZN(new_n763));
  INV_X1    g577(.A(new_n442), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n480), .A2(new_n499), .ZN(new_n765));
  INV_X1    g579(.A(new_n500), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n480), .A2(new_n499), .A3(new_n500), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n764), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n769), .A2(KEYINPUT108), .A3(new_n749), .A4(new_n750), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n763), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n758), .A2(new_n590), .A3(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(KEYINPUT109), .B(G119), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n772), .B(new_n773), .ZN(G21));
  OAI21_X1  g588(.A(new_n696), .B1(new_n375), .B2(new_n381), .ZN(new_n775));
  OAI211_X1 g589(.A(new_n390), .B(new_n750), .C1(new_n760), .C2(new_n761), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n775), .A2(new_n503), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n556), .A2(new_n565), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n580), .A2(new_n571), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n568), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NOR3_X1   g594(.A1(new_n634), .A2(new_n667), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n777), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G122), .ZN(G24));
  OAI21_X1  g597(.A(G472), .B1(new_n566), .B2(G902), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n779), .B1(new_n574), .B2(new_n575), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n567), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n784), .A2(new_n708), .A3(new_n786), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n787), .A2(new_n740), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n771), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G125), .ZN(G27));
  NAND2_X1  g604(.A1(G469), .A2(G902), .ZN(new_n791));
  XOR2_X1   g605(.A(new_n791), .B(KEYINPUT110), .Z(new_n792));
  NAND2_X1  g606(.A1(new_n296), .A2(new_n297), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n792), .B1(new_n793), .B2(new_n299), .ZN(new_n794));
  AOI211_X1 g608(.A(G902), .B(new_n288), .C1(new_n660), .C2(new_n661), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n189), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n767), .A2(new_n442), .A3(new_n768), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n741), .A2(new_n590), .A3(new_n631), .A4(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT42), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n642), .A2(KEYINPUT42), .A3(new_n741), .A4(new_n798), .ZN(new_n802));
  AND3_X1   g616(.A1(new_n801), .A2(KEYINPUT111), .A3(new_n802), .ZN(new_n803));
  AOI21_X1  g617(.A(KEYINPUT111), .B1(new_n801), .B2(new_n802), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G131), .ZN(G33));
  NAND4_X1  g620(.A1(new_n590), .A2(new_n631), .A3(new_n718), .A4(new_n798), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(G134), .ZN(G36));
  NAND2_X1  g622(.A1(new_n382), .A2(new_n738), .ZN(new_n809));
  XOR2_X1   g623(.A(new_n809), .B(KEYINPUT43), .Z(new_n810));
  NOR2_X1   g624(.A1(new_n668), .A2(new_n714), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  OR2_X1    g626(.A1(new_n812), .A2(KEYINPUT44), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(KEYINPUT44), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT45), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n299), .B1(new_n793), .B2(new_n815), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n816), .B1(new_n815), .B2(new_n793), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(new_n792), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT46), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n795), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n820), .B1(new_n819), .B2(new_n818), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(new_n189), .ZN(new_n822));
  INV_X1    g636(.A(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(new_n721), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n824), .A2(new_n797), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n813), .A2(new_n814), .A3(new_n825), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(G137), .ZN(G39));
  INV_X1    g641(.A(KEYINPUT47), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n822), .B(new_n828), .ZN(new_n829));
  NOR4_X1   g643(.A1(new_n590), .A2(new_n740), .A3(new_n631), .A4(new_n797), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(new_n321), .ZN(G42));
  NOR4_X1   g646(.A1(new_n809), .A2(new_n190), .A3(new_n764), .A4(new_n634), .ZN(new_n833));
  XOR2_X1   g647(.A(new_n833), .B(KEYINPUT112), .Z(new_n834));
  NAND2_X1  g648(.A1(new_n749), .A2(new_n294), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n733), .B1(KEYINPUT49), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n836), .B1(KEYINPUT49), .B2(new_n835), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n834), .A2(new_n731), .A3(new_n837), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n810), .A2(new_n384), .ZN(new_n839));
  AND4_X1   g653(.A1(new_n764), .A2(new_n733), .A3(new_n749), .A4(new_n750), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n839), .A2(new_n781), .A3(new_n840), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n841), .B(KEYINPUT50), .ZN(new_n842));
  INV_X1    g656(.A(new_n829), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n843), .B1(new_n189), .B2(new_n835), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n501), .A2(new_n502), .A3(new_n764), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n844), .A2(new_n781), .A3(new_n845), .A4(new_n839), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n762), .A2(new_n797), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n839), .A2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(new_n848), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n667), .A2(new_n714), .A3(new_n780), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  AND4_X1   g665(.A1(new_n384), .A2(new_n731), .A3(new_n631), .A4(new_n847), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n852), .A2(new_n382), .A3(new_n679), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n842), .A2(new_n846), .A3(new_n851), .A4(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT51), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n839), .A2(new_n771), .A3(new_n781), .ZN(new_n857));
  XOR2_X1   g671(.A(new_n383), .B(KEYINPUT115), .Z(new_n858));
  AOI21_X1  g672(.A(new_n858), .B1(new_n852), .B2(new_n684), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(KEYINPUT116), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n848), .A2(new_n632), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n862), .B(KEYINPUT48), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n860), .A2(KEYINPUT116), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n856), .A2(new_n861), .A3(new_n865), .ZN(new_n866));
  OAI211_X1 g680(.A(new_n189), .B(new_n739), .C1(new_n794), .C2(new_n795), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n867), .A2(new_n708), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n730), .A2(new_n868), .A3(new_n724), .A4(new_n769), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n789), .A2(new_n742), .A3(new_n719), .A4(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(KEYINPUT52), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n769), .A2(new_n708), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n872), .B1(new_n638), .B2(new_n641), .ZN(new_n873));
  OAI211_X1 g687(.A(new_n873), .B(new_n666), .C1(new_n718), .C2(new_n741), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT52), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n874), .A2(new_n875), .A3(new_n789), .A4(new_n869), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n871), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n741), .A2(new_n850), .A3(new_n798), .ZN(new_n878));
  AND2_X1   g692(.A1(new_n807), .A2(new_n878), .ZN(new_n879));
  OAI211_X1 g693(.A(new_n440), .B(new_n739), .C1(new_n379), .C2(new_n380), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n880), .B1(new_n680), .B2(new_n693), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n881), .A2(new_n708), .A3(new_n845), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n302), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(KEYINPUT113), .B1(new_n883), .B2(new_n590), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n881), .A2(new_n708), .A3(new_n845), .ZN(new_n885));
  AND4_X1   g699(.A1(KEYINPUT113), .A2(new_n885), .A3(new_n666), .A4(new_n590), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n879), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  AOI22_X1  g701(.A1(new_n752), .A2(new_n698), .B1(new_n777), .B2(new_n781), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n888), .A2(new_n753), .A3(new_n772), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n382), .A2(new_n440), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n679), .B1(new_n375), .B2(new_n381), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n893), .A2(new_n685), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n670), .A2(new_n894), .A3(new_n672), .ZN(new_n895));
  AND3_X1   g709(.A1(new_n645), .A2(new_n710), .A3(new_n895), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n877), .A2(new_n805), .A3(new_n890), .A4(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT53), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n897), .B(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(KEYINPUT54), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n897), .A2(new_n898), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT54), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n807), .A2(new_n878), .ZN(new_n903));
  INV_X1    g717(.A(new_n886), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n885), .A2(new_n666), .A3(new_n590), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT113), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n903), .B1(new_n904), .B2(new_n907), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n642), .B(new_n643), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n504), .B1(new_n909), .B2(new_n709), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT114), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n908), .A2(new_n910), .A3(new_n911), .A4(new_n895), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n645), .A2(new_n895), .A3(new_n710), .ZN(new_n913));
  OAI21_X1  g727(.A(KEYINPUT114), .B1(new_n913), .B2(new_n887), .ZN(new_n914));
  AND2_X1   g728(.A1(new_n801), .A2(new_n802), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n915), .A2(new_n889), .A3(new_n898), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n912), .A2(new_n914), .A3(new_n877), .A4(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n901), .A2(new_n902), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n900), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n854), .A2(new_n855), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n866), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  NOR2_X1   g735(.A1(G952), .A2(G953), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n838), .B1(new_n921), .B2(new_n922), .ZN(G75));
  NOR2_X1   g737(.A1(new_n276), .A2(G952), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n287), .B1(new_n901), .B2(new_n917), .ZN(new_n925));
  AOI21_X1  g739(.A(KEYINPUT56), .B1(new_n925), .B2(G210), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n472), .A2(new_n474), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(new_n479), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT55), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n926), .A2(new_n929), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n926), .A2(new_n929), .ZN(new_n931));
  OR2_X1    g745(.A1(new_n931), .A2(KEYINPUT117), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(KEYINPUT117), .ZN(new_n933));
  AOI211_X1 g747(.A(new_n924), .B(new_n930), .C1(new_n932), .C2(new_n933), .ZN(G51));
  AOI211_X1 g748(.A(new_n287), .B(new_n817), .C1(new_n901), .C2(new_n917), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n292), .A2(new_n293), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n792), .B(KEYINPUT57), .Z(new_n937));
  AND3_X1   g751(.A1(new_n901), .A2(new_n902), .A3(new_n917), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n902), .B1(new_n901), .B2(new_n917), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n937), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(KEYINPUT118), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT118), .ZN(new_n942));
  OAI211_X1 g756(.A(new_n942), .B(new_n937), .C1(new_n938), .C2(new_n939), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n936), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT119), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n935), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(new_n936), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n901), .A2(new_n917), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n948), .A2(KEYINPUT54), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(new_n918), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n942), .B1(new_n950), .B2(new_n937), .ZN(new_n951));
  INV_X1    g765(.A(new_n943), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n947), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(KEYINPUT119), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n924), .B1(new_n946), .B2(new_n954), .ZN(G54));
  NAND3_X1  g769(.A1(new_n925), .A2(KEYINPUT58), .A3(G475), .ZN(new_n956));
  AND2_X1   g770(.A1(new_n372), .A2(new_n373), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  AND3_X1   g772(.A1(new_n956), .A2(KEYINPUT120), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(KEYINPUT120), .B1(new_n956), .B2(new_n958), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n956), .A2(new_n958), .ZN(new_n961));
  NOR4_X1   g775(.A1(new_n959), .A2(new_n960), .A3(new_n961), .A4(new_n924), .ZN(G60));
  OR2_X1    g776(.A1(new_n675), .A2(new_n676), .ZN(new_n963));
  NAND2_X1  g777(.A1(G478), .A2(G902), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(KEYINPUT122), .ZN(new_n965));
  XNOR2_X1  g779(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n965), .B(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n963), .B1(new_n919), .B2(new_n968), .ZN(new_n969));
  AND3_X1   g783(.A1(new_n950), .A2(new_n963), .A3(new_n968), .ZN(new_n970));
  NOR3_X1   g784(.A1(new_n969), .A2(new_n970), .A3(new_n924), .ZN(G63));
  NAND2_X1  g785(.A1(G217), .A2(G902), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n972), .B(KEYINPUT60), .Z(new_n973));
  NAND2_X1  g787(.A1(new_n948), .A2(new_n973), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n626), .B(KEYINPUT124), .Z(new_n975));
  AOI21_X1  g789(.A(new_n924), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(new_n974), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT123), .ZN(new_n978));
  AND3_X1   g792(.A1(new_n977), .A2(new_n978), .A3(new_n704), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n978), .B1(new_n977), .B2(new_n704), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n976), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT61), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n981), .B(new_n982), .ZN(G66));
  INV_X1    g797(.A(G224), .ZN(new_n984));
  OAI21_X1  g798(.A(G953), .B1(new_n388), .B2(new_n984), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n913), .A2(new_n889), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n985), .B1(new_n986), .B2(G953), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n927), .B1(G898), .B2(new_n276), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n987), .B(new_n988), .ZN(G69));
  OAI21_X1  g803(.A(new_n544), .B1(new_n558), .B2(new_n559), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n359), .A2(new_n360), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n990), .B(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(G900), .A2(G953), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n874), .A2(new_n789), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n642), .A2(new_n769), .A3(new_n724), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n807), .B1(new_n824), .B2(new_n995), .ZN(new_n996));
  NOR3_X1   g810(.A1(new_n831), .A2(new_n994), .A3(new_n996), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n997), .A2(new_n805), .A3(new_n826), .ZN(new_n998));
  OAI211_X1 g812(.A(new_n992), .B(new_n993), .C1(new_n998), .C2(G953), .ZN(new_n999));
  NOR3_X1   g813(.A1(new_n722), .A2(new_n893), .A3(new_n797), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n909), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n826), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1002), .A2(KEYINPUT125), .ZN(new_n1003));
  INV_X1    g817(.A(KEYINPUT125), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n826), .A2(new_n1004), .A3(new_n1001), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  AND3_X1   g820(.A1(new_n736), .A2(new_n789), .A3(new_n874), .ZN(new_n1007));
  OR2_X1    g821(.A1(new_n1007), .A2(KEYINPUT62), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1007), .A2(KEYINPUT62), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n831), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g824(.A(G953), .B1(new_n1006), .B2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n999), .B1(new_n1011), .B2(new_n992), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n276), .B1(G227), .B2(G900), .ZN(new_n1013));
  INV_X1    g827(.A(KEYINPUT126), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1013), .B1(new_n999), .B2(new_n1014), .ZN(new_n1015));
  XOR2_X1   g829(.A(new_n1012), .B(new_n1015), .Z(G72));
  AOI21_X1  g830(.A(new_n571), .B1(new_n560), .B2(new_n531), .ZN(new_n1017));
  AND3_X1   g831(.A1(new_n1006), .A2(new_n986), .A3(new_n1010), .ZN(new_n1018));
  NAND2_X1  g832(.A1(G472), .A2(G902), .ZN(new_n1019));
  XOR2_X1   g833(.A(new_n1019), .B(KEYINPUT63), .Z(new_n1020));
  INV_X1    g834(.A(new_n1020), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n1017), .B1(new_n1018), .B2(new_n1021), .ZN(new_n1022));
  OAI211_X1 g836(.A(new_n899), .B(new_n1020), .C1(new_n584), .C2(new_n726), .ZN(new_n1023));
  INV_X1    g837(.A(new_n986), .ZN(new_n1024));
  OAI21_X1  g838(.A(new_n1020), .B1(new_n998), .B2(new_n1024), .ZN(new_n1025));
  AND3_X1   g839(.A1(new_n560), .A2(new_n571), .A3(new_n531), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n924), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g841(.A1(new_n1022), .A2(new_n1023), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g842(.A(KEYINPUT127), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND4_X1  g844(.A1(new_n1022), .A2(KEYINPUT127), .A3(new_n1023), .A4(new_n1027), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1030), .A2(new_n1031), .ZN(G57));
endmodule


