//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 1 0 1 1 0 1 1 1 1 1 1 0 0 0 0 0 0 1 0 1 0 0 1 1 0 0 0 1 0 0 0 1 1 1 1 1 1 0 0 0 0 1 0 0 0 0 1 0 0 1 0 0 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:25 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016;
  INV_X1    g000(.A(G478), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(KEYINPUT15), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT86), .ZN(new_n189));
  INV_X1    g003(.A(G134), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT82), .ZN(new_n191));
  INV_X1    g005(.A(G128), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n191), .B1(new_n192), .B2(G143), .ZN(new_n193));
  INV_X1    g007(.A(G143), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n194), .A2(KEYINPUT82), .A3(G128), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT83), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n192), .A2(G143), .ZN(new_n198));
  AND3_X1   g012(.A1(new_n196), .A2(new_n197), .A3(new_n198), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n197), .B1(new_n196), .B2(new_n198), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n190), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  AND2_X1   g016(.A1(KEYINPUT73), .A2(G107), .ZN(new_n203));
  NOR2_X1   g017(.A1(KEYINPUT73), .A2(G107), .ZN(new_n204));
  OR2_X1    g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  XNOR2_X1  g019(.A(G116), .B(G122), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n205), .A2(new_n206), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT13), .ZN(new_n211));
  AOI22_X1  g025(.A1(new_n196), .A2(new_n211), .B1(new_n192), .B2(G143), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n193), .A2(KEYINPUT13), .A3(new_n195), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n190), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NOR3_X1   g028(.A1(new_n202), .A2(new_n210), .A3(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  AND3_X1   g030(.A1(new_n194), .A2(KEYINPUT82), .A3(G128), .ZN(new_n217));
  AOI21_X1  g031(.A(KEYINPUT82), .B1(new_n194), .B2(G128), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n198), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(KEYINPUT83), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n196), .A2(new_n197), .A3(new_n198), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n220), .A2(G134), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n201), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G122), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT14), .B1(new_n224), .B2(G116), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(G116), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NOR3_X1   g041(.A1(new_n224), .A2(KEYINPUT14), .A3(G116), .ZN(new_n228));
  OAI21_X1  g042(.A(G107), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT84), .ZN(new_n230));
  XNOR2_X1  g044(.A(new_n229), .B(new_n230), .ZN(new_n231));
  AND4_X1   g045(.A1(KEYINPUT85), .A2(new_n223), .A3(new_n207), .A4(new_n231), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n208), .B1(new_n201), .B2(new_n222), .ZN(new_n233));
  AOI21_X1  g047(.A(KEYINPUT85), .B1(new_n233), .B2(new_n231), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n216), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  XOR2_X1   g049(.A(KEYINPUT9), .B(G234), .Z(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G217), .ZN(new_n238));
  NOR3_X1   g052(.A1(new_n237), .A2(new_n238), .A3(G953), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n235), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n223), .A2(new_n207), .A3(new_n231), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT85), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n233), .A2(KEYINPUT85), .A3(new_n231), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n246), .A2(new_n216), .A3(new_n239), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n241), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(G902), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n189), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  AOI211_X1 g064(.A(KEYINPUT86), .B(G902), .C1(new_n241), .C2(new_n247), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n188), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  OAI21_X1  g066(.A(G221), .B1(new_n237), .B2(G902), .ZN(new_n253));
  XOR2_X1   g067(.A(new_n253), .B(KEYINPUT72), .Z(new_n254));
  INV_X1    g068(.A(KEYINPUT10), .ZN(new_n255));
  OAI211_X1 g069(.A(new_n194), .B(G146), .C1(new_n192), .C2(KEYINPUT1), .ZN(new_n256));
  INV_X1    g070(.A(G146), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n192), .A2(new_n257), .A3(G143), .ZN(new_n258));
  AND3_X1   g072(.A1(new_n256), .A2(KEYINPUT64), .A3(new_n258), .ZN(new_n259));
  AOI21_X1  g073(.A(KEYINPUT64), .B1(new_n256), .B2(new_n258), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  XNOR2_X1  g075(.A(G143), .B(G146), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n192), .A2(KEYINPUT1), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n255), .B1(new_n261), .B2(new_n264), .ZN(new_n265));
  NOR3_X1   g079(.A1(new_n203), .A2(new_n204), .A3(G104), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT74), .ZN(new_n267));
  INV_X1    g081(.A(G104), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n267), .B1(new_n268), .B2(G107), .ZN(new_n269));
  INV_X1    g083(.A(G107), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n270), .A2(KEYINPUT74), .A3(G104), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(G101), .B1(new_n266), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT3), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n274), .B(G104), .C1(new_n203), .C2(new_n204), .ZN(new_n275));
  INV_X1    g089(.A(G101), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n268), .A2(G107), .ZN(new_n277));
  OAI21_X1  g091(.A(KEYINPUT3), .B1(new_n268), .B2(G107), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n275), .A2(new_n276), .A3(new_n277), .A4(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n273), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n264), .A2(new_n256), .A3(new_n258), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n282), .A2(new_n273), .A3(new_n279), .ZN(new_n283));
  AOI22_X1  g097(.A1(new_n265), .A2(new_n281), .B1(new_n255), .B2(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n275), .A2(new_n277), .A3(new_n278), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(G101), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n286), .A2(KEYINPUT4), .A3(new_n279), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT0), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n262), .B1(new_n288), .B2(new_n192), .ZN(new_n289));
  XOR2_X1   g103(.A(KEYINPUT0), .B(G128), .Z(new_n290));
  OAI21_X1  g104(.A(new_n289), .B1(new_n262), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT4), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n285), .A2(new_n292), .A3(G101), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n287), .A2(new_n291), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n284), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT11), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n296), .B1(new_n190), .B2(G137), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n190), .A2(G137), .ZN(new_n298));
  INV_X1    g112(.A(G137), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n299), .A2(KEYINPUT11), .A3(G134), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n297), .A2(new_n298), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(G131), .ZN(new_n302));
  INV_X1    g116(.A(G131), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n297), .A2(new_n300), .A3(new_n303), .A4(new_n298), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n295), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n265), .A2(new_n281), .ZN(new_n307));
  INV_X1    g121(.A(new_n305), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n283), .A2(new_n255), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n294), .A2(new_n307), .A3(new_n308), .A4(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(G110), .B(G140), .ZN(new_n311));
  INV_X1    g125(.A(G953), .ZN(new_n312));
  AND2_X1   g126(.A1(new_n312), .A2(G227), .ZN(new_n313));
  XOR2_X1   g127(.A(new_n311), .B(new_n313), .Z(new_n314));
  NAND2_X1  g128(.A1(new_n310), .A2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n257), .A2(G143), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n194), .A2(G146), .ZN(new_n318));
  AND3_X1   g132(.A1(new_n263), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  NOR3_X1   g133(.A1(new_n259), .A2(new_n260), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n280), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(new_n283), .ZN(new_n322));
  AOI21_X1  g136(.A(KEYINPUT12), .B1(new_n322), .B2(new_n305), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT12), .ZN(new_n324));
  AOI211_X1 g138(.A(new_n324), .B(new_n308), .C1(new_n321), .C2(new_n283), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n310), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(new_n314), .ZN(new_n327));
  AOI22_X1  g141(.A1(new_n306), .A2(new_n316), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  OAI21_X1  g142(.A(G469), .B1(new_n328), .B2(G902), .ZN(new_n329));
  INV_X1    g143(.A(new_n310), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n308), .B1(new_n284), .B2(new_n294), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n327), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n310), .B(new_n314), .C1(new_n323), .C2(new_n325), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(G469), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n334), .A2(new_n335), .A3(new_n249), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n254), .B1(new_n329), .B2(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(G902), .B1(new_n241), .B2(new_n247), .ZN(new_n338));
  OAI22_X1  g152(.A1(new_n338), .A2(new_n189), .B1(KEYINPUT15), .B2(new_n187), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n252), .A2(new_n337), .A3(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT78), .ZN(new_n341));
  INV_X1    g155(.A(G237), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n342), .A2(new_n312), .A3(G214), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n194), .A2(KEYINPUT77), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n343), .B(new_n344), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n341), .B1(new_n345), .B2(new_n303), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n343), .A2(KEYINPUT77), .A3(new_n194), .ZN(new_n347));
  NOR2_X1   g161(.A1(G237), .A2(G953), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n344), .A2(G214), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n350), .A2(KEYINPUT78), .A3(G131), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n346), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(G125), .ZN(new_n353));
  NOR3_X1   g167(.A1(new_n353), .A2(KEYINPUT16), .A3(G140), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(G140), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(G125), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n353), .A2(G140), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT16), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n355), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(new_n257), .ZN(new_n362));
  XNOR2_X1  g176(.A(G125), .B(G140), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n354), .B1(new_n363), .B2(KEYINPUT16), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(G146), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT70), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n362), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n364), .A2(KEYINPUT70), .A3(G146), .ZN(new_n368));
  AOI22_X1  g182(.A1(new_n352), .A2(KEYINPUT17), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT17), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n345), .A2(new_n303), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n346), .A2(new_n370), .A3(new_n371), .A4(new_n351), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(KEYINPUT80), .ZN(new_n373));
  AOI21_X1  g187(.A(KEYINPUT78), .B1(new_n350), .B2(G131), .ZN(new_n374));
  AOI211_X1 g188(.A(new_n341), .B(new_n303), .C1(new_n347), .C2(new_n349), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT80), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n376), .A2(new_n377), .A3(new_n370), .A4(new_n371), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n369), .A2(new_n373), .A3(new_n378), .ZN(new_n379));
  XNOR2_X1  g193(.A(G113), .B(G122), .ZN(new_n380));
  XNOR2_X1  g194(.A(new_n380), .B(new_n268), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT18), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n345), .B1(new_n382), .B2(new_n303), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n350), .A2(KEYINPUT18), .A3(G131), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n359), .A2(G146), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n363), .A2(new_n257), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n383), .B(new_n384), .C1(new_n385), .C2(new_n386), .ZN(new_n387));
  AND3_X1   g201(.A1(new_n379), .A2(new_n381), .A3(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n381), .B1(new_n379), .B2(new_n387), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n249), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(KEYINPUT81), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT81), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n392), .B(new_n249), .C1(new_n388), .C2(new_n389), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n391), .A2(G475), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(G234), .A2(G237), .ZN(new_n395));
  AND3_X1   g209(.A1(new_n395), .A2(G952), .A3(new_n312), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  AND3_X1   g211(.A1(new_n395), .A2(G902), .A3(G953), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  XOR2_X1   g213(.A(KEYINPUT21), .B(G898), .Z(new_n400));
  OAI21_X1  g214(.A(new_n397), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n379), .A2(new_n381), .A3(new_n387), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n361), .A2(new_n257), .ZN(new_n403));
  OR2_X1    g217(.A1(new_n359), .A2(KEYINPUT19), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n359), .A2(KEYINPUT19), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n404), .A2(new_n257), .A3(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT79), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n403), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n346), .A2(new_n371), .A3(new_n351), .ZN(new_n409));
  OAI211_X1 g223(.A(new_n408), .B(new_n409), .C1(new_n407), .C2(new_n406), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(new_n387), .ZN(new_n411));
  INV_X1    g225(.A(new_n381), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n402), .A2(new_n413), .ZN(new_n414));
  NOR2_X1   g228(.A1(G475), .A2(G902), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(KEYINPUT20), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT20), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n414), .A2(new_n418), .A3(new_n415), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n394), .A2(new_n401), .A3(new_n420), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n340), .A2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT32), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n256), .A2(new_n258), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT64), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n256), .A2(KEYINPUT64), .A3(new_n258), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n426), .A2(new_n264), .A3(new_n427), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n299), .A2(G134), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n190), .A2(G137), .ZN(new_n430));
  OAI21_X1  g244(.A(G131), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  AND2_X1   g245(.A1(new_n304), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n305), .A2(new_n291), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT30), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AOI22_X1  g251(.A1(new_n432), .A2(new_n428), .B1(new_n305), .B2(new_n291), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(KEYINPUT30), .ZN(new_n439));
  INV_X1    g253(.A(G119), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(G116), .ZN(new_n441));
  INV_X1    g255(.A(G116), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(G119), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  XNOR2_X1  g258(.A(KEYINPUT2), .B(G113), .ZN(new_n445));
  XOR2_X1   g259(.A(new_n444), .B(new_n445), .Z(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n437), .A2(new_n439), .A3(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n433), .A2(new_n434), .A3(new_n446), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(KEYINPUT65), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT65), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n438), .A2(new_n451), .A3(new_n446), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n448), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n348), .A2(G210), .ZN(new_n455));
  XOR2_X1   g269(.A(new_n455), .B(KEYINPUT27), .Z(new_n456));
  XNOR2_X1  g270(.A(new_n456), .B(KEYINPUT26), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n457), .B(G101), .ZN(new_n458));
  NOR3_X1   g272(.A1(new_n454), .A2(new_n458), .A3(KEYINPUT31), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT31), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT28), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n449), .A2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n435), .A2(new_n447), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n451), .B1(new_n438), .B2(new_n446), .ZN(new_n465));
  AND4_X1   g279(.A1(new_n451), .A2(new_n433), .A3(new_n446), .A4(new_n434), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n463), .B1(new_n467), .B2(KEYINPUT28), .ZN(new_n468));
  INV_X1    g282(.A(new_n458), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n460), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n454), .A2(new_n458), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n459), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g287(.A1(G472), .A2(G902), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n423), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n459), .ZN(new_n477));
  AOI22_X1  g291(.A1(new_n450), .A2(new_n452), .B1(new_n447), .B2(new_n435), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n462), .B1(new_n478), .B2(new_n461), .ZN(new_n479));
  AOI21_X1  g293(.A(KEYINPUT31), .B1(new_n479), .B2(new_n458), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n477), .B1(new_n480), .B2(new_n471), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n481), .A2(KEYINPUT32), .A3(new_n474), .ZN(new_n482));
  AOI21_X1  g296(.A(KEYINPUT29), .B1(new_n454), .B2(new_n458), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n483), .B1(new_n458), .B2(new_n479), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n468), .A2(KEYINPUT29), .A3(new_n469), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n484), .A2(new_n249), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(G472), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n476), .A2(new_n482), .A3(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n312), .A2(G221), .A3(G234), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n489), .B(KEYINPUT22), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n490), .B(G137), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n403), .A2(new_n385), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT68), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n494), .A2(KEYINPUT23), .ZN(new_n495));
  OAI21_X1  g309(.A(KEYINPUT68), .B1(new_n440), .B2(G128), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n495), .B1(new_n496), .B2(KEYINPUT23), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n440), .A2(G128), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT69), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n192), .A2(G119), .ZN(new_n500));
  AOI22_X1  g314(.A1(new_n497), .A2(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  OR3_X1    g315(.A1(new_n500), .A2(new_n499), .A3(KEYINPUT23), .ZN(new_n502));
  AOI21_X1  g316(.A(G110), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  XOR2_X1   g317(.A(KEYINPUT24), .B(G110), .Z(new_n504));
  XNOR2_X1  g318(.A(new_n498), .B(KEYINPUT67), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n504), .B1(new_n505), .B2(new_n500), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n493), .B1(new_n503), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n505), .A2(new_n500), .A3(new_n504), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n497), .A2(new_n498), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n500), .A2(new_n499), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n509), .A2(G110), .A3(new_n510), .A4(new_n502), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n367), .A2(new_n508), .A3(new_n368), .A4(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT71), .ZN(new_n513));
  AND3_X1   g327(.A1(new_n507), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n513), .B1(new_n507), .B2(new_n512), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n492), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n507), .A2(new_n512), .A3(new_n491), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n516), .A2(new_n249), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(KEYINPUT25), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n238), .B1(G234), .B2(new_n249), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT66), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT25), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n516), .A2(new_n523), .A3(new_n249), .A4(new_n517), .ZN(new_n524));
  OR2_X1    g338(.A1(new_n520), .A2(new_n521), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n519), .A2(new_n522), .A3(new_n524), .A4(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n516), .A2(new_n517), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n520), .A2(G902), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n526), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(G210), .B1(G237), .B2(G902), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n287), .A2(new_n447), .A3(new_n293), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n441), .A2(new_n443), .A3(KEYINPUT5), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n536), .B1(KEYINPUT5), .B2(new_n441), .ZN(new_n537));
  INV_X1    g351(.A(G113), .ZN(new_n538));
  OAI22_X1  g352(.A1(new_n537), .A2(new_n538), .B1(new_n444), .B2(new_n445), .ZN(new_n539));
  OR2_X1    g353(.A1(new_n539), .A2(new_n280), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n535), .A2(new_n540), .ZN(new_n541));
  XOR2_X1   g355(.A(G110), .B(G122), .Z(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n542), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n535), .A2(new_n540), .A3(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n543), .A2(KEYINPUT6), .A3(new_n545), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n289), .B(G125), .C1(new_n262), .C2(new_n290), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n547), .B1(new_n428), .B2(G125), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(KEYINPUT75), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT75), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(G224), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n553), .A2(G953), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n554), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n549), .A2(new_n556), .A3(new_n551), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT6), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n541), .A2(new_n559), .A3(new_n542), .ZN(new_n560));
  AND3_X1   g374(.A1(new_n546), .A2(new_n558), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n556), .A2(KEYINPUT7), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n563), .B1(new_n549), .B2(new_n551), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n549), .A2(new_n551), .A3(new_n563), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n539), .A2(new_n280), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n539), .A2(new_n280), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(KEYINPUT76), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT76), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n539), .A2(new_n280), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n568), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  XOR2_X1   g387(.A(new_n542), .B(KEYINPUT8), .Z(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n545), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n249), .B1(new_n567), .B2(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n534), .B1(new_n561), .B2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n576), .ZN(new_n579));
  INV_X1    g393(.A(new_n566), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n580), .A2(new_n564), .ZN(new_n581));
  AOI21_X1  g395(.A(G902), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n546), .A2(new_n558), .A3(new_n560), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n582), .A2(new_n533), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n578), .A2(new_n584), .ZN(new_n585));
  OAI21_X1  g399(.A(G214), .B1(G237), .B2(G902), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n422), .A2(new_n488), .A3(new_n532), .A4(new_n588), .ZN(new_n589));
  XOR2_X1   g403(.A(KEYINPUT87), .B(G101), .Z(new_n590));
  XNOR2_X1  g404(.A(new_n589), .B(new_n590), .ZN(G3));
  NAND3_X1  g405(.A1(new_n578), .A2(new_n584), .A3(KEYINPUT88), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT88), .ZN(new_n593));
  OAI211_X1 g407(.A(new_n593), .B(new_n534), .C1(new_n561), .C2(new_n577), .ZN(new_n594));
  AND3_X1   g408(.A1(new_n592), .A2(new_n586), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n248), .A2(new_n249), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(new_n187), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT33), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n248), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n241), .A2(new_n247), .A3(KEYINPUT33), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n599), .A2(G478), .A3(new_n249), .A4(new_n600), .ZN(new_n601));
  AOI22_X1  g415(.A1(new_n597), .A2(new_n601), .B1(new_n394), .B2(new_n420), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n595), .A2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n254), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n326), .A2(new_n327), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n306), .A2(new_n310), .A3(new_n314), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n605), .A2(G469), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(G469), .A2(G902), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  AOI211_X1 g423(.A(G469), .B(G902), .C1(new_n332), .C2(new_n333), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n604), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n401), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n481), .A2(new_n474), .ZN(new_n614));
  OAI21_X1  g428(.A(G472), .B1(new_n473), .B2(G902), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n613), .A2(new_n532), .A3(new_n614), .A4(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n603), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(KEYINPUT89), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(KEYINPUT34), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(new_n268), .ZN(G6));
  AOI21_X1  g434(.A(KEYINPUT90), .B1(new_n416), .B2(KEYINPUT20), .ZN(new_n621));
  INV_X1    g435(.A(new_n415), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n622), .B1(new_n402), .B2(new_n413), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT90), .ZN(new_n624));
  NOR3_X1   g438(.A1(new_n623), .A2(new_n624), .A3(new_n418), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT91), .ZN(new_n626));
  AND4_X1   g440(.A1(new_n626), .A2(new_n414), .A3(new_n418), .A4(new_n415), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n626), .B1(new_n623), .B2(new_n418), .ZN(new_n628));
  OAI22_X1  g442(.A1(new_n621), .A2(new_n625), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT92), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n416), .A2(KEYINPUT90), .A3(KEYINPUT20), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n624), .B1(new_n623), .B2(new_n418), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n419), .A2(KEYINPUT91), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n623), .A2(new_n626), .A3(new_n418), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n634), .A2(new_n637), .A3(KEYINPUT92), .ZN(new_n638));
  AND3_X1   g452(.A1(new_n631), .A2(new_n394), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n252), .A2(new_n339), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n639), .A2(new_n640), .A3(new_n595), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n641), .A2(new_n616), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(KEYINPUT93), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(KEYINPUT35), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(new_n270), .ZN(G9));
  NOR2_X1   g459(.A1(new_n492), .A2(KEYINPUT36), .ZN(new_n646));
  XOR2_X1   g460(.A(new_n646), .B(KEYINPUT94), .Z(new_n647));
  OR2_X1    g461(.A1(new_n514), .A2(new_n515), .ZN(new_n648));
  AND2_X1   g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n647), .A2(new_n648), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n529), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n526), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n615), .A2(new_n652), .A3(new_n614), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT95), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n615), .A2(new_n652), .A3(KEYINPUT95), .A4(new_n614), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n655), .A2(new_n422), .A3(new_n588), .A4(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(KEYINPUT96), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT37), .B(G110), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G12));
  INV_X1    g474(.A(G900), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n396), .B1(new_n398), .B2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n639), .A2(new_n640), .A3(new_n663), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n488), .A2(new_n595), .A3(new_n337), .A4(new_n652), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(new_n192), .ZN(G30));
  XOR2_X1   g481(.A(new_n662), .B(KEYINPUT39), .Z(new_n668));
  NAND2_X1  g482(.A1(new_n337), .A2(new_n668), .ZN(new_n669));
  OR2_X1    g483(.A1(new_n669), .A2(KEYINPUT40), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(KEYINPUT40), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n585), .B(KEYINPUT38), .ZN(new_n672));
  AND4_X1   g486(.A1(new_n586), .A2(new_n670), .A3(new_n671), .A4(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n652), .ZN(new_n674));
  AND2_X1   g488(.A1(new_n476), .A2(new_n482), .ZN(new_n675));
  INV_X1    g489(.A(new_n454), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n676), .A2(new_n458), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n249), .B1(new_n469), .B2(new_n467), .ZN(new_n678));
  OAI21_X1  g492(.A(G472), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n675), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n250), .A2(new_n188), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n596), .A2(KEYINPUT86), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n338), .A2(new_n189), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n681), .B1(new_n684), .B2(new_n188), .ZN(new_n685));
  AND2_X1   g499(.A1(new_n394), .A2(new_n420), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n673), .A2(new_n674), .A3(new_n680), .A4(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(KEYINPUT97), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(new_n194), .ZN(G45));
  AND3_X1   g504(.A1(new_n488), .A2(new_n337), .A3(new_n652), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n601), .A2(new_n597), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n394), .A2(new_n420), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n694), .A2(new_n662), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n691), .A2(KEYINPUT98), .A3(new_n595), .A4(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT98), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n602), .A2(new_n663), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n697), .B1(new_n665), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G146), .ZN(G48));
  AND2_X1   g515(.A1(new_n488), .A2(new_n532), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n592), .A2(new_n594), .A3(new_n586), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n694), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n334), .A2(new_n249), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(G469), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n706), .A2(new_n401), .A3(new_n604), .A4(new_n336), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n702), .A2(KEYINPUT99), .A3(new_n704), .A4(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT99), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n488), .A2(new_n532), .A3(new_n708), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n710), .B1(new_n711), .B2(new_n603), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n709), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(KEYINPUT41), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G113), .ZN(G15));
  OAI21_X1  g529(.A(KEYINPUT100), .B1(new_n641), .B2(new_n711), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n631), .A2(new_n640), .A3(new_n394), .A4(new_n638), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n717), .A2(new_n703), .ZN(new_n718));
  INV_X1    g532(.A(new_n711), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT100), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n718), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n716), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G116), .ZN(G18));
  AND3_X1   g537(.A1(new_n706), .A2(new_n604), .A3(new_n336), .ZN(new_n724));
  AND4_X1   g538(.A1(new_n488), .A2(new_n595), .A3(new_n652), .A4(new_n724), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n640), .A2(new_n421), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G119), .ZN(G21));
  OAI211_X1 g542(.A(KEYINPUT101), .B(new_n477), .C1(new_n480), .C2(new_n471), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT101), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n470), .A2(new_n730), .A3(new_n472), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n729), .A2(new_n474), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n615), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT102), .ZN(new_n734));
  AND3_X1   g548(.A1(new_n526), .A2(new_n734), .A3(new_n530), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n734), .B1(new_n526), .B2(new_n530), .ZN(new_n736));
  NOR4_X1   g550(.A1(new_n733), .A2(new_n735), .A3(new_n736), .A4(new_n707), .ZN(new_n737));
  NOR3_X1   g551(.A1(new_n685), .A2(new_n703), .A3(new_n686), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(KEYINPUT103), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G122), .ZN(G24));
  NAND3_X1  g555(.A1(new_n732), .A2(new_n615), .A3(new_n652), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT104), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n732), .A2(new_n615), .A3(KEYINPUT104), .A4(new_n652), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n698), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(new_n724), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n747), .A2(new_n703), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G125), .ZN(G27));
  INV_X1    g564(.A(KEYINPUT107), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n611), .A2(KEYINPUT105), .ZN(new_n752));
  AND3_X1   g566(.A1(new_n578), .A2(new_n584), .A3(new_n586), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n336), .A2(new_n608), .A3(new_n607), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT105), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n754), .A2(new_n755), .A3(new_n604), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n752), .A2(new_n753), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(KEYINPUT106), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT106), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n752), .A2(new_n759), .A3(new_n756), .A4(new_n753), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(new_n488), .ZN(new_n762));
  INV_X1    g576(.A(new_n736), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n526), .A2(new_n734), .A3(new_n530), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n761), .A2(new_n766), .A3(KEYINPUT42), .A4(new_n695), .ZN(new_n767));
  INV_X1    g581(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n488), .A2(new_n532), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n769), .B1(new_n758), .B2(new_n760), .ZN(new_n770));
  AOI21_X1  g584(.A(KEYINPUT42), .B1(new_n770), .B2(new_n695), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n751), .B1(new_n768), .B2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n761), .A2(new_n702), .A3(new_n695), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT42), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n775), .A2(KEYINPUT107), .A3(new_n767), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n772), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G131), .ZN(G33));
  INV_X1    g592(.A(KEYINPUT108), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n664), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n717), .A2(new_n662), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(KEYINPUT108), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n780), .A2(new_n770), .A3(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G134), .ZN(G36));
  INV_X1    g598(.A(new_n753), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n686), .A2(new_n692), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT43), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n473), .A2(new_n475), .ZN(new_n789));
  INV_X1    g603(.A(G472), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n790), .B1(new_n481), .B2(new_n249), .ZN(new_n791));
  OAI211_X1 g605(.A(new_n788), .B(new_n652), .C1(new_n789), .C2(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(new_n792), .ZN(new_n793));
  OR2_X1    g607(.A1(new_n793), .A2(KEYINPUT44), .ZN(new_n794));
  XOR2_X1   g608(.A(new_n328), .B(KEYINPUT45), .Z(new_n795));
  OAI21_X1  g609(.A(G469), .B1(new_n795), .B2(G902), .ZN(new_n796));
  OR3_X1    g610(.A1(new_n796), .A2(KEYINPUT109), .A3(KEYINPUT46), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(KEYINPUT46), .ZN(new_n798));
  OAI21_X1  g612(.A(KEYINPUT109), .B1(new_n796), .B2(KEYINPUT46), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n797), .A2(new_n336), .A3(new_n798), .A4(new_n799), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n800), .A2(new_n604), .A3(new_n668), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n794), .A2(new_n801), .ZN(new_n802));
  AOI211_X1 g616(.A(new_n785), .B(new_n802), .C1(KEYINPUT44), .C2(new_n793), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(KEYINPUT110), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(new_n299), .ZN(G39));
  INV_X1    g619(.A(KEYINPUT111), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(KEYINPUT47), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n807), .B1(new_n800), .B2(new_n604), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n800), .A2(new_n604), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n809), .B1(new_n806), .B2(KEYINPUT47), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n808), .B1(new_n810), .B2(new_n807), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n811), .A2(new_n695), .A3(new_n753), .ZN(new_n812));
  NOR3_X1   g626(.A1(new_n812), .A2(new_n488), .A3(new_n532), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(new_n356), .ZN(G42));
  NAND2_X1  g628(.A1(new_n312), .A2(G952), .ZN(new_n815));
  INV_X1    g629(.A(new_n680), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n747), .A2(new_n785), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n816), .A2(new_n532), .A3(new_n817), .A4(new_n396), .ZN(new_n818));
  INV_X1    g632(.A(new_n818), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n815), .B1(new_n819), .B2(new_n602), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n788), .A2(new_n396), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n821), .A2(new_n817), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(new_n766), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT48), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(KEYINPUT118), .ZN(new_n825));
  XOR2_X1   g639(.A(new_n823), .B(new_n825), .Z(new_n826));
  OAI21_X1  g640(.A(new_n826), .B1(KEYINPUT118), .B2(new_n824), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n765), .A2(new_n733), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n821), .A2(new_n828), .ZN(new_n829));
  NOR4_X1   g643(.A1(new_n829), .A2(new_n586), .A3(new_n672), .A4(new_n747), .ZN(new_n830));
  XOR2_X1   g644(.A(new_n830), .B(KEYINPUT50), .Z(new_n831));
  NOR3_X1   g645(.A1(new_n818), .A2(new_n693), .A3(new_n692), .ZN(new_n832));
  INV_X1    g646(.A(new_n829), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n706), .A2(new_n336), .ZN(new_n834));
  INV_X1    g648(.A(new_n834), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n835), .A2(new_n604), .ZN(new_n836));
  OAI211_X1 g650(.A(new_n753), .B(new_n833), .C1(new_n811), .C2(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n744), .A2(new_n745), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n822), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n831), .A2(new_n832), .A3(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT51), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n842), .B1(new_n837), .B2(KEYINPUT117), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n820), .B(new_n827), .C1(new_n841), .C2(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n844), .B1(new_n843), .B2(new_n841), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n833), .A2(new_n748), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n685), .A2(new_n693), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n754), .A2(new_n401), .A3(new_n604), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n848), .A2(new_n791), .A3(new_n789), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n847), .A2(new_n849), .A3(new_n532), .A4(new_n588), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT113), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n657), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n851), .B1(new_n657), .B2(new_n850), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n849), .A2(new_n532), .A3(new_n588), .A4(new_n602), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT112), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n589), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n855), .B1(new_n589), .B2(new_n854), .ZN(new_n857));
  OAI22_X1  g671(.A1(new_n852), .A2(new_n853), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  AOI22_X1  g672(.A1(new_n726), .A2(new_n725), .B1(new_n737), .B2(new_n738), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n720), .B1(new_n718), .B2(new_n719), .ZN(new_n860));
  NOR4_X1   g674(.A1(new_n711), .A2(new_n717), .A3(KEYINPUT100), .A4(new_n703), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n713), .B(new_n859), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n761), .A2(new_n838), .A3(new_n602), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n762), .A2(new_n674), .ZN(new_n864));
  INV_X1    g678(.A(new_n340), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n864), .A2(new_n639), .A3(new_n865), .A4(new_n753), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n662), .B1(new_n863), .B2(new_n866), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n858), .A2(new_n862), .A3(new_n867), .ZN(new_n868));
  AND4_X1   g682(.A1(new_n488), .A2(new_n595), .A3(new_n337), .A4(new_n652), .ZN(new_n869));
  AOI22_X1  g683(.A1(new_n746), .A2(new_n748), .B1(new_n781), .B2(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n611), .A2(new_n662), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n738), .A2(new_n680), .A3(new_n674), .A4(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n870), .A2(new_n700), .A3(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT52), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n870), .A2(new_n700), .A3(KEYINPUT52), .A4(new_n872), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(new_n783), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n878), .B1(new_n772), .B2(new_n776), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n868), .A2(new_n877), .A3(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT53), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n880), .A2(new_n881), .ZN(new_n884));
  OAI21_X1  g698(.A(KEYINPUT54), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n882), .A2(KEYINPUT114), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT114), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n880), .A2(new_n887), .A3(new_n881), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n657), .A2(new_n850), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(KEYINPUT113), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n657), .A2(new_n850), .A3(new_n851), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(new_n421), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n685), .A2(new_n893), .A3(new_n588), .A4(new_n337), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n894), .A2(new_n769), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n616), .A2(new_n587), .A3(new_n694), .ZN(new_n896));
  OAI21_X1  g710(.A(KEYINPUT112), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n589), .A2(new_n854), .A3(new_n855), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n892), .A2(KEYINPUT53), .A3(new_n899), .A4(new_n783), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT115), .ZN(new_n901));
  AOI211_X1 g715(.A(new_n774), .B(new_n698), .C1(new_n758), .C2(new_n760), .ZN(new_n902));
  AOI22_X1  g716(.A1(new_n766), .A2(new_n902), .B1(new_n773), .B2(new_n774), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n901), .B1(new_n862), .B2(new_n903), .ZN(new_n904));
  AND2_X1   g718(.A1(new_n713), .A2(new_n859), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n775), .A2(new_n767), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n905), .A2(new_n906), .A3(KEYINPUT115), .A4(new_n722), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n900), .B1(new_n904), .B2(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n867), .B1(new_n875), .B2(new_n876), .ZN(new_n909));
  AOI21_X1  g723(.A(KEYINPUT116), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n904), .A2(new_n907), .ZN(new_n911));
  INV_X1    g725(.A(new_n900), .ZN(new_n912));
  AND4_X1   g726(.A1(KEYINPUT116), .A2(new_n911), .A3(new_n912), .A4(new_n909), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n886), .B(new_n888), .C1(new_n910), .C2(new_n913), .ZN(new_n914));
  OR2_X1    g728(.A1(new_n914), .A2(KEYINPUT54), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n845), .A2(new_n846), .A3(new_n885), .A4(new_n915), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n916), .B1(G952), .B2(G953), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT49), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n604), .B1(new_n834), .B2(new_n918), .ZN(new_n919));
  AOI211_X1 g733(.A(new_n919), .B(new_n786), .C1(new_n918), .C2(new_n834), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n765), .A2(new_n672), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n920), .A2(new_n586), .A3(new_n816), .A4(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n917), .A2(new_n922), .ZN(G75));
  NOR2_X1   g737(.A1(new_n312), .A2(G952), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(KEYINPUT120), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n886), .A2(new_n888), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n913), .A2(new_n910), .ZN(new_n927));
  OAI21_X1  g741(.A(G902), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(KEYINPUT56), .B1(new_n929), .B2(G210), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n546), .A2(new_n560), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(new_n558), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT55), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n925), .B1(new_n930), .B2(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT56), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n928), .A2(KEYINPUT119), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT119), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n914), .A2(new_n938), .A3(G902), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n936), .B1(new_n940), .B2(new_n534), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n934), .A2(new_n941), .ZN(G51));
  INV_X1    g756(.A(KEYINPUT122), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n795), .A2(G469), .ZN(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n943), .B1(new_n940), .B2(new_n945), .ZN(new_n946));
  AOI211_X1 g760(.A(KEYINPUT122), .B(new_n944), .C1(new_n937), .C2(new_n939), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n914), .A2(KEYINPUT54), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n915), .A2(new_n949), .A3(KEYINPUT121), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT121), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n914), .A2(new_n951), .A3(KEYINPUT54), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n608), .B(KEYINPUT57), .Z(new_n953));
  NAND3_X1  g767(.A1(new_n950), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n334), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n924), .B1(new_n948), .B2(new_n955), .ZN(G54));
  NAND3_X1  g770(.A1(new_n940), .A2(KEYINPUT58), .A3(G475), .ZN(new_n957));
  INV_X1    g771(.A(new_n414), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(new_n924), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n940), .A2(KEYINPUT58), .A3(G475), .A4(new_n414), .ZN(new_n961));
  AND3_X1   g775(.A1(new_n959), .A2(new_n960), .A3(new_n961), .ZN(G60));
  AND2_X1   g776(.A1(new_n599), .A2(new_n600), .ZN(new_n963));
  NAND2_X1  g777(.A1(G478), .A2(G902), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(KEYINPUT59), .Z(new_n965));
  INV_X1    g779(.A(new_n965), .ZN(new_n966));
  AND4_X1   g780(.A1(new_n963), .A2(new_n950), .A3(new_n952), .A4(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n965), .B1(new_n915), .B2(new_n885), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n925), .B1(new_n968), .B2(new_n963), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n967), .A2(new_n969), .ZN(G63));
  XNOR2_X1  g784(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n238), .A2(new_n249), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n971), .B(new_n972), .ZN(new_n973));
  OAI211_X1 g787(.A(new_n914), .B(new_n973), .C1(new_n650), .C2(new_n649), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n914), .A2(new_n973), .ZN(new_n975));
  OAI211_X1 g789(.A(new_n974), .B(new_n925), .C1(new_n975), .C2(new_n528), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n976), .B(KEYINPUT61), .Z(G66));
  AOI21_X1  g791(.A(new_n312), .B1(new_n400), .B2(G224), .ZN(new_n978));
  OR2_X1    g792(.A1(new_n858), .A2(new_n862), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n978), .B1(new_n979), .B2(new_n312), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n931), .B1(G898), .B2(new_n312), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n981), .B(KEYINPUT124), .Z(new_n982));
  XNOR2_X1  g796(.A(new_n980), .B(new_n982), .ZN(G69));
  NAND2_X1  g797(.A1(G900), .A2(G953), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n437), .A2(new_n439), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n404), .A2(new_n405), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n985), .B(new_n986), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n803), .A2(new_n813), .ZN(new_n988));
  AND2_X1   g802(.A1(new_n870), .A2(new_n700), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n801), .A2(new_n738), .A3(new_n766), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n988), .A2(new_n989), .A3(new_n879), .A4(new_n990), .ZN(new_n991));
  OAI211_X1 g805(.A(new_n984), .B(new_n987), .C1(new_n991), .C2(G953), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n702), .B1(new_n602), .B2(new_n847), .ZN(new_n993));
  OR3_X1    g807(.A1(new_n993), .A2(new_n669), .A3(new_n785), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT62), .ZN(new_n995));
  OAI211_X1 g809(.A(new_n989), .B(new_n688), .C1(KEYINPUT126), .C2(new_n995), .ZN(new_n996));
  AND2_X1   g810(.A1(new_n995), .A2(KEYINPUT126), .ZN(new_n997));
  AND2_X1   g811(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n996), .A2(new_n997), .ZN(new_n999));
  OAI211_X1 g813(.A(new_n988), .B(new_n994), .C1(new_n998), .C2(new_n999), .ZN(new_n1000));
  AND2_X1   g814(.A1(new_n1000), .A2(new_n312), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n987), .B(KEYINPUT125), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n992), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n312), .B1(G227), .B2(G900), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1003), .B(new_n1004), .ZN(G72));
  XNOR2_X1  g819(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n790), .A2(new_n249), .ZN(new_n1007));
  XNOR2_X1  g821(.A(new_n1006), .B(new_n1007), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n1008), .B1(new_n1000), .B2(new_n979), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n924), .B1(new_n1009), .B2(new_n677), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n1008), .B1(new_n991), .B2(new_n979), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n469), .A2(new_n454), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g827(.A(new_n1008), .ZN(new_n1014));
  NOR2_X1   g828(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1015));
  OAI221_X1 g829(.A(new_n1015), .B1(new_n676), .B2(new_n458), .C1(new_n883), .C2(new_n884), .ZN(new_n1016));
  AND3_X1   g830(.A1(new_n1010), .A2(new_n1013), .A3(new_n1016), .ZN(G57));
endmodule


