

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U560 ( .A1(G164), .A2(G1384), .ZN(n790) );
  NAND2_X2 U561 ( .A1(n790), .A2(n788), .ZN(n746) );
  INV_X1 U562 ( .A(KEYINPUT96), .ZN(n715) );
  INV_X1 U563 ( .A(KEYINPUT29), .ZN(n725) );
  XNOR2_X1 U564 ( .A(n726), .B(n725), .ZN(n732) );
  AND2_X1 U565 ( .A1(n697), .A2(G40), .ZN(n788) );
  NOR2_X1 U566 ( .A1(G2105), .A2(G2104), .ZN(n525) );
  INV_X1 U567 ( .A(G651), .ZN(n551) );
  NOR2_X2 U568 ( .A1(G2105), .A2(n529), .ZN(n898) );
  NOR2_X1 U569 ( .A1(n820), .A2(n819), .ZN(n822) );
  XOR2_X1 U570 ( .A(KEYINPUT71), .B(n601), .Z(n934) );
  XOR2_X1 U571 ( .A(KEYINPUT66), .B(n525), .Z(n526) );
  XNOR2_X2 U572 ( .A(n526), .B(KEYINPUT17), .ZN(n899) );
  NAND2_X1 U573 ( .A1(n899), .A2(G138), .ZN(n534) );
  INV_X1 U574 ( .A(G2104), .ZN(n529) );
  AND2_X1 U575 ( .A1(n529), .A2(G2105), .ZN(n906) );
  NAND2_X1 U576 ( .A1(G126), .A2(n906), .ZN(n528) );
  AND2_X1 U577 ( .A1(G2105), .A2(G2104), .ZN(n903) );
  NAND2_X1 U578 ( .A1(G114), .A2(n903), .ZN(n527) );
  AND2_X1 U579 ( .A1(n528), .A2(n527), .ZN(n532) );
  NAND2_X1 U580 ( .A1(G102), .A2(n898), .ZN(n530) );
  XOR2_X1 U581 ( .A(KEYINPUT87), .B(n530), .Z(n531) );
  AND2_X1 U582 ( .A1(n532), .A2(n531), .ZN(n533) );
  AND2_X1 U583 ( .A1(n534), .A2(n533), .ZN(G164) );
  XNOR2_X1 U584 ( .A(G2451), .B(G2443), .ZN(n544) );
  XOR2_X1 U585 ( .A(G2446), .B(KEYINPUT105), .Z(n536) );
  XNOR2_X1 U586 ( .A(KEYINPUT106), .B(G2438), .ZN(n535) );
  XNOR2_X1 U587 ( .A(n536), .B(n535), .ZN(n540) );
  XOR2_X1 U588 ( .A(G2435), .B(G2454), .Z(n538) );
  XNOR2_X1 U589 ( .A(G1341), .B(G1348), .ZN(n537) );
  XNOR2_X1 U590 ( .A(n538), .B(n537), .ZN(n539) );
  XOR2_X1 U591 ( .A(n540), .B(n539), .Z(n542) );
  XNOR2_X1 U592 ( .A(G2430), .B(G2427), .ZN(n541) );
  XNOR2_X1 U593 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U594 ( .A(n544), .B(n543), .ZN(n545) );
  AND2_X1 U595 ( .A1(n545), .A2(G14), .ZN(G401) );
  XOR2_X1 U596 ( .A(G543), .B(KEYINPUT0), .Z(n662) );
  NOR2_X1 U597 ( .A1(G651), .A2(n662), .ZN(n546) );
  XOR2_X1 U598 ( .A(KEYINPUT65), .B(n546), .Z(n667) );
  NAND2_X1 U599 ( .A1(n667), .A2(G52), .ZN(n550) );
  NOR2_X1 U600 ( .A1(G543), .A2(n551), .ZN(n547) );
  XOR2_X1 U601 ( .A(KEYINPUT68), .B(n547), .Z(n548) );
  XNOR2_X2 U602 ( .A(KEYINPUT1), .B(n548), .ZN(n666) );
  NAND2_X1 U603 ( .A1(G64), .A2(n666), .ZN(n549) );
  NAND2_X1 U604 ( .A1(n550), .A2(n549), .ZN(n557) );
  NOR2_X1 U605 ( .A1(n662), .A2(n551), .ZN(n652) );
  NAND2_X1 U606 ( .A1(G77), .A2(n652), .ZN(n554) );
  NOR2_X1 U607 ( .A1(G543), .A2(G651), .ZN(n552) );
  XNOR2_X1 U608 ( .A(n552), .B(KEYINPUT64), .ZN(n655) );
  NAND2_X1 U609 ( .A1(G90), .A2(n655), .ZN(n553) );
  NAND2_X1 U610 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U611 ( .A(KEYINPUT9), .B(n555), .Z(n556) );
  NOR2_X1 U612 ( .A1(n557), .A2(n556), .ZN(G171) );
  AND2_X1 U613 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U614 ( .A1(n903), .A2(G113), .ZN(n560) );
  NAND2_X1 U615 ( .A1(G101), .A2(n898), .ZN(n558) );
  XOR2_X1 U616 ( .A(KEYINPUT23), .B(n558), .Z(n559) );
  NAND2_X1 U617 ( .A1(n560), .A2(n559), .ZN(n564) );
  NAND2_X1 U618 ( .A1(G125), .A2(n906), .ZN(n562) );
  NAND2_X1 U619 ( .A1(G137), .A2(n899), .ZN(n561) );
  NAND2_X1 U620 ( .A1(n562), .A2(n561), .ZN(n563) );
  NOR2_X1 U621 ( .A1(n564), .A2(n563), .ZN(n697) );
  BUF_X1 U622 ( .A(n697), .Z(G160) );
  INV_X1 U623 ( .A(G57), .ZN(G237) );
  INV_X1 U624 ( .A(G132), .ZN(G219) );
  INV_X1 U625 ( .A(G82), .ZN(G220) );
  NAND2_X1 U626 ( .A1(G75), .A2(n652), .ZN(n566) );
  NAND2_X1 U627 ( .A1(G88), .A2(n655), .ZN(n565) );
  NAND2_X1 U628 ( .A1(n566), .A2(n565), .ZN(n570) );
  NAND2_X1 U629 ( .A1(n667), .A2(G50), .ZN(n568) );
  NAND2_X1 U630 ( .A1(G62), .A2(n666), .ZN(n567) );
  NAND2_X1 U631 ( .A1(n568), .A2(n567), .ZN(n569) );
  NOR2_X1 U632 ( .A1(n570), .A2(n569), .ZN(G166) );
  NAND2_X1 U633 ( .A1(n667), .A2(G51), .ZN(n572) );
  NAND2_X1 U634 ( .A1(G63), .A2(n666), .ZN(n571) );
  NAND2_X1 U635 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U636 ( .A(n573), .B(KEYINPUT6), .ZN(n574) );
  XNOR2_X1 U637 ( .A(n574), .B(KEYINPUT75), .ZN(n581) );
  XNOR2_X1 U638 ( .A(KEYINPUT74), .B(KEYINPUT5), .ZN(n579) );
  NAND2_X1 U639 ( .A1(G89), .A2(n655), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n575), .B(KEYINPUT4), .ZN(n577) );
  NAND2_X1 U641 ( .A1(G76), .A2(n652), .ZN(n576) );
  NAND2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n579), .B(n578), .ZN(n580) );
  NAND2_X1 U644 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U645 ( .A(KEYINPUT7), .B(n582), .ZN(G168) );
  XOR2_X1 U646 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U647 ( .A1(n667), .A2(G53), .ZN(n584) );
  NAND2_X1 U648 ( .A1(G91), .A2(n655), .ZN(n583) );
  NAND2_X1 U649 ( .A1(n584), .A2(n583), .ZN(n587) );
  NAND2_X1 U650 ( .A1(n652), .A2(G78), .ZN(n585) );
  XOR2_X1 U651 ( .A(KEYINPUT70), .B(n585), .Z(n586) );
  NOR2_X1 U652 ( .A1(n587), .A2(n586), .ZN(n589) );
  NAND2_X1 U653 ( .A1(G65), .A2(n666), .ZN(n588) );
  NAND2_X1 U654 ( .A1(n589), .A2(n588), .ZN(G299) );
  NAND2_X1 U655 ( .A1(G7), .A2(G661), .ZN(n590) );
  XNOR2_X1 U656 ( .A(n590), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U657 ( .A(G223), .ZN(n841) );
  NAND2_X1 U658 ( .A1(n841), .A2(G567), .ZN(n591) );
  XOR2_X1 U659 ( .A(KEYINPUT11), .B(n591), .Z(G234) );
  NAND2_X1 U660 ( .A1(G81), .A2(n655), .ZN(n592) );
  XNOR2_X1 U661 ( .A(n592), .B(KEYINPUT12), .ZN(n594) );
  NAND2_X1 U662 ( .A1(G68), .A2(n652), .ZN(n593) );
  NAND2_X1 U663 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U664 ( .A(n595), .B(KEYINPUT13), .ZN(n597) );
  NAND2_X1 U665 ( .A1(G43), .A2(n667), .ZN(n596) );
  NAND2_X1 U666 ( .A1(n597), .A2(n596), .ZN(n600) );
  AND2_X1 U667 ( .A1(n666), .A2(G56), .ZN(n598) );
  XNOR2_X1 U668 ( .A(KEYINPUT14), .B(n598), .ZN(n599) );
  NOR2_X1 U669 ( .A1(n600), .A2(n599), .ZN(n601) );
  NAND2_X1 U670 ( .A1(G860), .A2(n934), .ZN(n602) );
  XNOR2_X1 U671 ( .A(n602), .B(KEYINPUT72), .ZN(G153) );
  XNOR2_X1 U672 ( .A(G171), .B(KEYINPUT73), .ZN(G301) );
  NAND2_X1 U673 ( .A1(G868), .A2(G301), .ZN(n611) );
  NAND2_X1 U674 ( .A1(G79), .A2(n652), .ZN(n604) );
  NAND2_X1 U675 ( .A1(G92), .A2(n655), .ZN(n603) );
  NAND2_X1 U676 ( .A1(n604), .A2(n603), .ZN(n608) );
  NAND2_X1 U677 ( .A1(n667), .A2(G54), .ZN(n606) );
  NAND2_X1 U678 ( .A1(G66), .A2(n666), .ZN(n605) );
  NAND2_X1 U679 ( .A1(n606), .A2(n605), .ZN(n607) );
  NOR2_X1 U680 ( .A1(n608), .A2(n607), .ZN(n609) );
  XOR2_X1 U681 ( .A(KEYINPUT15), .B(n609), .Z(n849) );
  INV_X1 U682 ( .A(n849), .ZN(n944) );
  INV_X1 U683 ( .A(G868), .ZN(n681) );
  NAND2_X1 U684 ( .A1(n944), .A2(n681), .ZN(n610) );
  NAND2_X1 U685 ( .A1(n611), .A2(n610), .ZN(G284) );
  NOR2_X1 U686 ( .A1(G286), .A2(n681), .ZN(n613) );
  NOR2_X1 U687 ( .A1(G868), .A2(G299), .ZN(n612) );
  NOR2_X1 U688 ( .A1(n613), .A2(n612), .ZN(G297) );
  INV_X1 U689 ( .A(G860), .ZN(n614) );
  NAND2_X1 U690 ( .A1(G559), .A2(n614), .ZN(n615) );
  XNOR2_X1 U691 ( .A(KEYINPUT76), .B(n615), .ZN(n616) );
  NAND2_X1 U692 ( .A1(n616), .A2(n849), .ZN(n617) );
  XNOR2_X1 U693 ( .A(KEYINPUT16), .B(n617), .ZN(G148) );
  NOR2_X1 U694 ( .A1(G559), .A2(n681), .ZN(n618) );
  NAND2_X1 U695 ( .A1(n849), .A2(n618), .ZN(n619) );
  XNOR2_X1 U696 ( .A(n619), .B(KEYINPUT77), .ZN(n621) );
  INV_X1 U697 ( .A(n934), .ZN(n633) );
  NOR2_X1 U698 ( .A1(n633), .A2(G868), .ZN(n620) );
  NOR2_X1 U699 ( .A1(n621), .A2(n620), .ZN(G282) );
  XNOR2_X1 U700 ( .A(G2100), .B(KEYINPUT79), .ZN(n631) );
  NAND2_X1 U701 ( .A1(G99), .A2(n898), .ZN(n623) );
  NAND2_X1 U702 ( .A1(G111), .A2(n903), .ZN(n622) );
  NAND2_X1 U703 ( .A1(n623), .A2(n622), .ZN(n624) );
  XNOR2_X1 U704 ( .A(KEYINPUT78), .B(n624), .ZN(n629) );
  NAND2_X1 U705 ( .A1(n906), .A2(G123), .ZN(n625) );
  XNOR2_X1 U706 ( .A(n625), .B(KEYINPUT18), .ZN(n627) );
  NAND2_X1 U707 ( .A1(G135), .A2(n899), .ZN(n626) );
  NAND2_X1 U708 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U709 ( .A1(n629), .A2(n628), .ZN(n1008) );
  XNOR2_X1 U710 ( .A(n1008), .B(G2096), .ZN(n630) );
  NAND2_X1 U711 ( .A1(n631), .A2(n630), .ZN(n632) );
  XNOR2_X1 U712 ( .A(KEYINPUT80), .B(n632), .ZN(G156) );
  NAND2_X1 U713 ( .A1(G559), .A2(n849), .ZN(n634) );
  XNOR2_X1 U714 ( .A(n634), .B(n633), .ZN(n677) );
  NOR2_X1 U715 ( .A1(n677), .A2(G860), .ZN(n643) );
  NAND2_X1 U716 ( .A1(G80), .A2(n652), .ZN(n636) );
  NAND2_X1 U717 ( .A1(G93), .A2(n655), .ZN(n635) );
  NAND2_X1 U718 ( .A1(n636), .A2(n635), .ZN(n639) );
  NAND2_X1 U719 ( .A1(G55), .A2(n667), .ZN(n637) );
  XNOR2_X1 U720 ( .A(KEYINPUT81), .B(n637), .ZN(n638) );
  NOR2_X1 U721 ( .A1(n639), .A2(n638), .ZN(n641) );
  NAND2_X1 U722 ( .A1(G67), .A2(n666), .ZN(n640) );
  NAND2_X1 U723 ( .A1(n641), .A2(n640), .ZN(n680) );
  XOR2_X1 U724 ( .A(n680), .B(KEYINPUT82), .Z(n642) );
  XNOR2_X1 U725 ( .A(n643), .B(n642), .ZN(G145) );
  NAND2_X1 U726 ( .A1(G61), .A2(n666), .ZN(n645) );
  NAND2_X1 U727 ( .A1(G86), .A2(n655), .ZN(n644) );
  NAND2_X1 U728 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U729 ( .A(KEYINPUT84), .B(n646), .ZN(n649) );
  NAND2_X1 U730 ( .A1(n652), .A2(G73), .ZN(n647) );
  XOR2_X1 U731 ( .A(KEYINPUT2), .B(n647), .Z(n648) );
  NOR2_X1 U732 ( .A1(n649), .A2(n648), .ZN(n651) );
  NAND2_X1 U733 ( .A1(n667), .A2(G48), .ZN(n650) );
  NAND2_X1 U734 ( .A1(n651), .A2(n650), .ZN(G305) );
  NAND2_X1 U735 ( .A1(n652), .A2(G72), .ZN(n654) );
  NAND2_X1 U736 ( .A1(G60), .A2(n666), .ZN(n653) );
  NAND2_X1 U737 ( .A1(n654), .A2(n653), .ZN(n658) );
  NAND2_X1 U738 ( .A1(G85), .A2(n655), .ZN(n656) );
  XNOR2_X1 U739 ( .A(KEYINPUT67), .B(n656), .ZN(n657) );
  NOR2_X1 U740 ( .A1(n658), .A2(n657), .ZN(n661) );
  NAND2_X1 U741 ( .A1(G47), .A2(n667), .ZN(n659) );
  XOR2_X1 U742 ( .A(KEYINPUT69), .B(n659), .Z(n660) );
  NAND2_X1 U743 ( .A1(n661), .A2(n660), .ZN(G290) );
  NAND2_X1 U744 ( .A1(G87), .A2(n662), .ZN(n664) );
  NAND2_X1 U745 ( .A1(G74), .A2(G651), .ZN(n663) );
  NAND2_X1 U746 ( .A1(n664), .A2(n663), .ZN(n665) );
  NOR2_X1 U747 ( .A1(n666), .A2(n665), .ZN(n670) );
  NAND2_X1 U748 ( .A1(G49), .A2(n667), .ZN(n668) );
  XOR2_X1 U749 ( .A(KEYINPUT83), .B(n668), .Z(n669) );
  NAND2_X1 U750 ( .A1(n670), .A2(n669), .ZN(G288) );
  XNOR2_X1 U751 ( .A(KEYINPUT85), .B(KEYINPUT19), .ZN(n672) );
  XNOR2_X1 U752 ( .A(G305), .B(G166), .ZN(n671) );
  XNOR2_X1 U753 ( .A(n672), .B(n671), .ZN(n673) );
  XNOR2_X1 U754 ( .A(n673), .B(G290), .ZN(n674) );
  XNOR2_X1 U755 ( .A(n674), .B(n680), .ZN(n675) );
  XNOR2_X1 U756 ( .A(n675), .B(G299), .ZN(n676) );
  XNOR2_X1 U757 ( .A(n676), .B(G288), .ZN(n848) );
  XOR2_X1 U758 ( .A(n848), .B(n677), .Z(n678) );
  NAND2_X1 U759 ( .A1(n678), .A2(G868), .ZN(n679) );
  XNOR2_X1 U760 ( .A(n679), .B(KEYINPUT86), .ZN(n683) );
  NAND2_X1 U761 ( .A1(n681), .A2(n680), .ZN(n682) );
  NAND2_X1 U762 ( .A1(n683), .A2(n682), .ZN(G295) );
  NAND2_X1 U763 ( .A1(G2078), .A2(G2084), .ZN(n684) );
  XOR2_X1 U764 ( .A(KEYINPUT20), .B(n684), .Z(n685) );
  NAND2_X1 U765 ( .A1(G2090), .A2(n685), .ZN(n686) );
  XNOR2_X1 U766 ( .A(KEYINPUT21), .B(n686), .ZN(n687) );
  NAND2_X1 U767 ( .A1(n687), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U768 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U769 ( .A1(G220), .A2(G219), .ZN(n688) );
  XOR2_X1 U770 ( .A(KEYINPUT22), .B(n688), .Z(n689) );
  NOR2_X1 U771 ( .A1(G218), .A2(n689), .ZN(n690) );
  NAND2_X1 U772 ( .A1(G96), .A2(n690), .ZN(n846) );
  NAND2_X1 U773 ( .A1(n846), .A2(G2106), .ZN(n694) );
  NAND2_X1 U774 ( .A1(G69), .A2(G120), .ZN(n691) );
  NOR2_X1 U775 ( .A1(G237), .A2(n691), .ZN(n692) );
  NAND2_X1 U776 ( .A1(G108), .A2(n692), .ZN(n847) );
  NAND2_X1 U777 ( .A1(n847), .A2(G567), .ZN(n693) );
  NAND2_X1 U778 ( .A1(n694), .A2(n693), .ZN(n922) );
  NAND2_X1 U779 ( .A1(G661), .A2(G483), .ZN(n695) );
  NOR2_X1 U780 ( .A1(n922), .A2(n695), .ZN(n845) );
  NAND2_X1 U781 ( .A1(n845), .A2(G36), .ZN(G176) );
  INV_X1 U782 ( .A(G166), .ZN(G303) );
  INV_X1 U783 ( .A(n746), .ZN(n728) );
  NAND2_X1 U784 ( .A1(G1996), .A2(n728), .ZN(n698) );
  XNOR2_X1 U785 ( .A(KEYINPUT26), .B(n698), .ZN(n699) );
  NAND2_X1 U786 ( .A1(n699), .A2(n934), .ZN(n702) );
  NAND2_X1 U787 ( .A1(G1341), .A2(n746), .ZN(n700) );
  XNOR2_X1 U788 ( .A(KEYINPUT95), .B(n700), .ZN(n701) );
  NOR2_X1 U789 ( .A1(n702), .A2(n701), .ZN(n707) );
  NAND2_X1 U790 ( .A1(n849), .A2(n707), .ZN(n706) );
  XOR2_X1 U791 ( .A(KEYINPUT93), .B(n746), .Z(n712) );
  INV_X1 U792 ( .A(n712), .ZN(n710) );
  NAND2_X1 U793 ( .A1(G2067), .A2(n710), .ZN(n704) );
  NAND2_X1 U794 ( .A1(G1348), .A2(n746), .ZN(n703) );
  NAND2_X1 U795 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U796 ( .A1(n706), .A2(n705), .ZN(n709) );
  OR2_X1 U797 ( .A1(n849), .A2(n707), .ZN(n708) );
  NAND2_X1 U798 ( .A1(n709), .A2(n708), .ZN(n718) );
  NAND2_X1 U799 ( .A1(n710), .A2(G2072), .ZN(n711) );
  XOR2_X1 U800 ( .A(n711), .B(KEYINPUT27), .Z(n720) );
  NAND2_X1 U801 ( .A1(G1956), .A2(n712), .ZN(n719) );
  INV_X1 U802 ( .A(G299), .ZN(n713) );
  AND2_X1 U803 ( .A1(n719), .A2(n713), .ZN(n714) );
  AND2_X1 U804 ( .A1(n720), .A2(n714), .ZN(n716) );
  XNOR2_X1 U805 ( .A(n716), .B(n715), .ZN(n717) );
  NAND2_X1 U806 ( .A1(n718), .A2(n717), .ZN(n724) );
  NAND2_X1 U807 ( .A1(n720), .A2(n719), .ZN(n721) );
  NAND2_X1 U808 ( .A1(G299), .A2(n721), .ZN(n722) );
  XNOR2_X1 U809 ( .A(n722), .B(KEYINPUT28), .ZN(n723) );
  NAND2_X1 U810 ( .A1(n724), .A2(n723), .ZN(n726) );
  XNOR2_X1 U811 ( .A(G2078), .B(KEYINPUT25), .ZN(n727) );
  XNOR2_X1 U812 ( .A(n727), .B(KEYINPUT94), .ZN(n955) );
  NAND2_X1 U813 ( .A1(n710), .A2(n955), .ZN(n730) );
  OR2_X1 U814 ( .A1(G1961), .A2(n728), .ZN(n729) );
  NAND2_X1 U815 ( .A1(n730), .A2(n729), .ZN(n738) );
  NAND2_X1 U816 ( .A1(n738), .A2(G171), .ZN(n731) );
  NAND2_X1 U817 ( .A1(n732), .A2(n731), .ZN(n743) );
  NAND2_X1 U818 ( .A1(G8), .A2(n746), .ZN(n778) );
  NOR2_X1 U819 ( .A1(G1966), .A2(n778), .ZN(n758) );
  NOR2_X1 U820 ( .A1(n746), .A2(G2084), .ZN(n733) );
  XNOR2_X1 U821 ( .A(n733), .B(KEYINPUT92), .ZN(n755) );
  NOR2_X1 U822 ( .A1(n758), .A2(n755), .ZN(n734) );
  NAND2_X1 U823 ( .A1(n734), .A2(G8), .ZN(n735) );
  XOR2_X1 U824 ( .A(KEYINPUT30), .B(n735), .Z(n736) );
  XNOR2_X1 U825 ( .A(KEYINPUT97), .B(n736), .ZN(n737) );
  NOR2_X1 U826 ( .A1(G168), .A2(n737), .ZN(n740) );
  NOR2_X1 U827 ( .A1(G171), .A2(n738), .ZN(n739) );
  NOR2_X1 U828 ( .A1(n740), .A2(n739), .ZN(n741) );
  XOR2_X1 U829 ( .A(KEYINPUT31), .B(n741), .Z(n742) );
  NAND2_X1 U830 ( .A1(n743), .A2(n742), .ZN(n744) );
  XNOR2_X1 U831 ( .A(n744), .B(KEYINPUT98), .ZN(n756) );
  AND2_X1 U832 ( .A1(n756), .A2(G286), .ZN(n753) );
  INV_X1 U833 ( .A(G8), .ZN(n751) );
  NOR2_X1 U834 ( .A1(G1971), .A2(n778), .ZN(n745) );
  XNOR2_X1 U835 ( .A(KEYINPUT99), .B(n745), .ZN(n749) );
  NOR2_X1 U836 ( .A1(G2090), .A2(n746), .ZN(n747) );
  NOR2_X1 U837 ( .A1(G166), .A2(n747), .ZN(n748) );
  NAND2_X1 U838 ( .A1(n749), .A2(n748), .ZN(n750) );
  NOR2_X1 U839 ( .A1(n751), .A2(n750), .ZN(n752) );
  NOR2_X1 U840 ( .A1(n753), .A2(n752), .ZN(n754) );
  XNOR2_X1 U841 ( .A(n754), .B(KEYINPUT32), .ZN(n762) );
  NAND2_X1 U842 ( .A1(n755), .A2(G8), .ZN(n760) );
  INV_X1 U843 ( .A(n756), .ZN(n757) );
  NOR2_X1 U844 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U845 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U846 ( .A1(n762), .A2(n761), .ZN(n776) );
  NOR2_X1 U847 ( .A1(G1976), .A2(G288), .ZN(n923) );
  NOR2_X1 U848 ( .A1(G1971), .A2(G303), .ZN(n763) );
  NOR2_X1 U849 ( .A1(n923), .A2(n763), .ZN(n765) );
  INV_X1 U850 ( .A(KEYINPUT33), .ZN(n764) );
  AND2_X1 U851 ( .A1(n765), .A2(n764), .ZN(n766) );
  NAND2_X1 U852 ( .A1(n776), .A2(n766), .ZN(n772) );
  INV_X1 U853 ( .A(n778), .ZN(n784) );
  NAND2_X1 U854 ( .A1(G1976), .A2(G288), .ZN(n924) );
  AND2_X1 U855 ( .A1(n784), .A2(n924), .ZN(n767) );
  NOR2_X1 U856 ( .A1(KEYINPUT33), .A2(n767), .ZN(n770) );
  NAND2_X1 U857 ( .A1(n923), .A2(KEYINPUT33), .ZN(n768) );
  NOR2_X1 U858 ( .A1(n768), .A2(n778), .ZN(n769) );
  NOR2_X1 U859 ( .A1(n770), .A2(n769), .ZN(n771) );
  AND2_X1 U860 ( .A1(n772), .A2(n771), .ZN(n773) );
  XOR2_X1 U861 ( .A(G1981), .B(G305), .Z(n939) );
  NAND2_X1 U862 ( .A1(n773), .A2(n939), .ZN(n781) );
  NOR2_X1 U863 ( .A1(G2090), .A2(G303), .ZN(n774) );
  XNOR2_X1 U864 ( .A(n774), .B(KEYINPUT100), .ZN(n775) );
  NAND2_X1 U865 ( .A1(n775), .A2(G8), .ZN(n777) );
  NAND2_X1 U866 ( .A1(n777), .A2(n776), .ZN(n779) );
  NAND2_X1 U867 ( .A1(n779), .A2(n778), .ZN(n780) );
  NAND2_X1 U868 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U869 ( .A(n782), .B(KEYINPUT101), .ZN(n787) );
  NOR2_X1 U870 ( .A1(G1981), .A2(G305), .ZN(n783) );
  XNOR2_X1 U871 ( .A(n783), .B(KEYINPUT24), .ZN(n785) );
  NAND2_X1 U872 ( .A1(n785), .A2(n784), .ZN(n786) );
  AND2_X1 U873 ( .A1(n787), .A2(n786), .ZN(n820) );
  INV_X1 U874 ( .A(n788), .ZN(n789) );
  NOR2_X1 U875 ( .A1(n790), .A2(n789), .ZN(n835) );
  NAND2_X1 U876 ( .A1(G95), .A2(n898), .ZN(n792) );
  NAND2_X1 U877 ( .A1(G131), .A2(n899), .ZN(n791) );
  NAND2_X1 U878 ( .A1(n792), .A2(n791), .ZN(n796) );
  NAND2_X1 U879 ( .A1(G119), .A2(n906), .ZN(n794) );
  NAND2_X1 U880 ( .A1(G107), .A2(n903), .ZN(n793) );
  NAND2_X1 U881 ( .A1(n794), .A2(n793), .ZN(n795) );
  OR2_X1 U882 ( .A1(n796), .A2(n795), .ZN(n881) );
  AND2_X1 U883 ( .A1(n881), .A2(G1991), .ZN(n1007) );
  NAND2_X1 U884 ( .A1(G129), .A2(n906), .ZN(n798) );
  NAND2_X1 U885 ( .A1(G117), .A2(n903), .ZN(n797) );
  NAND2_X1 U886 ( .A1(n798), .A2(n797), .ZN(n801) );
  NAND2_X1 U887 ( .A1(n898), .A2(G105), .ZN(n799) );
  XOR2_X1 U888 ( .A(KEYINPUT38), .B(n799), .Z(n800) );
  NOR2_X1 U889 ( .A1(n801), .A2(n800), .ZN(n803) );
  NAND2_X1 U890 ( .A1(G141), .A2(n899), .ZN(n802) );
  NAND2_X1 U891 ( .A1(n803), .A2(n802), .ZN(n895) );
  AND2_X1 U892 ( .A1(n895), .A2(G1996), .ZN(n1009) );
  OR2_X1 U893 ( .A1(n1007), .A2(n1009), .ZN(n804) );
  NAND2_X1 U894 ( .A1(n835), .A2(n804), .ZN(n823) );
  XNOR2_X1 U895 ( .A(KEYINPUT89), .B(KEYINPUT36), .ZN(n815) );
  NAND2_X1 U896 ( .A1(G128), .A2(n906), .ZN(n806) );
  NAND2_X1 U897 ( .A1(G116), .A2(n903), .ZN(n805) );
  NAND2_X1 U898 ( .A1(n806), .A2(n805), .ZN(n807) );
  XNOR2_X1 U899 ( .A(KEYINPUT35), .B(n807), .ZN(n813) );
  NAND2_X1 U900 ( .A1(G104), .A2(n898), .ZN(n809) );
  NAND2_X1 U901 ( .A1(G140), .A2(n899), .ZN(n808) );
  NAND2_X1 U902 ( .A1(n809), .A2(n808), .ZN(n811) );
  XOR2_X1 U903 ( .A(KEYINPUT88), .B(KEYINPUT34), .Z(n810) );
  XNOR2_X1 U904 ( .A(n811), .B(n810), .ZN(n812) );
  NAND2_X1 U905 ( .A1(n813), .A2(n812), .ZN(n814) );
  XNOR2_X1 U906 ( .A(n815), .B(n814), .ZN(n882) );
  XNOR2_X1 U907 ( .A(KEYINPUT37), .B(G2067), .ZN(n833) );
  NOR2_X1 U908 ( .A1(n882), .A2(n833), .ZN(n816) );
  XNOR2_X1 U909 ( .A(n816), .B(KEYINPUT90), .ZN(n1026) );
  NAND2_X1 U910 ( .A1(n1026), .A2(n835), .ZN(n817) );
  XNOR2_X1 U911 ( .A(n817), .B(KEYINPUT91), .ZN(n831) );
  INV_X1 U912 ( .A(n831), .ZN(n818) );
  NAND2_X1 U913 ( .A1(n823), .A2(n818), .ZN(n819) );
  XNOR2_X1 U914 ( .A(G1986), .B(G290), .ZN(n928) );
  NAND2_X1 U915 ( .A1(n928), .A2(n835), .ZN(n821) );
  NAND2_X1 U916 ( .A1(n822), .A2(n821), .ZN(n838) );
  NOR2_X1 U917 ( .A1(G1996), .A2(n895), .ZN(n1003) );
  INV_X1 U918 ( .A(n823), .ZN(n827) );
  NOR2_X1 U919 ( .A1(G1991), .A2(n881), .ZN(n1006) );
  NOR2_X1 U920 ( .A1(G1986), .A2(G290), .ZN(n824) );
  XNOR2_X1 U921 ( .A(KEYINPUT102), .B(n824), .ZN(n825) );
  NOR2_X1 U922 ( .A1(n1006), .A2(n825), .ZN(n826) );
  NOR2_X1 U923 ( .A1(n827), .A2(n826), .ZN(n828) );
  NOR2_X1 U924 ( .A1(n1003), .A2(n828), .ZN(n829) );
  XOR2_X1 U925 ( .A(KEYINPUT39), .B(n829), .Z(n830) );
  NOR2_X1 U926 ( .A1(n831), .A2(n830), .ZN(n832) );
  XNOR2_X1 U927 ( .A(n832), .B(KEYINPUT103), .ZN(n834) );
  NAND2_X1 U928 ( .A1(n833), .A2(n882), .ZN(n1014) );
  NAND2_X1 U929 ( .A1(n834), .A2(n1014), .ZN(n836) );
  NAND2_X1 U930 ( .A1(n836), .A2(n835), .ZN(n837) );
  NAND2_X1 U931 ( .A1(n838), .A2(n837), .ZN(n840) );
  XNOR2_X1 U932 ( .A(KEYINPUT40), .B(KEYINPUT104), .ZN(n839) );
  XNOR2_X1 U933 ( .A(n840), .B(n839), .ZN(G329) );
  NAND2_X1 U934 ( .A1(G2106), .A2(n841), .ZN(G217) );
  NAND2_X1 U935 ( .A1(G15), .A2(G2), .ZN(n842) );
  XNOR2_X1 U936 ( .A(KEYINPUT107), .B(n842), .ZN(n843) );
  NAND2_X1 U937 ( .A1(n843), .A2(G661), .ZN(G259) );
  NAND2_X1 U938 ( .A1(G3), .A2(G1), .ZN(n844) );
  NAND2_X1 U939 ( .A1(n845), .A2(n844), .ZN(G188) );
  NOR2_X1 U940 ( .A1(n847), .A2(n846), .ZN(G325) );
  XOR2_X1 U941 ( .A(KEYINPUT108), .B(G325), .Z(G261) );
  INV_X1 U943 ( .A(G120), .ZN(G236) );
  INV_X1 U944 ( .A(G96), .ZN(G221) );
  INV_X1 U945 ( .A(G69), .ZN(G235) );
  XOR2_X1 U946 ( .A(n848), .B(G286), .Z(n851) );
  XNOR2_X1 U947 ( .A(G171), .B(n849), .ZN(n850) );
  XNOR2_X1 U948 ( .A(n851), .B(n850), .ZN(n852) );
  XNOR2_X1 U949 ( .A(n852), .B(n934), .ZN(n853) );
  NOR2_X1 U950 ( .A1(G37), .A2(n853), .ZN(G397) );
  XOR2_X1 U951 ( .A(G2096), .B(G2100), .Z(n855) );
  XNOR2_X1 U952 ( .A(KEYINPUT42), .B(G2678), .ZN(n854) );
  XNOR2_X1 U953 ( .A(n855), .B(n854), .ZN(n859) );
  XOR2_X1 U954 ( .A(KEYINPUT43), .B(G2072), .Z(n857) );
  XNOR2_X1 U955 ( .A(G2067), .B(G2090), .ZN(n856) );
  XNOR2_X1 U956 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U957 ( .A(n859), .B(n858), .Z(n861) );
  XNOR2_X1 U958 ( .A(G2078), .B(G2084), .ZN(n860) );
  XNOR2_X1 U959 ( .A(n861), .B(n860), .ZN(G227) );
  XOR2_X1 U960 ( .A(G1976), .B(G1971), .Z(n863) );
  XNOR2_X1 U961 ( .A(G1986), .B(G1956), .ZN(n862) );
  XNOR2_X1 U962 ( .A(n863), .B(n862), .ZN(n864) );
  XOR2_X1 U963 ( .A(n864), .B(KEYINPUT41), .Z(n866) );
  XNOR2_X1 U964 ( .A(G1996), .B(G1991), .ZN(n865) );
  XNOR2_X1 U965 ( .A(n866), .B(n865), .ZN(n870) );
  XOR2_X1 U966 ( .A(G2474), .B(G1961), .Z(n868) );
  XNOR2_X1 U967 ( .A(G1981), .B(G1966), .ZN(n867) );
  XNOR2_X1 U968 ( .A(n868), .B(n867), .ZN(n869) );
  XNOR2_X1 U969 ( .A(n870), .B(n869), .ZN(G229) );
  NAND2_X1 U970 ( .A1(n906), .A2(G124), .ZN(n871) );
  XNOR2_X1 U971 ( .A(n871), .B(KEYINPUT44), .ZN(n873) );
  NAND2_X1 U972 ( .A1(G136), .A2(n899), .ZN(n872) );
  NAND2_X1 U973 ( .A1(n873), .A2(n872), .ZN(n874) );
  XNOR2_X1 U974 ( .A(n874), .B(KEYINPUT109), .ZN(n876) );
  NAND2_X1 U975 ( .A1(G112), .A2(n903), .ZN(n875) );
  NAND2_X1 U976 ( .A1(n876), .A2(n875), .ZN(n879) );
  NAND2_X1 U977 ( .A1(n898), .A2(G100), .ZN(n877) );
  XOR2_X1 U978 ( .A(KEYINPUT110), .B(n877), .Z(n878) );
  NOR2_X1 U979 ( .A1(n879), .A2(n878), .ZN(n880) );
  XOR2_X1 U980 ( .A(KEYINPUT111), .B(n880), .Z(G162) );
  XNOR2_X1 U981 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n884) );
  XOR2_X1 U982 ( .A(n882), .B(n881), .Z(n883) );
  XNOR2_X1 U983 ( .A(n884), .B(n883), .ZN(n894) );
  NAND2_X1 U984 ( .A1(G127), .A2(n906), .ZN(n886) );
  NAND2_X1 U985 ( .A1(G115), .A2(n903), .ZN(n885) );
  NAND2_X1 U986 ( .A1(n886), .A2(n885), .ZN(n887) );
  XNOR2_X1 U987 ( .A(n887), .B(KEYINPUT47), .ZN(n892) );
  NAND2_X1 U988 ( .A1(G103), .A2(n898), .ZN(n889) );
  NAND2_X1 U989 ( .A1(G139), .A2(n899), .ZN(n888) );
  NAND2_X1 U990 ( .A1(n889), .A2(n888), .ZN(n890) );
  XNOR2_X1 U991 ( .A(KEYINPUT113), .B(n890), .ZN(n891) );
  NAND2_X1 U992 ( .A1(n892), .A2(n891), .ZN(n893) );
  XNOR2_X1 U993 ( .A(n893), .B(KEYINPUT114), .ZN(n1016) );
  XOR2_X1 U994 ( .A(n894), .B(n1016), .Z(n897) );
  XOR2_X1 U995 ( .A(G160), .B(n895), .Z(n896) );
  XNOR2_X1 U996 ( .A(n897), .B(n896), .ZN(n911) );
  NAND2_X1 U997 ( .A1(G106), .A2(n898), .ZN(n901) );
  NAND2_X1 U998 ( .A1(G142), .A2(n899), .ZN(n900) );
  NAND2_X1 U999 ( .A1(n901), .A2(n900), .ZN(n902) );
  XNOR2_X1 U1000 ( .A(n902), .B(KEYINPUT45), .ZN(n905) );
  NAND2_X1 U1001 ( .A1(G118), .A2(n903), .ZN(n904) );
  NAND2_X1 U1002 ( .A1(n905), .A2(n904), .ZN(n909) );
  NAND2_X1 U1003 ( .A1(n906), .A2(G130), .ZN(n907) );
  XOR2_X1 U1004 ( .A(KEYINPUT112), .B(n907), .Z(n908) );
  NOR2_X1 U1005 ( .A1(n909), .A2(n908), .ZN(n910) );
  XOR2_X1 U1006 ( .A(n911), .B(n910), .Z(n913) );
  XNOR2_X1 U1007 ( .A(G164), .B(n1008), .ZN(n912) );
  XNOR2_X1 U1008 ( .A(n913), .B(n912), .ZN(n914) );
  XOR2_X1 U1009 ( .A(G162), .B(n914), .Z(n915) );
  NOR2_X1 U1010 ( .A1(G37), .A2(n915), .ZN(G395) );
  NOR2_X1 U1011 ( .A1(G401), .A2(n922), .ZN(n919) );
  NOR2_X1 U1012 ( .A1(G227), .A2(G229), .ZN(n916) );
  XNOR2_X1 U1013 ( .A(KEYINPUT49), .B(n916), .ZN(n917) );
  NOR2_X1 U1014 ( .A1(G397), .A2(n917), .ZN(n918) );
  NAND2_X1 U1015 ( .A1(n919), .A2(n918), .ZN(n920) );
  NOR2_X1 U1016 ( .A1(n920), .A2(G395), .ZN(n921) );
  XNOR2_X1 U1017 ( .A(n921), .B(KEYINPUT115), .ZN(G225) );
  INV_X1 U1018 ( .A(G225), .ZN(G308) );
  INV_X1 U1019 ( .A(n922), .ZN(G319) );
  INV_X1 U1020 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1021 ( .A(G166), .B(G1971), .ZN(n930) );
  INV_X1 U1022 ( .A(n923), .ZN(n925) );
  NAND2_X1 U1023 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1024 ( .A(KEYINPUT122), .B(n926), .ZN(n927) );
  NOR2_X1 U1025 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1026 ( .A1(n930), .A2(n929), .ZN(n932) );
  XNOR2_X1 U1027 ( .A(G1956), .B(G299), .ZN(n931) );
  NOR2_X1 U1028 ( .A1(n932), .A2(n931), .ZN(n933) );
  XOR2_X1 U1029 ( .A(KEYINPUT123), .B(n933), .Z(n936) );
  XNOR2_X1 U1030 ( .A(n934), .B(G1341), .ZN(n935) );
  NAND2_X1 U1031 ( .A1(n936), .A2(n935), .ZN(n943) );
  XOR2_X1 U1032 ( .A(KEYINPUT57), .B(KEYINPUT121), .Z(n941) );
  XNOR2_X1 U1033 ( .A(G1966), .B(G168), .ZN(n937) );
  XNOR2_X1 U1034 ( .A(n937), .B(KEYINPUT120), .ZN(n938) );
  NAND2_X1 U1035 ( .A1(n939), .A2(n938), .ZN(n940) );
  XOR2_X1 U1036 ( .A(n941), .B(n940), .Z(n942) );
  NOR2_X1 U1037 ( .A1(n943), .A2(n942), .ZN(n948) );
  XOR2_X1 U1038 ( .A(G171), .B(G1961), .Z(n946) );
  XNOR2_X1 U1039 ( .A(n944), .B(G1348), .ZN(n945) );
  NOR2_X1 U1040 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1041 ( .A1(n948), .A2(n947), .ZN(n951) );
  XOR2_X1 U1042 ( .A(G16), .B(KEYINPUT56), .Z(n949) );
  XNOR2_X1 U1043 ( .A(KEYINPUT119), .B(n949), .ZN(n950) );
  NAND2_X1 U1044 ( .A1(n951), .A2(n950), .ZN(n1000) );
  XNOR2_X1 U1045 ( .A(G2067), .B(G26), .ZN(n953) );
  XNOR2_X1 U1046 ( .A(G33), .B(G2072), .ZN(n952) );
  NOR2_X1 U1047 ( .A1(n953), .A2(n952), .ZN(n961) );
  XOR2_X1 U1048 ( .A(G32), .B(G1996), .Z(n954) );
  NAND2_X1 U1049 ( .A1(n954), .A2(G28), .ZN(n959) );
  XNOR2_X1 U1050 ( .A(G27), .B(n955), .ZN(n957) );
  XOR2_X1 U1051 ( .A(G1991), .B(G25), .Z(n956) );
  NAND2_X1 U1052 ( .A1(n957), .A2(n956), .ZN(n958) );
  NOR2_X1 U1053 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1054 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1055 ( .A(n962), .B(KEYINPUT53), .ZN(n965) );
  XOR2_X1 U1056 ( .A(G2084), .B(G34), .Z(n963) );
  XNOR2_X1 U1057 ( .A(KEYINPUT54), .B(n963), .ZN(n964) );
  NAND2_X1 U1058 ( .A1(n965), .A2(n964), .ZN(n967) );
  XNOR2_X1 U1059 ( .A(G35), .B(G2090), .ZN(n966) );
  NOR2_X1 U1060 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1061 ( .A(KEYINPUT55), .B(n968), .ZN(n970) );
  INV_X1 U1062 ( .A(G29), .ZN(n969) );
  NAND2_X1 U1063 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1064 ( .A1(n971), .A2(G11), .ZN(n972) );
  XNOR2_X1 U1065 ( .A(KEYINPUT118), .B(n972), .ZN(n998) );
  XOR2_X1 U1066 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n994) );
  XNOR2_X1 U1067 ( .A(G1981), .B(G6), .ZN(n974) );
  XNOR2_X1 U1068 ( .A(G1341), .B(G19), .ZN(n973) );
  NOR2_X1 U1069 ( .A1(n974), .A2(n973), .ZN(n980) );
  XOR2_X1 U1070 ( .A(KEYINPUT124), .B(G4), .Z(n976) );
  XNOR2_X1 U1071 ( .A(G1348), .B(KEYINPUT59), .ZN(n975) );
  XNOR2_X1 U1072 ( .A(n976), .B(n975), .ZN(n978) );
  XNOR2_X1 U1073 ( .A(G1956), .B(G20), .ZN(n977) );
  NOR2_X1 U1074 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1075 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1076 ( .A(n981), .B(KEYINPUT60), .ZN(n988) );
  XNOR2_X1 U1077 ( .A(G1971), .B(G22), .ZN(n983) );
  XNOR2_X1 U1078 ( .A(G23), .B(G1976), .ZN(n982) );
  NOR2_X1 U1079 ( .A1(n983), .A2(n982), .ZN(n985) );
  XOR2_X1 U1080 ( .A(G1986), .B(G24), .Z(n984) );
  NAND2_X1 U1081 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1082 ( .A(KEYINPUT58), .B(n986), .ZN(n987) );
  NOR2_X1 U1083 ( .A1(n988), .A2(n987), .ZN(n992) );
  XNOR2_X1 U1084 ( .A(G1966), .B(G21), .ZN(n990) );
  XNOR2_X1 U1085 ( .A(G5), .B(G1961), .ZN(n989) );
  NOR2_X1 U1086 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1087 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1088 ( .A(n994), .B(n993), .ZN(n995) );
  NOR2_X1 U1089 ( .A1(G16), .A2(n995), .ZN(n996) );
  XNOR2_X1 U1090 ( .A(n996), .B(KEYINPUT126), .ZN(n997) );
  NOR2_X1 U1091 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1092 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1093 ( .A(n1001), .B(KEYINPUT127), .ZN(n1032) );
  XOR2_X1 U1094 ( .A(G2090), .B(G162), .Z(n1002) );
  NOR2_X1 U1095 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XOR2_X1 U1096 ( .A(KEYINPUT116), .B(n1004), .Z(n1005) );
  XNOR2_X1 U1097 ( .A(KEYINPUT51), .B(n1005), .ZN(n1024) );
  NOR2_X1 U1098 ( .A1(n1007), .A2(n1006), .ZN(n1011) );
  NOR2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1013) );
  XOR2_X1 U1101 ( .A(G160), .B(G2084), .Z(n1012) );
  NOR2_X1 U1102 ( .A1(n1013), .A2(n1012), .ZN(n1015) );
  NAND2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1022) );
  XOR2_X1 U1104 ( .A(G2072), .B(n1016), .Z(n1018) );
  XNOR2_X1 U1105 ( .A(G164), .B(G2078), .ZN(n1017) );
  NAND2_X1 U1106 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XOR2_X1 U1107 ( .A(KEYINPUT117), .B(n1019), .Z(n1020) );
  XNOR2_X1 U1108 ( .A(KEYINPUT50), .B(n1020), .ZN(n1021) );
  NOR2_X1 U1109 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1110 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NOR2_X1 U1111 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1112 ( .A(KEYINPUT52), .B(n1027), .ZN(n1029) );
  INV_X1 U1113 ( .A(KEYINPUT55), .ZN(n1028) );
  NAND2_X1 U1114 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NAND2_X1 U1115 ( .A1(n1030), .A2(G29), .ZN(n1031) );
  NAND2_X1 U1116 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XOR2_X1 U1117 ( .A(KEYINPUT62), .B(n1033), .Z(G311) );
  INV_X1 U1118 ( .A(G311), .ZN(G150) );
endmodule

