//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 1 1 0 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 0 1 0 1 1 0 0 1 1 1 1 0 0 0 0 1 1 1 0 1 1 0 0 1 1 0 0 1 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n653, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n673, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n713, new_n714, new_n716,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n819, new_n820, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n868, new_n869, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n884,
    new_n885, new_n886, new_n887, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929;
  NOR2_X1   g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT64), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n204), .B1(G169gat), .B2(G176gat), .ZN(new_n205));
  AOI21_X1  g004(.A(KEYINPUT26), .B1(new_n203), .B2(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(G169gat), .A2(G176gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT26), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n207), .B1(new_n202), .B2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G183gat), .ZN(new_n210));
  INV_X1    g009(.A(G190gat), .ZN(new_n211));
  OAI22_X1  g010(.A1(new_n206), .A2(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n210), .A2(KEYINPUT27), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n210), .A2(KEYINPUT27), .ZN(new_n215));
  AND4_X1   g014(.A1(KEYINPUT28), .A2(new_n214), .A3(new_n215), .A4(new_n211), .ZN(new_n216));
  AOI21_X1  g015(.A(G190gat), .B1(new_n213), .B2(KEYINPUT69), .ZN(new_n217));
  NAND2_X1  g016(.A1(KEYINPUT69), .A2(G183gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT68), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n218), .A2(new_n219), .A3(KEYINPUT27), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT27), .ZN(new_n221));
  OAI21_X1  g020(.A(KEYINPUT68), .B1(new_n221), .B2(G183gat), .ZN(new_n222));
  NAND4_X1  g021(.A1(new_n217), .A2(KEYINPUT70), .A3(new_n220), .A4(new_n222), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n221), .A2(KEYINPUT69), .A3(G183gat), .ZN(new_n224));
  NAND4_X1  g023(.A1(new_n220), .A2(new_n222), .A3(new_n211), .A4(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT70), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT28), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n223), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n216), .B1(new_n229), .B2(KEYINPUT71), .ZN(new_n230));
  AOI21_X1  g029(.A(KEYINPUT28), .B1(new_n225), .B2(new_n226), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT71), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n231), .A2(new_n232), .A3(new_n223), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n212), .B1(new_n230), .B2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT65), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT23), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n236), .B1(new_n203), .B2(new_n205), .ZN(new_n237));
  INV_X1    g036(.A(new_n207), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n235), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT67), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n210), .A2(new_n211), .ZN(new_n241));
  NAND3_X1  g040(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n242));
  AOI21_X1  g041(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT66), .ZN(new_n244));
  OAI211_X1 g043(.A(new_n241), .B(new_n242), .C1(new_n243), .C2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n243), .A2(new_n244), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n240), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n243), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(KEYINPUT66), .ZN(new_n250));
  AND2_X1   g049(.A1(new_n241), .A2(new_n242), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n250), .A2(new_n251), .A3(KEYINPUT67), .A4(new_n246), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n239), .A2(new_n248), .A3(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n236), .B1(G169gat), .B2(G176gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(KEYINPUT25), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n237), .A2(new_n238), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n256), .B1(new_n257), .B2(KEYINPUT65), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT25), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n251), .A2(new_n249), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n238), .B1(KEYINPUT23), .B2(new_n202), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n260), .A2(new_n255), .A3(new_n261), .ZN(new_n262));
  AOI22_X1  g061(.A1(new_n254), .A2(new_n258), .B1(new_n259), .B2(new_n262), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n234), .A2(new_n263), .ZN(new_n264));
  XOR2_X1   g063(.A(G113gat), .B(G120gat), .Z(new_n265));
  INV_X1    g064(.A(KEYINPUT1), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(G127gat), .B(G134gat), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n265), .A2(new_n266), .A3(new_n268), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(KEYINPUT72), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT72), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n264), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(G227gat), .A2(G233gat), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n277), .B1(new_n234), .B2(new_n263), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(KEYINPUT34), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT34), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n279), .A2(new_n284), .A3(new_n280), .A4(new_n281), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  XOR2_X1   g086(.A(G15gat), .B(G43gat), .Z(new_n288));
  XNOR2_X1  g087(.A(G71gat), .B(G99gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n288), .B(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n280), .B1(new_n279), .B2(new_n281), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n290), .B1(new_n291), .B2(KEYINPUT33), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT32), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  AND2_X1   g093(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n292), .A2(new_n294), .ZN(new_n296));
  OAI211_X1 g095(.A(KEYINPUT73), .B(new_n287), .C1(new_n295), .C2(new_n296), .ZN(new_n297));
  OR2_X1    g096(.A1(new_n292), .A2(new_n294), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT73), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n286), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n283), .A2(KEYINPUT73), .A3(new_n285), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n292), .A2(new_n294), .ZN(new_n302));
  NAND4_X1  g101(.A1(new_n298), .A2(new_n300), .A3(new_n301), .A4(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n297), .A2(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(new_n304), .B(KEYINPUT36), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  OAI21_X1  g105(.A(KEYINPUT76), .B1(new_n234), .B2(new_n263), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT76), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n262), .A2(new_n259), .ZN(new_n309));
  INV_X1    g108(.A(new_n258), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n309), .B1(new_n310), .B2(new_n253), .ZN(new_n311));
  AND3_X1   g110(.A1(new_n231), .A2(new_n232), .A3(new_n223), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n232), .B1(new_n231), .B2(new_n223), .ZN(new_n313));
  NOR3_X1   g112(.A1(new_n312), .A2(new_n313), .A3(new_n216), .ZN(new_n314));
  OAI211_X1 g113(.A(new_n308), .B(new_n311), .C1(new_n314), .C2(new_n212), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n307), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(G226gat), .A2(G233gat), .ZN(new_n317));
  XOR2_X1   g116(.A(new_n317), .B(KEYINPUT75), .Z(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  XOR2_X1   g119(.A(KEYINPUT74), .B(G211gat), .Z(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(G218gat), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT22), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(G197gat), .B(G204gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  XOR2_X1   g125(.A(G211gat), .B(G218gat), .Z(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n327), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n324), .A2(new_n329), .A3(new_n325), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT29), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n332), .B1(new_n234), .B2(new_n263), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(new_n317), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n320), .A2(new_n331), .A3(new_n334), .ZN(new_n335));
  OR2_X1    g134(.A1(new_n264), .A2(new_n317), .ZN(new_n336));
  AOI21_X1  g135(.A(KEYINPUT29), .B1(new_n307), .B2(new_n315), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n336), .B1(new_n337), .B2(new_n319), .ZN(new_n338));
  INV_X1    g137(.A(new_n331), .ZN(new_n339));
  AOI22_X1  g138(.A1(KEYINPUT77), .A2(new_n335), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  AND3_X1   g139(.A1(new_n338), .A2(KEYINPUT77), .A3(new_n339), .ZN(new_n341));
  OAI21_X1  g140(.A(KEYINPUT78), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(G8gat), .B(G36gat), .ZN(new_n343));
  XNOR2_X1  g142(.A(G64gat), .B(G92gat), .ZN(new_n344));
  XNOR2_X1  g143(.A(new_n343), .B(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT78), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n338), .A2(KEYINPUT77), .A3(new_n339), .ZN(new_n347));
  AND2_X1   g146(.A1(new_n338), .A2(new_n339), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT77), .ZN(new_n349));
  AOI22_X1  g148(.A1(new_n316), .A2(new_n319), .B1(new_n317), .B2(new_n333), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n349), .B1(new_n350), .B2(new_n331), .ZN(new_n351));
  OAI211_X1 g150(.A(new_n346), .B(new_n347), .C1(new_n348), .C2(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n342), .A2(new_n345), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(KEYINPUT79), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT79), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n342), .A2(new_n352), .A3(new_n355), .A4(new_n345), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  NOR2_X1   g156(.A1(KEYINPUT80), .A2(KEYINPUT30), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n335), .A2(KEYINPUT77), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n338), .A2(new_n339), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n345), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n361), .A2(new_n362), .A3(new_n347), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n363), .A2(KEYINPUT80), .A3(KEYINPUT30), .ZN(new_n364));
  NAND2_X1  g163(.A1(KEYINPUT80), .A2(KEYINPUT30), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n361), .A2(new_n362), .A3(new_n347), .A4(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n358), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n357), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(G225gat), .A2(G233gat), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  XOR2_X1   g169(.A(G141gat), .B(G148gat), .Z(new_n371));
  XNOR2_X1  g170(.A(G155gat), .B(G162gat), .ZN(new_n372));
  INV_X1    g171(.A(G155gat), .ZN(new_n373));
  INV_X1    g172(.A(G162gat), .ZN(new_n374));
  OAI21_X1  g173(.A(KEYINPUT2), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  AND3_X1   g174(.A1(new_n371), .A2(new_n372), .A3(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n372), .B1(new_n371), .B2(new_n375), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(KEYINPUT4), .B1(new_n278), .B2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n378), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(KEYINPUT3), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n273), .A2(KEYINPUT81), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT81), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n272), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT3), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n378), .A2(new_n385), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n381), .A2(new_n382), .A3(new_n384), .A4(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT4), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n273), .A2(new_n378), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n387), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n370), .B1(new_n379), .B2(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n382), .A2(new_n380), .A3(new_n384), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(new_n389), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n391), .B(KEYINPUT39), .C1(new_n370), .C2(new_n393), .ZN(new_n394));
  XNOR2_X1  g193(.A(G1gat), .B(G29gat), .ZN(new_n395));
  INV_X1    g194(.A(G85gat), .ZN(new_n396));
  XNOR2_X1  g195(.A(new_n395), .B(new_n396), .ZN(new_n397));
  XNOR2_X1  g196(.A(KEYINPUT0), .B(G57gat), .ZN(new_n398));
  XOR2_X1   g197(.A(new_n397), .B(new_n398), .Z(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  OAI211_X1 g199(.A(new_n394), .B(new_n400), .C1(KEYINPUT39), .C2(new_n391), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT40), .ZN(new_n402));
  OR2_X1    g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n379), .A2(new_n390), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n370), .A2(KEYINPUT5), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  NOR3_X1   g206(.A1(new_n277), .A2(new_n388), .A3(new_n380), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n370), .B1(new_n389), .B2(new_n388), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n387), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g209(.A(KEYINPUT5), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n393), .A2(new_n370), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(KEYINPUT82), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT82), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n393), .A2(new_n414), .A3(new_n370), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n411), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n399), .B1(new_n407), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n418));
  AND3_X1   g217(.A1(new_n403), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n368), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n331), .A2(new_n332), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n378), .B1(new_n421), .B2(new_n385), .ZN(new_n422));
  INV_X1    g221(.A(G228gat), .ZN(new_n423));
  INV_X1    g222(.A(G233gat), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT29), .B1(new_n378), .B2(new_n385), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n331), .A2(new_n427), .ZN(new_n428));
  NOR3_X1   g227(.A1(new_n422), .A2(new_n426), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n339), .A2(KEYINPUT83), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n330), .A2(KEYINPUT83), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n431), .A2(KEYINPUT29), .ZN(new_n432));
  AOI21_X1  g231(.A(KEYINPUT3), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n433), .A2(new_n378), .ZN(new_n434));
  OAI211_X1 g233(.A(KEYINPUT84), .B(new_n426), .C1(new_n434), .C2(new_n428), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT84), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT83), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n432), .B1(new_n437), .B2(new_n331), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(new_n385), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n428), .B1(new_n439), .B2(new_n380), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n436), .B1(new_n440), .B2(new_n425), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n429), .B1(new_n435), .B2(new_n441), .ZN(new_n442));
  XNOR2_X1  g241(.A(G78gat), .B(G106gat), .ZN(new_n443));
  INV_X1    g242(.A(G22gat), .ZN(new_n444));
  XNOR2_X1  g243(.A(new_n443), .B(new_n444), .ZN(new_n445));
  XNOR2_X1  g244(.A(KEYINPUT31), .B(G50gat), .ZN(new_n446));
  XOR2_X1   g245(.A(new_n445), .B(new_n446), .Z(new_n447));
  NOR2_X1   g246(.A1(new_n442), .A2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n447), .ZN(new_n449));
  AOI211_X1 g248(.A(new_n429), .B(new_n449), .C1(new_n435), .C2(new_n441), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n342), .A2(KEYINPUT37), .A3(new_n352), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT37), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n361), .A2(new_n453), .A3(new_n347), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n452), .A2(new_n345), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(KEYINPUT38), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT6), .ZN(new_n457));
  AND2_X1   g256(.A1(new_n413), .A2(new_n415), .ZN(new_n458));
  OAI211_X1 g257(.A(new_n400), .B(new_n406), .C1(new_n458), .C2(new_n411), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n417), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  OAI211_X1 g259(.A(KEYINPUT6), .B(new_n399), .C1(new_n407), .C2(new_n416), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n453), .B1(new_n350), .B2(new_n339), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n338), .A2(new_n331), .ZN(new_n465));
  AOI211_X1 g264(.A(KEYINPUT38), .B(new_n362), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(new_n454), .ZN(new_n467));
  AND3_X1   g266(.A1(new_n463), .A2(new_n363), .A3(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n451), .B1(new_n456), .B2(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n306), .B1(new_n420), .B2(new_n469), .ZN(new_n470));
  XOR2_X1   g269(.A(new_n451), .B(KEYINPUT85), .Z(new_n471));
  OAI21_X1  g270(.A(new_n471), .B1(new_n368), .B2(new_n463), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n451), .B1(new_n297), .B2(new_n303), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n357), .A2(new_n462), .A3(new_n367), .A4(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT35), .ZN(new_n475));
  AND3_X1   g274(.A1(new_n297), .A2(new_n303), .A3(KEYINPUT86), .ZN(new_n476));
  AOI21_X1  g275(.A(KEYINPUT86), .B1(new_n297), .B2(new_n303), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT35), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n478), .B1(new_n448), .B2(new_n450), .ZN(new_n479));
  NOR3_X1   g278(.A1(new_n476), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n480), .A2(new_n462), .A3(new_n357), .A4(new_n367), .ZN(new_n481));
  AOI22_X1  g280(.A1(new_n470), .A2(new_n472), .B1(new_n475), .B2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  XNOR2_X1  g282(.A(G120gat), .B(G148gat), .ZN(new_n484));
  XNOR2_X1  g283(.A(G176gat), .B(G204gat), .ZN(new_n485));
  XNOR2_X1  g284(.A(new_n484), .B(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(G230gat), .A2(G233gat), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(G71gat), .ZN(new_n490));
  INV_X1    g289(.A(G78gat), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n490), .A2(new_n491), .A3(KEYINPUT9), .ZN(new_n492));
  NAND2_X1  g291(.A1(G71gat), .A2(G78gat), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(G64gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(G57gat), .ZN(new_n496));
  INV_X1    g295(.A(G57gat), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(G64gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n494), .B1(new_n499), .B2(KEYINPUT94), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n500), .B1(KEYINPUT94), .B2(new_n499), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT95), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n501), .B(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n490), .A2(new_n491), .ZN(new_n504));
  XNOR2_X1  g303(.A(G57gat), .B(G64gat), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT92), .ZN(new_n506));
  OAI21_X1  g305(.A(KEYINPUT9), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n499), .A2(KEYINPUT92), .ZN(new_n508));
  OAI211_X1 g307(.A(new_n493), .B(new_n504), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n509), .B(KEYINPUT93), .ZN(new_n510));
  NAND2_X1  g309(.A1(G99gat), .A2(G106gat), .ZN(new_n511));
  INV_X1    g310(.A(G92gat), .ZN(new_n512));
  AOI22_X1  g311(.A1(KEYINPUT8), .A2(new_n511), .B1(new_n396), .B2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT7), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n514), .B1(new_n396), .B2(new_n512), .ZN(new_n515));
  NAND3_X1  g314(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n513), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  XNOR2_X1  g316(.A(G99gat), .B(G106gat), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n517), .B(new_n518), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n503), .A2(new_n510), .A3(KEYINPUT10), .A4(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n520), .B(KEYINPUT99), .ZN(new_n521));
  INV_X1    g320(.A(new_n518), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(KEYINPUT98), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n503), .A2(new_n510), .A3(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n519), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT10), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n503), .A2(new_n510), .A3(new_n519), .A4(new_n523), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n489), .B1(new_n521), .B2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT101), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n530), .B(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n526), .A2(new_n528), .ZN(new_n533));
  AND3_X1   g332(.A1(new_n533), .A2(KEYINPUT100), .A3(new_n489), .ZN(new_n534));
  AOI21_X1  g333(.A(KEYINPUT100), .B1(new_n533), .B2(new_n489), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n487), .B1(new_n532), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n529), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(new_n488), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n536), .A2(new_n539), .A3(new_n487), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  NAND3_X1  g342(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n544));
  NAND2_X1  g343(.A1(G29gat), .A2(G36gat), .ZN(new_n545));
  OAI21_X1  g344(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  NOR3_X1   g346(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n545), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(G43gat), .B(G50gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(KEYINPUT88), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(KEYINPUT15), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n550), .A2(KEYINPUT88), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n549), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n552), .A2(new_n553), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT15), .ZN(new_n556));
  XNOR2_X1  g355(.A(KEYINPUT89), .B(G50gat), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(G43gat), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n560), .B1(new_n559), .B2(G50gat), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n555), .B1(new_n556), .B2(new_n561), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n554), .B1(new_n562), .B2(new_n549), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n544), .B1(new_n563), .B2(new_n525), .ZN(new_n564));
  NOR3_X1   g363(.A1(new_n563), .A2(KEYINPUT90), .A3(KEYINPUT17), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  OAI21_X1  g365(.A(KEYINPUT90), .B1(new_n563), .B2(KEYINPUT17), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n519), .B1(new_n563), .B2(KEYINPUT17), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n564), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  XOR2_X1   g369(.A(G190gat), .B(G218gat), .Z(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(KEYINPUT97), .ZN(new_n573));
  XNOR2_X1  g372(.A(G134gat), .B(G162gat), .ZN(new_n574));
  AOI21_X1  g373(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n573), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n570), .B(new_n571), .ZN(new_n578));
  OR2_X1    g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n577), .A2(new_n578), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(G15gat), .B(G22gat), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT16), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n582), .B1(new_n583), .B2(G1gat), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n584), .B1(G1gat), .B2(new_n582), .ZN(new_n585));
  INV_X1    g384(.A(G8gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  AND2_X1   g387(.A1(new_n503), .A2(new_n510), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n588), .B1(new_n589), .B2(KEYINPUT21), .ZN(new_n590));
  XOR2_X1   g389(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  XOR2_X1   g391(.A(G127gat), .B(G155gat), .Z(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(KEYINPUT96), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n592), .B(new_n594), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n589), .A2(KEYINPUT21), .ZN(new_n596));
  NAND2_X1  g395(.A1(G231gat), .A2(G233gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(new_n210), .ZN(new_n598));
  INV_X1    g397(.A(G211gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n596), .B(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n595), .B(new_n601), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n563), .A2(new_n587), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n588), .B1(new_n563), .B2(KEYINPUT17), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n603), .B1(new_n568), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(G229gat), .A2(G233gat), .ZN(new_n606));
  AOI21_X1  g405(.A(KEYINPUT18), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n567), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n604), .B1(new_n608), .B2(new_n565), .ZN(new_n609));
  INV_X1    g408(.A(new_n603), .ZN(new_n610));
  NAND4_X1  g409(.A1(new_n609), .A2(KEYINPUT18), .A3(new_n606), .A4(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n563), .B(new_n587), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n606), .B(KEYINPUT13), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n607), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n611), .A2(KEYINPUT91), .A3(new_n615), .ZN(new_n618));
  XOR2_X1   g417(.A(G169gat), .B(G197gat), .Z(new_n619));
  XNOR2_X1  g418(.A(G113gat), .B(G141gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  XOR2_X1   g420(.A(KEYINPUT87), .B(KEYINPUT11), .Z(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XOR2_X1   g422(.A(new_n623), .B(KEYINPUT12), .Z(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n618), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n617), .A2(new_n626), .ZN(new_n627));
  OAI211_X1 g426(.A(new_n618), .B(new_n625), .C1(new_n607), .C2(new_n616), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NOR4_X1   g429(.A1(new_n543), .A2(new_n581), .A3(new_n602), .A4(new_n630), .ZN(new_n631));
  AND2_X1   g430(.A1(new_n483), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(new_n463), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g433(.A1(new_n632), .A2(new_n368), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  OAI21_X1  g435(.A(KEYINPUT42), .B1(new_n636), .B2(new_n586), .ZN(new_n637));
  NAND2_X1  g436(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n583), .A2(new_n586), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n636), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  MUX2_X1   g439(.A(KEYINPUT42), .B(new_n637), .S(new_n640), .Z(G1325gat));
  NAND3_X1  g440(.A1(new_n632), .A2(G15gat), .A3(new_n306), .ZN(new_n642));
  INV_X1    g441(.A(G15gat), .ZN(new_n643));
  INV_X1    g442(.A(new_n632), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n476), .A2(new_n477), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n643), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT102), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n642), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n649), .B1(new_n648), .B2(new_n647), .ZN(G1326gat));
  NAND2_X1  g449(.A1(new_n632), .A2(new_n471), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(new_n444), .ZN(new_n652));
  XNOR2_X1  g451(.A(KEYINPUT103), .B(KEYINPUT43), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(G1327gat));
  INV_X1    g453(.A(new_n581), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n482), .A2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n602), .ZN(new_n657));
  NOR3_X1   g456(.A1(new_n543), .A2(new_n657), .A3(new_n630), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  NOR3_X1   g458(.A1(new_n659), .A2(G29gat), .A3(new_n462), .ZN(new_n660));
  XOR2_X1   g459(.A(new_n660), .B(KEYINPUT45), .Z(new_n661));
  NAND2_X1  g460(.A1(new_n470), .A2(new_n472), .ZN(new_n662));
  AND3_X1   g461(.A1(new_n475), .A2(KEYINPUT104), .A3(new_n481), .ZN(new_n663));
  AOI21_X1  g462(.A(KEYINPUT104), .B1(new_n475), .B2(new_n481), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n662), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT44), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n665), .A2(new_n666), .A3(new_n581), .ZN(new_n667));
  OAI21_X1  g466(.A(KEYINPUT44), .B1(new_n482), .B2(new_n655), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(new_n658), .ZN(new_n670));
  OAI21_X1  g469(.A(G29gat), .B1(new_n670), .B2(new_n462), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n661), .A2(new_n671), .ZN(G1328gat));
  INV_X1    g471(.A(new_n368), .ZN(new_n673));
  NOR3_X1   g472(.A1(new_n659), .A2(G36gat), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(KEYINPUT46), .ZN(new_n675));
  OAI21_X1  g474(.A(G36gat), .B1(new_n670), .B2(new_n673), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(G1329gat));
  INV_X1    g476(.A(KEYINPUT106), .ZN(new_n678));
  NOR3_X1   g477(.A1(new_n659), .A2(G43gat), .A3(new_n646), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n669), .A2(new_n306), .A3(new_n658), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n679), .B1(new_n680), .B2(G43gat), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n678), .B1(new_n681), .B2(KEYINPUT105), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT47), .ZN(new_n683));
  OR2_X1    g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n682), .A2(new_n683), .ZN(new_n685));
  OR2_X1    g484(.A1(new_n681), .A2(new_n678), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n684), .A2(new_n685), .A3(new_n686), .ZN(G1330gat));
  INV_X1    g486(.A(new_n451), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n558), .B1(new_n670), .B2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n471), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n659), .A2(new_n690), .A3(new_n558), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n689), .A2(KEYINPUT48), .A3(new_n692), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n669), .A2(new_n471), .A3(new_n658), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n691), .B1(new_n694), .B2(new_n558), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n693), .B1(new_n695), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR2_X1   g495(.A1(new_n581), .A2(new_n602), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(new_n630), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n475), .A2(new_n481), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT104), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n475), .A2(new_n481), .A3(KEYINPUT104), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  AOI211_X1 g502(.A(new_n542), .B(new_n698), .C1(new_n703), .C2(new_n662), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(new_n463), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g505(.A1(new_n704), .A2(new_n368), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n707), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n708));
  XOR2_X1   g507(.A(KEYINPUT49), .B(G64gat), .Z(new_n709));
  OAI21_X1  g508(.A(new_n708), .B1(new_n707), .B2(new_n709), .ZN(G1333gat));
  NAND3_X1  g509(.A1(new_n704), .A2(G71gat), .A3(new_n306), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(KEYINPUT107), .ZN(new_n712));
  AND2_X1   g511(.A1(new_n704), .A2(new_n645), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n712), .B1(G71gat), .B2(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g514(.A1(new_n704), .A2(new_n471), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g516(.A1(new_n657), .A2(new_n629), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(new_n543), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n719), .B1(new_n667), .B2(new_n668), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  OAI21_X1  g520(.A(G85gat), .B1(new_n721), .B2(new_n462), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n655), .B1(new_n703), .B2(new_n662), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n723), .A2(KEYINPUT51), .A3(new_n718), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n665), .A2(new_n581), .A3(new_n718), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT51), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n728), .A2(new_n396), .A3(new_n463), .A4(new_n543), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n722), .A2(new_n729), .ZN(G1336gat));
  AOI21_X1  g529(.A(new_n512), .B1(new_n720), .B2(new_n368), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT52), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n673), .A2(G92gat), .ZN(new_n734));
  AOI21_X1  g533(.A(KEYINPUT51), .B1(new_n723), .B2(new_n718), .ZN(new_n735));
  AND4_X1   g534(.A1(KEYINPUT51), .A2(new_n665), .A3(new_n581), .A4(new_n718), .ZN(new_n736));
  OAI211_X1 g535(.A(new_n543), .B(new_n734), .C1(new_n735), .C2(new_n736), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n732), .A2(new_n733), .A3(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT108), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n731), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  NAND4_X1  g539(.A1(new_n728), .A2(KEYINPUT108), .A3(new_n543), .A4(new_n734), .ZN(new_n741));
  AOI211_X1 g540(.A(KEYINPUT109), .B(new_n733), .C1(new_n740), .C2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT109), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n737), .A2(new_n739), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n744), .A2(new_n741), .A3(new_n732), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n743), .B1(new_n745), .B2(KEYINPUT52), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n738), .B1(new_n742), .B2(new_n746), .ZN(G1337gat));
  NOR2_X1   g546(.A1(new_n646), .A2(G99gat), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n728), .A2(new_n543), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n720), .A2(new_n306), .ZN(new_n750));
  AND2_X1   g549(.A1(new_n750), .A2(KEYINPUT110), .ZN(new_n751));
  OAI21_X1  g550(.A(G99gat), .B1(new_n750), .B2(KEYINPUT110), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n749), .B1(new_n751), .B2(new_n752), .ZN(G1338gat));
  OAI21_X1  g552(.A(G106gat), .B1(new_n721), .B2(new_n690), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT111), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NOR3_X1   g555(.A1(new_n542), .A2(G106gat), .A3(new_n688), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(KEYINPUT112), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n728), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n756), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n754), .A2(new_n755), .ZN(new_n761));
  OAI21_X1  g560(.A(KEYINPUT53), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(G106gat), .B1(new_n721), .B2(new_n688), .ZN(new_n763));
  AOI21_X1  g562(.A(KEYINPUT53), .B1(new_n728), .B2(new_n757), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n762), .A2(new_n765), .ZN(G1339gat));
  NOR2_X1   g565(.A1(new_n698), .A2(new_n543), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT55), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n539), .A2(new_n531), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n530), .A2(KEYINPUT101), .ZN(new_n771));
  AOI21_X1  g570(.A(KEYINPUT54), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n521), .A2(new_n529), .A3(new_n489), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n539), .A2(KEYINPUT54), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(new_n486), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n769), .B1(new_n772), .B2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT54), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n530), .A2(new_n777), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n487), .B1(new_n778), .B2(new_n773), .ZN(new_n779));
  OAI211_X1 g578(.A(new_n779), .B(KEYINPUT55), .C1(new_n532), .C2(KEYINPUT54), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n629), .A2(new_n776), .A3(new_n780), .A4(new_n540), .ZN(new_n781));
  OR2_X1    g580(.A1(new_n605), .A2(new_n606), .ZN(new_n782));
  OR2_X1    g581(.A1(new_n612), .A2(new_n614), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(new_n623), .ZN(new_n785));
  AOI22_X1  g584(.A1(new_n617), .A2(new_n624), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n786), .B1(new_n537), .B2(new_n541), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n781), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(new_n655), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT113), .ZN(new_n790));
  AND2_X1   g589(.A1(new_n776), .A2(new_n540), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n791), .A2(new_n581), .A3(new_n780), .A4(new_n786), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n789), .A2(new_n790), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(new_n602), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n790), .B1(new_n789), .B2(new_n792), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n768), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(new_n690), .ZN(new_n797));
  OR2_X1    g596(.A1(new_n797), .A2(KEYINPUT114), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(KEYINPUT114), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n646), .A2(new_n368), .A3(new_n462), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  OAI21_X1  g601(.A(G113gat), .B1(new_n802), .B2(new_n630), .ZN(new_n803));
  AND2_X1   g602(.A1(new_n796), .A2(new_n473), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n368), .A2(new_n462), .ZN(new_n805));
  AND2_X1   g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n630), .A2(G113gat), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n807), .B(KEYINPUT115), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n803), .A2(new_n809), .ZN(G1340gat));
  INV_X1    g609(.A(G120gat), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n806), .A2(new_n811), .A3(new_n543), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT116), .ZN(new_n813));
  INV_X1    g612(.A(new_n802), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(new_n543), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n813), .B1(new_n815), .B2(G120gat), .ZN(new_n816));
  AOI211_X1 g615(.A(KEYINPUT116), .B(new_n811), .C1(new_n814), .C2(new_n543), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n812), .B1(new_n816), .B2(new_n817), .ZN(G1341gat));
  AOI21_X1  g617(.A(G127gat), .B1(new_n806), .B2(new_n657), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n657), .A2(G127gat), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n819), .B1(new_n814), .B2(new_n820), .ZN(G1342gat));
  OAI21_X1  g620(.A(G134gat), .B1(new_n802), .B2(new_n655), .ZN(new_n822));
  OR2_X1    g621(.A1(new_n822), .A2(KEYINPUT117), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(KEYINPUT117), .ZN(new_n824));
  INV_X1    g623(.A(G134gat), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n806), .A2(new_n825), .A3(new_n581), .ZN(new_n826));
  XOR2_X1   g625(.A(new_n826), .B(KEYINPUT56), .Z(new_n827));
  NAND3_X1  g626(.A1(new_n823), .A2(new_n824), .A3(new_n827), .ZN(G1343gat));
  NAND2_X1  g627(.A1(new_n805), .A2(new_n305), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n796), .A2(new_n451), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n831), .A2(KEYINPUT57), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT118), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n781), .A2(new_n833), .A3(new_n787), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(new_n655), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n833), .B1(new_n781), .B2(new_n787), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n792), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n767), .B1(new_n837), .B2(new_n602), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT57), .ZN(new_n839));
  NOR3_X1   g638(.A1(new_n838), .A2(new_n839), .A3(new_n690), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n830), .B1(new_n832), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(G141gat), .B1(new_n841), .B2(new_n630), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n831), .A2(new_n830), .ZN(new_n843));
  INV_X1    g642(.A(G141gat), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n843), .A2(new_n844), .A3(new_n629), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g645(.A(new_n846), .B(KEYINPUT58), .ZN(G1344gat));
  INV_X1    g646(.A(G148gat), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n843), .A2(new_n848), .A3(new_n543), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n848), .A2(KEYINPUT59), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n850), .B1(new_n841), .B2(new_n542), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT119), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n851), .B(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT59), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n837), .A2(new_n602), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(new_n768), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT120), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n690), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  AOI211_X1 g657(.A(new_n857), .B(new_n767), .C1(new_n837), .C2(new_n602), .ZN(new_n859));
  INV_X1    g658(.A(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(KEYINPUT57), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n796), .A2(KEYINPUT57), .A3(new_n451), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n543), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  OR2_X1    g663(.A1(new_n864), .A2(new_n829), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n854), .B1(new_n865), .B2(G148gat), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n849), .B1(new_n853), .B2(new_n866), .ZN(G1345gat));
  NOR3_X1   g666(.A1(new_n841), .A2(new_n373), .A3(new_n602), .ZN(new_n868));
  AOI21_X1  g667(.A(G155gat), .B1(new_n843), .B2(new_n657), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n868), .A2(new_n869), .ZN(G1346gat));
  OAI21_X1  g669(.A(G162gat), .B1(new_n841), .B2(new_n655), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n843), .A2(new_n374), .A3(new_n581), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g672(.A(new_n873), .B(KEYINPUT121), .ZN(G1347gat));
  INV_X1    g673(.A(G169gat), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n673), .A2(new_n463), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(new_n645), .ZN(new_n877));
  XNOR2_X1  g676(.A(new_n877), .B(KEYINPUT122), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n878), .B1(new_n798), .B2(new_n799), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n875), .B1(new_n879), .B2(new_n629), .ZN(new_n880));
  AND2_X1   g679(.A1(new_n804), .A2(new_n876), .ZN(new_n881));
  AND3_X1   g680(.A1(new_n881), .A2(new_n875), .A3(new_n629), .ZN(new_n882));
  OR2_X1    g681(.A1(new_n880), .A2(new_n882), .ZN(G1348gat));
  NAND3_X1  g682(.A1(new_n879), .A2(G176gat), .A3(new_n543), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n884), .A2(KEYINPUT123), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n884), .A2(KEYINPUT123), .ZN(new_n886));
  AOI21_X1  g685(.A(G176gat), .B1(new_n881), .B2(new_n543), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(G1349gat));
  AOI21_X1  g687(.A(new_n210), .B1(new_n879), .B2(new_n657), .ZN(new_n889));
  NAND4_X1  g688(.A1(new_n881), .A2(new_n214), .A3(new_n215), .A4(new_n657), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(KEYINPUT124), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT60), .ZN(new_n893));
  XNOR2_X1  g692(.A(new_n892), .B(new_n893), .ZN(G1350gat));
  NAND3_X1  g693(.A1(new_n881), .A2(new_n211), .A3(new_n581), .ZN(new_n895));
  XOR2_X1   g694(.A(new_n895), .B(KEYINPUT125), .Z(new_n896));
  AOI211_X1 g695(.A(KEYINPUT61), .B(new_n211), .C1(new_n879), .C2(new_n581), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT61), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n879), .A2(new_n581), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n898), .B1(new_n899), .B2(G190gat), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n896), .B1(new_n897), .B2(new_n900), .ZN(G1351gat));
  INV_X1    g700(.A(G197gat), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n673), .A2(new_n306), .A3(new_n463), .ZN(new_n903));
  XNOR2_X1  g702(.A(new_n903), .B(KEYINPUT126), .ZN(new_n904));
  INV_X1    g703(.A(new_n904), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n471), .B1(new_n838), .B2(KEYINPUT120), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n839), .B1(new_n906), .B2(new_n859), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n905), .B1(new_n907), .B2(new_n862), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n902), .B1(new_n908), .B2(new_n629), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n831), .A2(new_n903), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n910), .A2(G197gat), .A3(new_n630), .ZN(new_n911));
  OR2_X1    g710(.A1(new_n909), .A2(new_n911), .ZN(G1352gat));
  NOR3_X1   g711(.A1(new_n910), .A2(G204gat), .A3(new_n542), .ZN(new_n913));
  XNOR2_X1  g712(.A(new_n913), .B(KEYINPUT62), .ZN(new_n914));
  OAI21_X1  g713(.A(G204gat), .B1(new_n864), .B2(new_n905), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(G1353gat));
  OR3_X1    g715(.A1(new_n910), .A2(new_n321), .A3(new_n602), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT63), .ZN(new_n918));
  AOI211_X1 g717(.A(new_n918), .B(new_n599), .C1(new_n908), .C2(new_n657), .ZN(new_n919));
  OAI211_X1 g718(.A(new_n657), .B(new_n904), .C1(new_n861), .C2(new_n863), .ZN(new_n920));
  AOI21_X1  g719(.A(KEYINPUT63), .B1(new_n920), .B2(G211gat), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n917), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(KEYINPUT127), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT127), .ZN(new_n924));
  OAI211_X1 g723(.A(new_n924), .B(new_n917), .C1(new_n919), .C2(new_n921), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n923), .A2(new_n925), .ZN(G1354gat));
  INV_X1    g725(.A(new_n910), .ZN(new_n927));
  AOI21_X1  g726(.A(G218gat), .B1(new_n927), .B2(new_n581), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n581), .A2(G218gat), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n928), .B1(new_n908), .B2(new_n929), .ZN(G1355gat));
endmodule


