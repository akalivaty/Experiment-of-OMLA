//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 0 1 0 1 0 1 1 0 0 0 1 0 1 1 0 0 0 0 1 0 0 1 1 1 0 0 0 1 1 0 0 0 0 0 1 0 1 0 1 1 0 1 0 0 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:53 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n552, new_n554, new_n555, new_n556, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n619, new_n621, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1185;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT65), .B(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT66), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT68), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G125), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n462), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT69), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n465), .A2(G2105), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  AND2_X1   g046(.A1(new_n471), .A2(G2104), .ZN(new_n472));
  AOI22_X1  g047(.A1(new_n470), .A2(G137), .B1(G101), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n468), .A2(KEYINPUT69), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n474), .A2(new_n475), .ZN(G160));
  NAND2_X1  g051(.A1(new_n470), .A2(G136), .ZN(new_n477));
  MUX2_X1   g052(.A(G100), .B(G112), .S(G2105), .Z(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G2104), .ZN(new_n479));
  INV_X1    g054(.A(G124), .ZN(new_n480));
  XNOR2_X1  g055(.A(KEYINPUT3), .B(G2104), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n477), .B(new_n479), .C1(new_n480), .C2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  NAND2_X1  g059(.A1(G114), .A2(G2105), .ZN(new_n485));
  INV_X1    g060(.A(G102), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n485), .B1(new_n486), .B2(G2105), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G2104), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(KEYINPUT71), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT71), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n487), .A2(new_n490), .A3(G2104), .ZN(new_n491));
  OAI211_X1 g066(.A(G126), .B(G2105), .C1(new_n463), .C2(new_n464), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT70), .ZN(new_n494));
  AOI22_X1  g069(.A1(new_n489), .A2(new_n491), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  OAI211_X1 g070(.A(G138), .B(new_n471), .C1(new_n463), .C2(new_n464), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT72), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n481), .A2(KEYINPUT72), .A3(G138), .A4(new_n471), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n498), .A2(new_n499), .A3(KEYINPUT4), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n496), .A2(new_n497), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n492), .A2(KEYINPUT70), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n495), .A2(new_n500), .A3(new_n502), .A4(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(G164));
  AND2_X1   g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  NOR2_X1   g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  OAI211_X1 g082(.A(G50), .B(G543), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  NOR2_X1   g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  OAI22_X1  g086(.A1(new_n510), .A2(new_n511), .B1(new_n506), .B2(new_n507), .ZN(new_n512));
  INV_X1    g087(.A(G88), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n508), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  OAI21_X1  g090(.A(G62), .B1(new_n510), .B2(new_n511), .ZN(new_n516));
  NAND2_X1  g091(.A1(G75), .A2(G543), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n514), .A2(new_n518), .ZN(G166));
  NAND3_X1  g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n520), .B(KEYINPUT7), .ZN(new_n521));
  OR2_X1    g096(.A1(KEYINPUT6), .A2(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(KEYINPUT6), .A2(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G543), .ZN(new_n525));
  INV_X1    g100(.A(G51), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n521), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n510), .A2(new_n511), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n524), .A2(G89), .ZN(new_n529));
  NAND2_X1  g104(.A1(G63), .A2(G651), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n527), .A2(new_n531), .ZN(G168));
  OR2_X1    g107(.A1(KEYINPUT5), .A2(G543), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(new_n509), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n534), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n535), .A2(new_n515), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT73), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n536), .B(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(G52), .ZN(new_n539));
  INV_X1    g114(.A(G90), .ZN(new_n540));
  OAI22_X1  g115(.A1(new_n525), .A2(new_n539), .B1(new_n512), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n538), .A2(new_n541), .ZN(G171));
  AOI22_X1  g117(.A1(new_n534), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n543), .A2(new_n515), .ZN(new_n544));
  INV_X1    g119(.A(G43), .ZN(new_n545));
  INV_X1    g120(.A(G81), .ZN(new_n546));
  OAI22_X1  g121(.A1(new_n525), .A2(new_n545), .B1(new_n512), .B2(new_n546), .ZN(new_n547));
  OR2_X1    g122(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT74), .ZN(G153));
  AND3_X1   g126(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G36), .ZN(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  XOR2_X1   g131(.A(new_n556), .B(KEYINPUT75), .Z(G188));
  XOR2_X1   g132(.A(KEYINPUT76), .B(KEYINPUT9), .Z(new_n558));
  INV_X1    g133(.A(G53), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n525), .B2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(G543), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n561), .B1(new_n522), .B2(new_n523), .ZN(new_n562));
  NAND4_X1  g137(.A1(new_n562), .A2(KEYINPUT76), .A3(KEYINPUT9), .A4(G53), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(G78), .A2(G543), .ZN(new_n566));
  INV_X1    g141(.A(G65), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n566), .B1(new_n528), .B2(new_n567), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n533), .A2(new_n509), .B1(new_n522), .B2(new_n523), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n568), .A2(G651), .B1(new_n569), .B2(G91), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n565), .A2(new_n570), .ZN(G299));
  INV_X1    g146(.A(G171), .ZN(G301));
  INV_X1    g147(.A(G168), .ZN(G286));
  OAI21_X1  g148(.A(KEYINPUT77), .B1(new_n514), .B2(new_n518), .ZN(new_n574));
  INV_X1    g149(.A(G62), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n575), .B1(new_n533), .B2(new_n509), .ZN(new_n576));
  INV_X1    g151(.A(new_n517), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT77), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n534), .A2(new_n524), .A3(G88), .ZN(new_n580));
  NAND4_X1  g155(.A1(new_n578), .A2(new_n579), .A3(new_n580), .A4(new_n508), .ZN(new_n581));
  AND2_X1   g156(.A1(new_n574), .A2(new_n581), .ZN(G303));
  NAND2_X1  g157(.A1(new_n569), .A2(G87), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n562), .A2(G49), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n534), .B2(G74), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(G288));
  NAND2_X1  g161(.A1(new_n569), .A2(G86), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n562), .A2(G48), .ZN(new_n588));
  AND2_X1   g163(.A1(G73), .A2(G543), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n589), .B1(new_n534), .B2(G61), .ZN(new_n590));
  OAI211_X1 g165(.A(new_n587), .B(new_n588), .C1(new_n590), .C2(new_n515), .ZN(G305));
  AOI22_X1  g166(.A1(new_n534), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n592), .A2(new_n515), .ZN(new_n593));
  INV_X1    g168(.A(G47), .ZN(new_n594));
  INV_X1    g169(.A(G85), .ZN(new_n595));
  OAI22_X1  g170(.A1(new_n525), .A2(new_n594), .B1(new_n512), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(G290));
  NAND3_X1  g173(.A1(G301), .A2(KEYINPUT78), .A3(G868), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT78), .ZN(new_n600));
  INV_X1    g175(.A(G868), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(G171), .B2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(G92), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n512), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(KEYINPUT10), .ZN(new_n605));
  NAND2_X1  g180(.A1(G79), .A2(G543), .ZN(new_n606));
  INV_X1    g181(.A(G66), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n528), .B2(new_n607), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n608), .A2(G651), .B1(G54), .B2(new_n562), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n605), .A2(new_n609), .ZN(new_n610));
  AND2_X1   g185(.A1(new_n610), .A2(KEYINPUT79), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n610), .A2(KEYINPUT79), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(new_n613), .ZN(new_n614));
  OAI211_X1 g189(.A(new_n599), .B(new_n602), .C1(new_n614), .C2(G868), .ZN(G284));
  XNOR2_X1  g190(.A(G284), .B(KEYINPUT80), .ZN(G321));
  MUX2_X1   g191(.A(G286), .B(G299), .S(new_n601), .Z(G297));
  MUX2_X1   g192(.A(G286), .B(G299), .S(new_n601), .Z(G280));
  INV_X1    g193(.A(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n614), .B1(new_n619), .B2(G860), .ZN(G148));
  NOR2_X1   g195(.A1(new_n548), .A2(G868), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n613), .A2(G559), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n621), .B1(new_n622), .B2(G868), .ZN(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g199(.A1(new_n470), .A2(G2104), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT12), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT13), .ZN(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT81), .B(G2100), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n627), .A2(new_n628), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n470), .A2(G135), .ZN(new_n631));
  MUX2_X1   g206(.A(G99), .B(G111), .S(G2105), .Z(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(G2104), .ZN(new_n633));
  INV_X1    g208(.A(G123), .ZN(new_n634));
  OAI211_X1 g209(.A(new_n631), .B(new_n633), .C1(new_n634), .C2(new_n482), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(G2096), .Z(new_n636));
  NAND3_X1  g211(.A1(new_n629), .A2(new_n630), .A3(new_n636), .ZN(G156));
  XNOR2_X1  g212(.A(G2451), .B(G2454), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT16), .ZN(new_n639));
  XOR2_X1   g214(.A(G2443), .B(G2446), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(G1341), .B(G1348), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  INV_X1    g218(.A(KEYINPUT14), .ZN(new_n644));
  XOR2_X1   g219(.A(KEYINPUT15), .B(G2435), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2438), .ZN(new_n646));
  XOR2_X1   g221(.A(G2427), .B(G2430), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT82), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n644), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n649), .B1(new_n646), .B2(new_n648), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n643), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n643), .A2(new_n650), .ZN(new_n652));
  AND3_X1   g227(.A1(new_n651), .A2(G14), .A3(new_n652), .ZN(G401));
  XNOR2_X1  g228(.A(G2067), .B(G2678), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT83), .ZN(new_n655));
  XOR2_X1   g230(.A(G2072), .B(G2078), .Z(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G2084), .B(G2090), .Z(new_n658));
  NAND3_X1  g233(.A1(new_n655), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(KEYINPUT18), .Z(new_n660));
  OR2_X1    g235(.A1(new_n655), .A2(new_n658), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n657), .B1(new_n661), .B2(KEYINPUT17), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n657), .A2(KEYINPUT17), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n655), .B1(new_n664), .B2(new_n658), .ZN(new_n665));
  INV_X1    g240(.A(new_n658), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n665), .B1(new_n666), .B2(new_n663), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n660), .B1(new_n662), .B2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(G2096), .ZN(new_n669));
  XNOR2_X1  g244(.A(KEYINPUT84), .B(G2100), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(G227));
  XOR2_X1   g246(.A(G1971), .B(G1976), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT19), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1956), .B(G2474), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1961), .B(G1966), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  AND2_X1   g251(.A1(new_n674), .A2(new_n675), .ZN(new_n677));
  NOR3_X1   g252(.A1(new_n673), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n673), .A2(new_n676), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT85), .B(KEYINPUT20), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  AOI211_X1 g256(.A(new_n678), .B(new_n681), .C1(new_n673), .C2(new_n677), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1981), .B(G1986), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT86), .ZN(new_n686));
  XOR2_X1   g261(.A(G1991), .B(G1996), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n684), .B(new_n688), .ZN(G229));
  INV_X1    g264(.A(G16), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(G5), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n691), .B1(G171), .B2(new_n690), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(G1961), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n690), .A2(G20), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n694), .B(KEYINPUT23), .Z(new_n695));
  AOI21_X1  g270(.A(new_n695), .B1(G299), .B2(G16), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(G1956), .ZN(new_n697));
  NOR2_X1   g272(.A1(G29), .A2(G35), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n698), .B1(G162), .B2(G29), .ZN(new_n699));
  XOR2_X1   g274(.A(new_n699), .B(KEYINPUT29), .Z(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(new_n701));
  OAI211_X1 g276(.A(new_n693), .B(new_n697), .C1(new_n701), .C2(G2090), .ZN(new_n702));
  INV_X1    g277(.A(G29), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(G33), .ZN(new_n704));
  NAND2_X1  g279(.A1(G115), .A2(G2104), .ZN(new_n705));
  INV_X1    g280(.A(G127), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n705), .B1(new_n465), .B2(new_n706), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n471), .B1(new_n707), .B2(KEYINPUT92), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(KEYINPUT92), .B2(new_n707), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n472), .A2(G103), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT25), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n472), .A2(KEYINPUT25), .A3(G103), .ZN(new_n713));
  AOI22_X1  g288(.A1(new_n712), .A2(new_n713), .B1(new_n470), .B2(G139), .ZN(new_n714));
  AND2_X1   g289(.A1(new_n709), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n704), .B1(new_n715), .B2(new_n703), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT93), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(G2072), .Z(new_n718));
  NOR2_X1   g293(.A1(G29), .A2(G32), .ZN(new_n719));
  INV_X1    g294(.A(new_n482), .ZN(new_n720));
  AOI22_X1  g295(.A1(new_n720), .A2(G129), .B1(new_n470), .B2(G141), .ZN(new_n721));
  NAND3_X1  g296(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT26), .ZN(new_n723));
  OR2_X1    g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n722), .A2(new_n723), .ZN(new_n725));
  AOI22_X1  g300(.A1(new_n724), .A2(new_n725), .B1(G105), .B2(new_n472), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n721), .A2(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT97), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n721), .A2(KEYINPUT97), .A3(new_n726), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n719), .B1(new_n732), .B2(G29), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT98), .Z(new_n734));
  XNOR2_X1  g309(.A(KEYINPUT27), .B(G1996), .ZN(new_n735));
  AOI211_X1 g310(.A(new_n702), .B(new_n718), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(G2090), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n700), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g313(.A1(G168), .A2(new_n690), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(new_n690), .B2(G21), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT99), .B(G1966), .Z(new_n741));
  OR2_X1    g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n740), .A2(new_n741), .ZN(new_n743));
  XOR2_X1   g318(.A(KEYINPUT31), .B(G11), .Z(new_n744));
  NOR2_X1   g319(.A1(new_n635), .A2(new_n703), .ZN(new_n745));
  XOR2_X1   g320(.A(KEYINPUT100), .B(G28), .Z(new_n746));
  OR2_X1    g321(.A1(new_n746), .A2(KEYINPUT30), .ZN(new_n747));
  AOI21_X1  g322(.A(G29), .B1(new_n746), .B2(KEYINPUT30), .ZN(new_n748));
  AOI211_X1 g323(.A(new_n744), .B(new_n745), .C1(new_n747), .C2(new_n748), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n742), .A2(new_n743), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(G164), .A2(G29), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G27), .B2(G29), .ZN(new_n752));
  INV_X1    g327(.A(G2078), .ZN(new_n753));
  AND2_X1   g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n752), .A2(new_n753), .ZN(new_n755));
  NOR4_X1   g330(.A1(new_n738), .A2(new_n750), .A3(new_n754), .A4(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT101), .ZN(new_n757));
  XNOR2_X1  g332(.A(KEYINPUT94), .B(KEYINPUT24), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G34), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n759), .A2(new_n703), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G160), .B2(new_n703), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT95), .Z(new_n762));
  INV_X1    g337(.A(G2084), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  OAI221_X1 g339(.A(new_n764), .B1(G1961), .B2(new_n692), .C1(new_n734), .C2(new_n735), .ZN(new_n765));
  OAI211_X1 g340(.A(new_n736), .B(new_n756), .C1(new_n757), .C2(new_n765), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(new_n757), .B2(new_n765), .ZN(new_n767));
  MUX2_X1   g342(.A(G6), .B(G305), .S(G16), .Z(new_n768));
  XOR2_X1   g343(.A(KEYINPUT32), .B(G1981), .Z(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n690), .A2(G23), .ZN(new_n771));
  INV_X1    g346(.A(G288), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n771), .B1(new_n772), .B2(new_n690), .ZN(new_n773));
  XOR2_X1   g348(.A(KEYINPUT33), .B(G1976), .Z(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT88), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n773), .B(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(G16), .A2(G22), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(G166), .B2(G16), .ZN(new_n778));
  INV_X1    g353(.A(G1971), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n770), .A2(new_n776), .A3(new_n780), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n781), .A2(KEYINPUT34), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n781), .A2(KEYINPUT34), .ZN(new_n783));
  NOR2_X1   g358(.A1(G25), .A2(G29), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n720), .A2(G119), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n470), .A2(G131), .ZN(new_n786));
  MUX2_X1   g361(.A(G95), .B(G107), .S(G2105), .Z(new_n787));
  NAND2_X1  g362(.A1(new_n787), .A2(G2104), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n785), .A2(new_n786), .A3(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(new_n789), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n784), .B1(new_n790), .B2(G29), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT87), .ZN(new_n792));
  XOR2_X1   g367(.A(KEYINPUT35), .B(G1991), .Z(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(G16), .A2(G24), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(new_n597), .B2(G16), .ZN(new_n796));
  INV_X1    g371(.A(G1986), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n782), .A2(new_n783), .A3(new_n794), .A4(new_n798), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT36), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n762), .A2(new_n763), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT96), .ZN(new_n802));
  NOR2_X1   g377(.A1(G4), .A2(G16), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(new_n614), .B2(G16), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n804), .A2(G1348), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n804), .A2(G1348), .ZN(new_n806));
  NOR2_X1   g381(.A1(G16), .A2(G19), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(new_n549), .B2(G16), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(G1341), .Z(new_n809));
  NAND2_X1  g384(.A1(new_n703), .A2(G26), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT89), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT28), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n720), .A2(G128), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n470), .A2(G140), .ZN(new_n814));
  MUX2_X1   g389(.A(G104), .B(G116), .S(G2105), .Z(new_n815));
  NAND2_X1  g390(.A1(new_n815), .A2(G2104), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n813), .A2(new_n814), .A3(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n812), .B1(new_n818), .B2(new_n703), .ZN(new_n819));
  XOR2_X1   g394(.A(KEYINPUT90), .B(G2067), .Z(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  NAND4_X1  g396(.A1(new_n805), .A2(new_n806), .A3(new_n809), .A4(new_n821), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT91), .ZN(new_n823));
  NAND4_X1  g398(.A1(new_n767), .A2(new_n800), .A3(new_n802), .A4(new_n823), .ZN(G150));
  INV_X1    g399(.A(G150), .ZN(G311));
  NOR2_X1   g400(.A1(new_n613), .A2(new_n619), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT38), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT104), .ZN(new_n828));
  AOI22_X1  g403(.A1(new_n534), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n829), .A2(new_n515), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT102), .ZN(new_n831));
  INV_X1    g406(.A(G55), .ZN(new_n832));
  INV_X1    g407(.A(G93), .ZN(new_n833));
  OAI22_X1  g408(.A1(new_n525), .A2(new_n832), .B1(new_n512), .B2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n831), .A2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT103), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n549), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n548), .A2(KEYINPUT103), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n836), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  NAND4_X1  g415(.A1(new_n831), .A2(new_n549), .A3(new_n837), .A4(new_n835), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n828), .B(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT39), .ZN(new_n845));
  AOI21_X1  g420(.A(G860), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n846), .B1(new_n845), .B2(new_n844), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n836), .A2(G860), .ZN(new_n848));
  XOR2_X1   g423(.A(KEYINPUT105), .B(KEYINPUT37), .Z(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n847), .A2(new_n850), .ZN(G145));
  INV_X1    g426(.A(KEYINPUT106), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n715), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(G164), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n731), .B(new_n818), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n854), .B(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n626), .B(new_n790), .ZN(new_n857));
  MUX2_X1   g432(.A(G106), .B(G118), .S(G2105), .Z(new_n858));
  AOI22_X1  g433(.A1(new_n720), .A2(G130), .B1(G2104), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n470), .A2(G142), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n857), .B(new_n861), .ZN(new_n862));
  OR2_X1    g437(.A1(new_n856), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n856), .A2(new_n862), .ZN(new_n864));
  XNOR2_X1  g439(.A(G160), .B(G162), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(new_n635), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n863), .A2(new_n864), .A3(new_n866), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n862), .A2(KEYINPUT107), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n866), .B1(new_n856), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n869), .B1(new_n856), .B2(new_n868), .ZN(new_n870));
  INV_X1    g445(.A(G37), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n867), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g448(.A1(new_n836), .A2(G868), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n843), .B(new_n622), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n610), .A2(new_n570), .A3(new_n565), .ZN(new_n876));
  OR2_X1    g451(.A1(new_n876), .A2(KEYINPUT108), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(KEYINPUT108), .ZN(new_n878));
  NAND3_X1  g453(.A1(G299), .A2(new_n605), .A3(new_n609), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n875), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n880), .B(KEYINPUT41), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n881), .B1(new_n882), .B2(new_n875), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT42), .ZN(new_n884));
  XOR2_X1   g459(.A(G305), .B(G166), .Z(new_n885));
  XNOR2_X1  g460(.A(new_n597), .B(new_n772), .ZN(new_n886));
  XOR2_X1   g461(.A(new_n885), .B(new_n886), .Z(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n884), .B(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n874), .B1(new_n889), .B2(G868), .ZN(G295));
  AOI21_X1  g465(.A(new_n874), .B1(new_n889), .B2(G868), .ZN(G331));
  INV_X1    g466(.A(KEYINPUT44), .ZN(new_n892));
  XNOR2_X1  g467(.A(G168), .B(KEYINPUT109), .ZN(new_n893));
  XNOR2_X1  g468(.A(G171), .B(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n843), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(KEYINPUT110), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT110), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n843), .A2(new_n894), .A3(new_n897), .ZN(new_n898));
  XOR2_X1   g473(.A(G171), .B(new_n893), .Z(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(new_n842), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n896), .A2(new_n898), .A3(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT41), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n880), .B(new_n902), .ZN(new_n903));
  AND2_X1   g478(.A1(new_n900), .A2(new_n895), .ZN(new_n904));
  AOI22_X1  g479(.A1(new_n901), .A2(new_n903), .B1(new_n904), .B2(new_n880), .ZN(new_n905));
  AOI21_X1  g480(.A(G37), .B1(new_n905), .B2(new_n888), .ZN(new_n906));
  INV_X1    g481(.A(new_n880), .ZN(new_n907));
  OAI22_X1  g482(.A1(new_n901), .A2(new_n907), .B1(new_n904), .B2(new_n882), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(new_n887), .ZN(new_n909));
  AND3_X1   g484(.A1(new_n906), .A2(KEYINPUT112), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(KEYINPUT112), .B1(new_n906), .B2(new_n909), .ZN(new_n911));
  OAI21_X1  g486(.A(KEYINPUT43), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT43), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n905), .A2(new_n888), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n901), .A2(new_n903), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n904), .A2(new_n880), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(new_n887), .ZN(new_n918));
  AOI21_X1  g493(.A(KEYINPUT111), .B1(new_n918), .B2(new_n871), .ZN(new_n919));
  OAI211_X1 g494(.A(KEYINPUT111), .B(new_n871), .C1(new_n905), .C2(new_n888), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  OAI211_X1 g496(.A(new_n913), .B(new_n914), .C1(new_n919), .C2(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n892), .B1(new_n912), .B2(new_n922), .ZN(new_n923));
  OAI211_X1 g498(.A(KEYINPUT43), .B(new_n914), .C1(new_n919), .C2(new_n921), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n906), .A2(new_n909), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(new_n913), .ZN(new_n926));
  AOI21_X1  g501(.A(KEYINPUT44), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n923), .A2(new_n927), .ZN(G397));
  INV_X1    g503(.A(KEYINPUT127), .ZN(new_n929));
  XOR2_X1   g504(.A(KEYINPUT113), .B(G1384), .Z(new_n930));
  NAND2_X1  g505(.A1(new_n504), .A2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT45), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n475), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n934), .A2(new_n469), .A3(G40), .A4(new_n473), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n731), .A2(G1996), .ZN(new_n937));
  XOR2_X1   g512(.A(new_n817), .B(G2067), .Z(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(G1996), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n939), .B1(new_n940), .B2(new_n732), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n789), .B(new_n793), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n597), .B(G1986), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n936), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(G8), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n574), .A2(new_n581), .A3(G8), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT55), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT115), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n574), .A2(new_n581), .A3(KEYINPUT55), .A4(G8), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n951), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  AND2_X1   g529(.A1(new_n953), .A2(new_n952), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(G1384), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n489), .A2(new_n491), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n481), .A2(new_n494), .A3(G126), .A4(G2105), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n958), .A2(new_n502), .A3(new_n503), .A4(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(new_n500), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n957), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT114), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT50), .ZN(new_n965));
  OAI211_X1 g540(.A(KEYINPUT114), .B(new_n957), .C1(new_n960), .C2(new_n961), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n935), .B1(new_n962), .B2(KEYINPUT50), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n967), .A2(new_n968), .A3(new_n737), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n962), .A2(new_n932), .ZN(new_n970));
  INV_X1    g545(.A(G40), .ZN(new_n971));
  NOR3_X1   g546(.A1(new_n474), .A2(new_n475), .A3(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n504), .A2(KEYINPUT45), .A3(new_n930), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n970), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(new_n779), .ZN(new_n975));
  AOI211_X1 g550(.A(new_n948), .B(new_n956), .C1(new_n969), .C2(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n964), .A2(new_n966), .A3(new_n972), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n772), .A2(G1976), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n977), .A2(G8), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(KEYINPUT52), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT116), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n981), .B1(new_n590), .B2(new_n515), .ZN(new_n982));
  NAND3_X1  g557(.A1(G305), .A2(G1981), .A3(new_n982), .ZN(new_n983));
  AND2_X1   g558(.A1(new_n534), .A2(G61), .ZN(new_n984));
  OAI21_X1  g559(.A(G651), .B1(new_n984), .B2(new_n589), .ZN(new_n985));
  AOI22_X1  g560(.A1(new_n569), .A2(G86), .B1(new_n562), .B2(G48), .ZN(new_n986));
  INV_X1    g561(.A(G1981), .ZN(new_n987));
  OAI211_X1 g562(.A(new_n985), .B(new_n986), .C1(new_n981), .C2(new_n987), .ZN(new_n988));
  AND2_X1   g563(.A1(new_n983), .A2(new_n988), .ZN(new_n989));
  OR2_X1    g564(.A1(new_n989), .A2(KEYINPUT49), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n983), .A2(KEYINPUT49), .A3(new_n988), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT117), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n983), .A2(new_n988), .A3(KEYINPUT117), .A4(KEYINPUT49), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n990), .A2(new_n995), .A3(new_n977), .A4(G8), .ZN(new_n996));
  INV_X1    g571(.A(G1976), .ZN(new_n997));
  AOI21_X1  g572(.A(KEYINPUT52), .B1(G288), .B2(new_n997), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n977), .A2(G8), .A3(new_n978), .A4(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n980), .A2(new_n996), .A3(new_n999), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n976), .A2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(KEYINPUT45), .B1(new_n964), .B2(new_n966), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n972), .B1(new_n962), .B2(new_n932), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1004), .A2(KEYINPUT53), .A3(new_n753), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n967), .A2(new_n968), .ZN(new_n1006));
  INV_X1    g581(.A(G1961), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT53), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n970), .A2(new_n753), .A3(new_n972), .A4(new_n973), .ZN(new_n1009));
  AOI22_X1  g584(.A1(new_n1006), .A2(new_n1007), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(G301), .B1(new_n1005), .B2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n965), .B1(new_n964), .B2(new_n966), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT118), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n504), .A2(new_n965), .A3(new_n957), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n972), .A2(new_n1014), .ZN(new_n1015));
  NOR3_X1   g590(.A1(new_n1012), .A2(new_n1013), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(new_n966), .ZN(new_n1017));
  AOI21_X1  g592(.A(KEYINPUT114), .B1(new_n504), .B2(new_n957), .ZN(new_n1018));
  OAI21_X1  g593(.A(KEYINPUT50), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  AND2_X1   g594(.A1(new_n972), .A2(new_n1014), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT118), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n737), .B1(new_n1016), .B2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n948), .B1(new_n1022), .B2(new_n975), .ZN(new_n1023));
  INV_X1    g598(.A(new_n956), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n1001), .B(new_n1011), .C1(new_n1023), .C2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT62), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT51), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n741), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n967), .A2(new_n968), .A3(new_n763), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1027), .B1(new_n1030), .B2(G286), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1028), .A2(G168), .A3(new_n1029), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(G8), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1027), .B1(new_n1032), .B2(G8), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1026), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1035), .ZN(new_n1037));
  AOI21_X1  g612(.A(G168), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1038));
  OAI211_X1 g613(.A(G8), .B(new_n1032), .C1(new_n1038), .C2(new_n1027), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1037), .A2(new_n1039), .A3(KEYINPUT62), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1025), .B1(new_n1036), .B2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n948), .B1(new_n969), .B2(new_n975), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(new_n1024), .ZN(new_n1043));
  AND2_X1   g618(.A1(new_n996), .A2(new_n999), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1043), .A2(new_n1044), .A3(new_n980), .ZN(new_n1045));
  NAND2_X1  g620(.A1(G168), .A2(G8), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1046), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1047), .B(KEYINPUT63), .C1(new_n1024), .C2(new_n1042), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1045), .A2(new_n1048), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n1001), .B(new_n1047), .C1(new_n1023), .C2(new_n1024), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT63), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1049), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NOR2_X1   g627(.A1(G305), .A2(G1981), .ZN(new_n1053));
  NOR2_X1   g628(.A1(G288), .A2(G1976), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1053), .B1(new_n996), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n977), .A2(G8), .ZN(new_n1056));
  OAI22_X1  g631(.A1(new_n1043), .A2(new_n1000), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  NOR3_X1   g632(.A1(new_n1041), .A2(new_n1052), .A3(new_n1057), .ZN(new_n1058));
  AOI21_X1  g633(.A(G1348), .B1(new_n967), .B2(new_n968), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n977), .A2(G2067), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n614), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  XOR2_X1   g637(.A(KEYINPUT56), .B(G2072), .Z(new_n1063));
  OR2_X1    g638(.A1(new_n974), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(G1956), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1065), .B1(new_n1012), .B2(new_n1015), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT120), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT119), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n564), .A2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n560), .A2(KEYINPUT119), .A3(new_n563), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1069), .A2(new_n570), .A3(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT57), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1067), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1070), .A2(new_n570), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT119), .B1(new_n560), .B2(new_n563), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n1067), .B(new_n1072), .C1(new_n1074), .C2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n565), .A2(KEYINPUT57), .A3(new_n570), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n1064), .B(new_n1066), .C1(new_n1073), .C2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1062), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT121), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1081), .B1(new_n1078), .B2(new_n1073), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1072), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(KEYINPUT120), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1084), .A2(KEYINPUT121), .A3(new_n1076), .A4(new_n1077), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1082), .A2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(G1956), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n974), .A2(new_n1063), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1086), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1080), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT123), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT61), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1093), .B1(new_n1094), .B2(new_n1086), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1092), .B1(new_n1095), .B2(new_n1079), .ZN(new_n1096));
  AND4_X1   g671(.A1(new_n1092), .A2(new_n1089), .A3(new_n1079), .A4(KEYINPUT61), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1078), .A2(new_n1073), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1099), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1079), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(new_n1093), .ZN(new_n1102));
  NOR3_X1   g677(.A1(new_n1059), .A2(new_n614), .A3(new_n1060), .ZN(new_n1103));
  OAI21_X1  g678(.A(KEYINPUT60), .B1(new_n1062), .B2(new_n1103), .ZN(new_n1104));
  XOR2_X1   g679(.A(KEYINPUT58), .B(G1341), .Z(new_n1105));
  XNOR2_X1  g680(.A(new_n1105), .B(KEYINPUT122), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n977), .A2(new_n1106), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n970), .A2(new_n940), .A3(new_n972), .A4(new_n973), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(new_n549), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(KEYINPUT59), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT59), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1109), .A2(new_n1112), .A3(new_n549), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n613), .A2(KEYINPUT60), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1102), .A2(new_n1104), .A3(new_n1114), .A4(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1091), .B1(new_n1098), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1022), .A2(new_n975), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(G8), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1045), .B1(new_n1121), .B2(new_n956), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT54), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n473), .A2(KEYINPUT53), .A3(G40), .A4(new_n753), .ZN(new_n1125));
  XNOR2_X1  g700(.A(new_n467), .B(KEYINPUT124), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1125), .B1(G2105), .B2(new_n1126), .ZN(new_n1127));
  AND2_X1   g702(.A1(new_n973), .A2(new_n1127), .ZN(new_n1128));
  AOI22_X1  g703(.A1(new_n1009), .A2(new_n1008), .B1(new_n1128), .B2(new_n933), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1124), .A2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1123), .B1(new_n1130), .B2(G171), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1005), .A2(new_n1010), .A3(G301), .ZN(new_n1132));
  AOI22_X1  g707(.A1(new_n1037), .A2(new_n1039), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  AND2_X1   g708(.A1(new_n1122), .A2(new_n1133), .ZN(new_n1134));
  AND3_X1   g709(.A1(new_n1124), .A2(new_n1129), .A3(G301), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1123), .B1(new_n1011), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT125), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  OAI211_X1 g713(.A(KEYINPUT125), .B(new_n1123), .C1(new_n1011), .C2(new_n1135), .ZN(new_n1139));
  AND2_X1   g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1119), .A2(new_n1134), .A3(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n947), .B1(new_n1058), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n943), .A2(new_n936), .ZN(new_n1143));
  XNOR2_X1  g718(.A(new_n1143), .B(KEYINPUT126), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n936), .A2(new_n797), .A3(new_n597), .ZN(new_n1145));
  XNOR2_X1  g720(.A(new_n1145), .B(KEYINPUT48), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n936), .A2(new_n940), .ZN(new_n1148));
  XNOR2_X1  g723(.A(new_n1148), .B(KEYINPUT46), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n938), .A2(new_n732), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(new_n936), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1152));
  XNOR2_X1  g727(.A(new_n1152), .B(KEYINPUT47), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n941), .A2(new_n790), .A3(new_n793), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1154), .B1(G2067), .B2(new_n817), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1155), .A2(new_n936), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1147), .A2(new_n1153), .A3(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n929), .B1(new_n1142), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1052), .ZN(new_n1159));
  NOR3_X1   g734(.A1(new_n1034), .A2(new_n1026), .A3(new_n1035), .ZN(new_n1160));
  AOI21_X1  g735(.A(KEYINPUT62), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1161));
  OAI211_X1 g736(.A(new_n1122), .B(new_n1011), .C1(new_n1160), .C2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1057), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1159), .A2(new_n1162), .A3(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT60), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1103), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1165), .B1(new_n1166), .B2(new_n1061), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1112), .B1(new_n1109), .B2(new_n549), .ZN(new_n1168));
  AOI211_X1 g743(.A(KEYINPUT59), .B(new_n548), .C1(new_n1107), .C2(new_n1108), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1117), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g745(.A(KEYINPUT61), .B1(new_n1079), .B2(new_n1100), .ZN(new_n1171));
  NOR3_X1   g746(.A1(new_n1167), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1089), .A2(new_n1079), .A3(KEYINPUT61), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1173), .A2(KEYINPUT123), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1095), .A2(new_n1092), .A3(new_n1079), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1090), .B1(new_n1172), .B2(new_n1176), .ZN(new_n1177));
  NAND4_X1  g752(.A1(new_n1122), .A2(new_n1133), .A3(new_n1138), .A4(new_n1139), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n946), .B1(new_n1164), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(new_n1157), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1180), .A2(KEYINPUT127), .A3(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1158), .A2(new_n1182), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g758(.A1(G229), .A2(new_n460), .A3(G401), .A4(G227), .ZN(new_n1185));
  NAND4_X1  g759(.A1(new_n924), .A2(new_n872), .A3(new_n926), .A4(new_n1185), .ZN(G225));
  INV_X1    g760(.A(G225), .ZN(G308));
endmodule


