//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 0 1 1 1 0 1 1 0 1 1 0 1 1 1 1 1 1 0 1 1 1 0 1 0 1 1 0 1 0 0 0 0 0 1 0 1 0 1 1 1 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:52 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n744, new_n745, new_n746, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n755, new_n756, new_n757,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n801,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n995, new_n996, new_n997, new_n998, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040;
  AND2_X1   g000(.A1(KEYINPUT70), .A2(G125), .ZN(new_n187));
  NOR2_X1   g001(.A1(KEYINPUT70), .A2(G125), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G143), .ZN(new_n191));
  INV_X1    g005(.A(G143), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G146), .ZN(new_n193));
  OR2_X1    g007(.A1(KEYINPUT0), .A2(G128), .ZN(new_n194));
  NAND2_X1  g008(.A1(KEYINPUT0), .A2(G128), .ZN(new_n195));
  AOI22_X1  g009(.A1(new_n191), .A2(new_n193), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  AND3_X1   g010(.A1(new_n191), .A2(new_n193), .A3(new_n195), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n189), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G953), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G224), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT83), .ZN(new_n201));
  XNOR2_X1  g015(.A(new_n200), .B(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT7), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT1), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n191), .A2(new_n193), .A3(new_n205), .A4(G128), .ZN(new_n206));
  INV_X1    g020(.A(new_n206), .ZN(new_n207));
  OAI21_X1  g021(.A(KEYINPUT1), .B1(new_n192), .B2(G146), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(KEYINPUT64), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT64), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n191), .A2(new_n210), .A3(KEYINPUT1), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n209), .A2(G128), .A3(new_n211), .ZN(new_n212));
  XNOR2_X1  g026(.A(G143), .B(G146), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n207), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  OAI211_X1 g029(.A(new_n198), .B(new_n204), .C1(new_n215), .C2(new_n189), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  XNOR2_X1  g031(.A(KEYINPUT70), .B(G125), .ZN(new_n218));
  INV_X1    g032(.A(G128), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n219), .B1(new_n208), .B2(KEYINPUT64), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n213), .B1(new_n220), .B2(new_n211), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n218), .B1(new_n221), .B2(new_n207), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n204), .B1(new_n222), .B2(new_n198), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n217), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g038(.A(G110), .B(G122), .ZN(new_n225));
  XNOR2_X1  g039(.A(new_n225), .B(KEYINPUT8), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G107), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n228), .A2(G104), .ZN(new_n229));
  INV_X1    g043(.A(G104), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n230), .A2(G107), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT75), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n232), .A2(KEYINPUT3), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n229), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  XOR2_X1   g048(.A(KEYINPUT76), .B(G101), .Z(new_n235));
  INV_X1    g049(.A(KEYINPUT3), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(KEYINPUT75), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n236), .A2(KEYINPUT75), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n228), .A2(G104), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n237), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n234), .A2(new_n235), .A3(new_n240), .ZN(new_n241));
  OAI21_X1  g055(.A(G101), .B1(new_n231), .B2(new_n229), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(G116), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n244), .A2(G119), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT65), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(new_n244), .ZN(new_n247));
  NAND2_X1  g061(.A1(KEYINPUT65), .A2(G116), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n245), .B1(new_n249), .B2(G119), .ZN(new_n250));
  XOR2_X1   g064(.A(KEYINPUT2), .B(G113), .Z(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n245), .ZN(new_n254));
  OAI21_X1  g068(.A(G113), .B1(new_n254), .B2(KEYINPUT5), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n255), .B1(new_n250), .B2(KEYINPUT5), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n243), .B1(new_n253), .B2(new_n256), .ZN(new_n257));
  AND2_X1   g071(.A1(KEYINPUT65), .A2(G116), .ZN(new_n258));
  NOR2_X1   g072(.A1(KEYINPUT65), .A2(G116), .ZN(new_n259));
  OAI21_X1  g073(.A(G119), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n260), .A2(KEYINPUT5), .A3(new_n254), .ZN(new_n261));
  OAI211_X1 g075(.A(new_n261), .B(G113), .C1(KEYINPUT5), .C2(new_n254), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n262), .A2(new_n252), .A3(new_n242), .A4(new_n241), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n227), .B1(new_n257), .B2(new_n263), .ZN(new_n264));
  OAI21_X1  g078(.A(KEYINPUT84), .B1(new_n224), .B2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(G101), .ZN(new_n266));
  AOI211_X1 g080(.A(KEYINPUT4), .B(new_n266), .C1(new_n234), .C2(new_n240), .ZN(new_n267));
  AND2_X1   g081(.A1(new_n241), .A2(KEYINPUT4), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n266), .B1(new_n234), .B2(new_n240), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n267), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n260), .A2(new_n254), .ZN(new_n272));
  XNOR2_X1  g086(.A(new_n272), .B(new_n251), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n271), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n275), .A2(new_n225), .A3(new_n263), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n257), .A2(new_n263), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(new_n226), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n198), .B1(new_n215), .B2(new_n189), .ZN(new_n279));
  INV_X1    g093(.A(new_n204), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(new_n216), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT84), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n278), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n265), .A2(new_n276), .A3(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(G902), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(KEYINPUT85), .ZN(new_n288));
  AND3_X1   g102(.A1(new_n275), .A2(new_n225), .A3(new_n263), .ZN(new_n289));
  XNOR2_X1  g103(.A(new_n225), .B(KEYINPUT82), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n290), .B1(new_n275), .B2(new_n263), .ZN(new_n291));
  OAI21_X1  g105(.A(KEYINPUT6), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT6), .ZN(new_n293));
  AND2_X1   g107(.A1(new_n275), .A2(new_n263), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n293), .B1(new_n294), .B2(new_n290), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n292), .A2(new_n295), .ZN(new_n296));
  XNOR2_X1  g110(.A(new_n279), .B(new_n202), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(G210), .B1(G237), .B2(G902), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT85), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n285), .A2(new_n301), .A3(new_n286), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n288), .A2(new_n299), .A3(new_n300), .A4(new_n302), .ZN(new_n303));
  AND3_X1   g117(.A1(new_n285), .A2(new_n301), .A3(new_n286), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n301), .B1(new_n285), .B2(new_n286), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n297), .B1(new_n292), .B2(new_n295), .ZN(new_n306));
  NOR3_X1   g120(.A1(new_n304), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  XNOR2_X1  g121(.A(new_n300), .B(KEYINPUT86), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n303), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(G214), .B1(G237), .B2(G902), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(KEYINPUT87), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT87), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n309), .A2(new_n313), .A3(new_n310), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT11), .ZN(new_n316));
  INV_X1    g130(.A(G134), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n316), .B1(new_n317), .B2(G137), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(G137), .ZN(new_n319));
  INV_X1    g133(.A(G137), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n320), .A2(KEYINPUT11), .A3(G134), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n318), .A2(new_n319), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G131), .ZN(new_n323));
  INV_X1    g137(.A(G131), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n318), .A2(new_n321), .A3(new_n324), .A4(new_n319), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n213), .A2(new_n195), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT66), .ZN(new_n328));
  AND2_X1   g142(.A1(new_n194), .A2(new_n195), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n327), .B(new_n328), .C1(new_n329), .C2(new_n213), .ZN(new_n330));
  OAI21_X1  g144(.A(KEYINPUT66), .B1(new_n196), .B2(new_n197), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n326), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n320), .A2(G134), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n317), .A2(G137), .ZN(new_n334));
  OAI21_X1  g148(.A(G131), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  AND2_X1   g149(.A1(new_n325), .A2(new_n335), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n336), .B1(new_n221), .B2(new_n207), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n332), .A2(new_n273), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(KEYINPUT28), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT28), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n332), .A2(new_n273), .A3(new_n337), .A4(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n327), .B1(new_n329), .B2(new_n213), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n326), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n337), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(new_n274), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n342), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(G237), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n348), .A2(new_n199), .A3(G210), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT27), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n349), .B(new_n350), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n351), .B(KEYINPUT26), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n352), .B(new_n266), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n347), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(new_n338), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n332), .A2(new_n337), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(KEYINPUT30), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT30), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n337), .A2(new_n359), .A3(new_n344), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n356), .B1(new_n361), .B2(new_n274), .ZN(new_n362));
  AOI21_X1  g176(.A(KEYINPUT31), .B1(new_n362), .B2(new_n353), .ZN(new_n363));
  AND3_X1   g177(.A1(new_n337), .A2(new_n359), .A3(new_n344), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n359), .B1(new_n332), .B2(new_n337), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n274), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n366), .A2(new_n353), .A3(KEYINPUT31), .A4(new_n338), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n355), .B1(new_n363), .B2(new_n368), .ZN(new_n369));
  NOR2_X1   g183(.A1(G472), .A2(G902), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n369), .A2(KEYINPUT67), .A3(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT67), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n366), .A2(new_n338), .A3(new_n353), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT31), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  AOI22_X1  g189(.A1(new_n375), .A2(new_n367), .B1(new_n347), .B2(new_n354), .ZN(new_n376));
  INV_X1    g190(.A(new_n370), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n372), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n371), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT32), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(G472), .ZN(new_n382));
  XOR2_X1   g196(.A(KEYINPUT68), .B(G902), .Z(new_n383));
  INV_X1    g197(.A(KEYINPUT29), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n354), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n357), .A2(new_n274), .ZN(new_n386));
  AND2_X1   g200(.A1(new_n342), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n383), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n342), .A2(new_n346), .A3(new_n353), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n389), .B(new_n384), .C1(new_n362), .C2(new_n353), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n382), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n376), .A2(new_n377), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n391), .B1(new_n392), .B2(KEYINPUT32), .ZN(new_n393));
  INV_X1    g207(.A(G217), .ZN(new_n394));
  INV_X1    g208(.A(new_n383), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n394), .B1(new_n395), .B2(G234), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n219), .A2(G119), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT23), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(G119), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(G128), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n219), .A2(KEYINPUT23), .A3(G119), .ZN(new_n403));
  AND3_X1   g217(.A1(new_n400), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(G110), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  XNOR2_X1  g220(.A(KEYINPUT24), .B(G110), .ZN(new_n407));
  AND3_X1   g221(.A1(new_n402), .A2(new_n398), .A3(KEYINPUT69), .ZN(new_n408));
  AOI21_X1  g222(.A(KEYINPUT69), .B1(new_n402), .B2(new_n398), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n407), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n406), .A2(new_n410), .ZN(new_n411));
  XNOR2_X1  g225(.A(G125), .B(G140), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(new_n190), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n413), .B(KEYINPUT72), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT16), .ZN(new_n415));
  INV_X1    g229(.A(G140), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n189), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  NOR2_X1   g231(.A1(G125), .A2(G140), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n418), .B1(new_n189), .B2(G140), .ZN(new_n419));
  OAI211_X1 g233(.A(G146), .B(new_n417), .C1(new_n419), .C2(new_n415), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n411), .A2(new_n414), .A3(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT73), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  OR2_X1    g237(.A1(KEYINPUT70), .A2(G125), .ZN(new_n424));
  NAND2_X1  g238(.A1(KEYINPUT70), .A2(G125), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n424), .A2(G140), .A3(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n418), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n415), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NOR3_X1   g242(.A1(new_n218), .A2(KEYINPUT16), .A3(G140), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n190), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n430), .A2(new_n420), .A3(KEYINPUT71), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT71), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n432), .B(new_n190), .C1(new_n428), .C2(new_n429), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n404), .A2(new_n405), .ZN(new_n434));
  NOR3_X1   g248(.A1(new_n408), .A2(new_n409), .A3(new_n407), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n431), .A2(new_n433), .A3(new_n436), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n411), .A2(new_n414), .A3(KEYINPUT73), .A4(new_n420), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n423), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n199), .A2(G221), .A3(G234), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n440), .B(KEYINPUT22), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n441), .B(G137), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n439), .A2(new_n443), .ZN(new_n444));
  NAND4_X1  g258(.A1(new_n423), .A2(new_n437), .A3(new_n438), .A4(new_n442), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n444), .A2(new_n395), .A3(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT25), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n444), .A2(KEYINPUT25), .A3(new_n395), .A4(new_n445), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n397), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  AND2_X1   g264(.A1(new_n444), .A2(new_n445), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n396), .A2(G902), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(KEYINPUT74), .B1(new_n450), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n448), .A2(new_n449), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(new_n396), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT74), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n457), .A2(new_n458), .A3(new_n453), .ZN(new_n459));
  AOI22_X1  g273(.A1(new_n381), .A2(new_n393), .B1(new_n455), .B2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(G475), .ZN(new_n461));
  XNOR2_X1  g275(.A(G113), .B(G122), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n462), .B(new_n230), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n431), .A2(new_n433), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n348), .A2(new_n199), .A3(G214), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n466), .B(G143), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT17), .ZN(new_n468));
  NOR3_X1   g282(.A1(new_n467), .A2(new_n468), .A3(new_n324), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(KEYINPUT91), .B1(new_n465), .B2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT91), .ZN(new_n472));
  AOI211_X1 g286(.A(new_n472), .B(new_n469), .C1(new_n431), .C2(new_n433), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT89), .ZN(new_n474));
  INV_X1    g288(.A(new_n467), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n474), .B1(new_n475), .B2(G131), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(G131), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n467), .A2(KEYINPUT89), .A3(new_n324), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n479), .A2(KEYINPUT17), .ZN(new_n480));
  NOR3_X1   g294(.A1(new_n471), .A2(new_n473), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n419), .A2(G146), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n482), .B(KEYINPUT88), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(new_n414), .ZN(new_n484));
  NAND2_X1  g298(.A1(KEYINPUT18), .A2(G131), .ZN(new_n485));
  XOR2_X1   g299(.A(new_n467), .B(new_n485), .Z(new_n486));
  NAND2_X1  g300(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n464), .B1(new_n481), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n465), .A2(new_n470), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(new_n472), .ZN(new_n491));
  INV_X1    g305(.A(new_n480), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n465), .A2(KEYINPUT91), .A3(new_n470), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n491), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n494), .A2(new_n463), .A3(new_n487), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n489), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n461), .B1(new_n496), .B2(new_n286), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n419), .A2(KEYINPUT19), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT19), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n412), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n498), .A2(new_n190), .A3(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT90), .ZN(new_n502));
  OR2_X1    g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n501), .A2(new_n502), .ZN(new_n504));
  AND4_X1   g318(.A1(new_n420), .A2(new_n503), .A3(new_n479), .A4(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n464), .B1(new_n488), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n495), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g321(.A1(G475), .A2(G902), .ZN(new_n508));
  AOI21_X1  g322(.A(KEYINPUT20), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT20), .ZN(new_n510));
  INV_X1    g324(.A(new_n508), .ZN(new_n511));
  AOI211_X1 g325(.A(new_n510), .B(new_n511), .C1(new_n495), .C2(new_n506), .ZN(new_n512));
  NOR3_X1   g326(.A1(new_n497), .A2(new_n509), .A3(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(G478), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n514), .A2(KEYINPUT15), .ZN(new_n515));
  XOR2_X1   g329(.A(KEYINPUT9), .B(G234), .Z(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  NOR3_X1   g331(.A1(new_n517), .A2(new_n394), .A3(G953), .ZN(new_n518));
  OAI21_X1  g332(.A(G122), .B1(new_n258), .B2(new_n259), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n519), .B1(new_n244), .B2(G122), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n520), .A2(G107), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT95), .ZN(new_n522));
  INV_X1    g336(.A(G122), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n523), .B1(new_n247), .B2(new_n248), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT14), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n522), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n244), .A2(G122), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n527), .B1(new_n524), .B2(new_n525), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n519), .A2(KEYINPUT95), .A3(KEYINPUT14), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n526), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n521), .B1(new_n530), .B2(G107), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n192), .A2(G128), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT92), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n533), .A2(new_n192), .A3(G128), .ZN(new_n534));
  OAI21_X1  g348(.A(KEYINPUT92), .B1(new_n219), .B2(G143), .ZN(new_n535));
  AOI211_X1 g349(.A(G134), .B(new_n532), .C1(new_n534), .C2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n534), .ZN(new_n537));
  INV_X1    g351(.A(new_n532), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n317), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(KEYINPUT94), .B1(new_n536), .B2(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n533), .B1(G128), .B2(new_n192), .ZN(new_n541));
  NOR3_X1   g355(.A1(new_n219), .A2(KEYINPUT92), .A3(G143), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n538), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(G134), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n537), .A2(new_n317), .A3(new_n538), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT94), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n540), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n531), .A2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT96), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n531), .A2(new_n548), .A3(KEYINPUT96), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n520), .B(G107), .ZN(new_n554));
  AOI21_X1  g368(.A(KEYINPUT13), .B1(new_n535), .B2(new_n534), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT93), .ZN(new_n556));
  OR3_X1    g370(.A1(new_n555), .A2(new_n556), .A3(new_n532), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n535), .A2(new_n534), .A3(KEYINPUT13), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n556), .B1(new_n555), .B2(new_n532), .ZN(new_n559));
  AND3_X1   g373(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n545), .B(new_n554), .C1(new_n560), .C2(new_n317), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n518), .B1(new_n553), .B2(new_n561), .ZN(new_n562));
  AND3_X1   g376(.A1(new_n531), .A2(KEYINPUT96), .A3(new_n548), .ZN(new_n563));
  AOI21_X1  g377(.A(KEYINPUT96), .B1(new_n531), .B2(new_n548), .ZN(new_n564));
  OAI211_X1 g378(.A(new_n561), .B(new_n518), .C1(new_n563), .C2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n395), .B1(new_n562), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT97), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n515), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n561), .B1(new_n563), .B2(new_n564), .ZN(new_n570));
  INV_X1    g384(.A(new_n518), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n383), .B1(new_n572), .B2(new_n565), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n573), .B(KEYINPUT97), .C1(KEYINPUT15), .C2(new_n514), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n569), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(G234), .A2(G237), .ZN(new_n577));
  AND3_X1   g391(.A1(new_n577), .A2(G952), .A3(new_n199), .ZN(new_n578));
  AND3_X1   g392(.A1(new_n383), .A2(G953), .A3(new_n577), .ZN(new_n579));
  XOR2_X1   g393(.A(KEYINPUT21), .B(G898), .Z(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n578), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n513), .A2(new_n576), .A3(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT79), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n585), .A2(KEYINPUT12), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n585), .A2(KEYINPUT12), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n219), .B1(new_n191), .B2(KEYINPUT1), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n206), .B1(new_n589), .B2(new_n213), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n241), .A2(new_n242), .A3(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT77), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n241), .A2(new_n590), .A3(KEYINPUT77), .A4(new_n242), .ZN(new_n594));
  AOI22_X1  g408(.A1(new_n593), .A2(new_n594), .B1(new_n215), .B2(new_n243), .ZN(new_n595));
  INV_X1    g409(.A(new_n326), .ZN(new_n596));
  OAI211_X1 g410(.A(new_n587), .B(new_n588), .C1(new_n595), .C2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n593), .A2(new_n594), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n215), .A2(new_n243), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n600), .A2(new_n326), .A3(new_n586), .ZN(new_n601));
  AND2_X1   g415(.A1(new_n597), .A2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT10), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n598), .A2(new_n603), .ZN(new_n604));
  AND2_X1   g418(.A1(new_n241), .A2(new_n242), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n212), .A2(new_n214), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(new_n206), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT78), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n605), .A2(new_n607), .A3(new_n608), .A4(KEYINPUT10), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n241), .A2(KEYINPUT10), .A3(new_n242), .ZN(new_n610));
  OAI21_X1  g424(.A(KEYINPUT78), .B1(new_n610), .B2(new_n215), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n268), .A2(new_n270), .ZN(new_n613));
  AND2_X1   g427(.A1(new_n330), .A2(new_n331), .ZN(new_n614));
  INV_X1    g428(.A(new_n267), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n604), .A2(new_n612), .A3(new_n596), .A4(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(G110), .B(G140), .ZN(new_n618));
  AND2_X1   g432(.A1(new_n199), .A2(G227), .ZN(new_n619));
  XOR2_X1   g433(.A(new_n618), .B(new_n619), .Z(new_n620));
  NAND4_X1  g434(.A1(new_n602), .A2(KEYINPUT81), .A3(new_n617), .A4(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n620), .ZN(new_n622));
  INV_X1    g436(.A(new_n617), .ZN(new_n623));
  AOI22_X1  g437(.A1(new_n603), .A2(new_n598), .B1(new_n271), .B2(new_n614), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n596), .B1(new_n624), .B2(new_n612), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n622), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n617), .A2(new_n597), .A3(new_n601), .A4(new_n620), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT81), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n621), .A2(new_n626), .A3(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(G469), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n630), .A2(new_n631), .A3(new_n395), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n617), .A2(new_n597), .A3(new_n601), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(KEYINPUT80), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT80), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n617), .A2(new_n597), .A3(new_n601), .A4(new_n635), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n620), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n620), .B1(new_n623), .B2(new_n625), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  OAI21_X1  g453(.A(G469), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(G469), .A2(G902), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n632), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  OAI21_X1  g456(.A(G221), .B1(new_n517), .B2(G902), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n584), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n315), .A2(new_n460), .A3(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(KEYINPUT98), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(new_n235), .ZN(G3));
  NAND2_X1  g462(.A1(new_n459), .A2(new_n455), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n382), .B1(new_n369), .B2(new_n395), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n650), .B1(new_n378), .B2(new_n371), .ZN(new_n651));
  AND4_X1   g465(.A1(new_n649), .A2(new_n651), .A3(new_n642), .A4(new_n643), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n304), .A2(new_n305), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n300), .B1(new_n653), .B2(new_n299), .ZN(new_n654));
  INV_X1    g468(.A(new_n303), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n310), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n656), .A2(new_n582), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT33), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n658), .B1(new_n571), .B2(KEYINPUT99), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n660), .B1(new_n562), .B2(new_n566), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n572), .A2(new_n565), .A3(new_n659), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n383), .A2(new_n514), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n661), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT100), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n665), .B1(new_n573), .B2(G478), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT101), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n661), .A2(new_n665), .A3(new_n662), .A4(new_n663), .ZN(new_n669));
  AND3_X1   g483(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n668), .B1(new_n667), .B2(new_n669), .ZN(new_n671));
  NOR3_X1   g485(.A1(new_n670), .A2(new_n671), .A3(new_n513), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n652), .A2(new_n657), .A3(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(KEYINPUT34), .B(G104), .Z(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G6));
  NOR2_X1   g489(.A1(new_n509), .A2(new_n512), .ZN(new_n676));
  INV_X1    g490(.A(new_n497), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n676), .A2(new_n677), .A3(new_n575), .ZN(new_n678));
  NOR3_X1   g492(.A1(new_n656), .A2(new_n678), .A3(new_n582), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(new_n652), .ZN(new_n680));
  XOR2_X1   g494(.A(KEYINPUT35), .B(G107), .Z(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G9));
  NOR2_X1   g496(.A1(new_n443), .A2(KEYINPUT36), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n439), .B(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(new_n452), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n457), .A2(new_n685), .ZN(new_n686));
  AOI21_X1  g500(.A(KEYINPUT102), .B1(new_n651), .B2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n650), .ZN(new_n688));
  AND4_X1   g502(.A1(KEYINPUT102), .A2(new_n379), .A3(new_n688), .A4(new_n686), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n315), .A2(new_n690), .A3(new_n645), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(KEYINPUT37), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(new_n405), .ZN(G12));
  AOI21_X1  g507(.A(KEYINPUT32), .B1(new_n371), .B2(new_n378), .ZN(new_n694));
  INV_X1    g508(.A(new_n391), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n369), .A2(KEYINPUT32), .A3(new_n370), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n686), .B1(new_n694), .B2(new_n697), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n698), .A2(new_n644), .ZN(new_n699));
  INV_X1    g513(.A(new_n656), .ZN(new_n700));
  INV_X1    g514(.A(new_n579), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n701), .A2(G900), .ZN(new_n702));
  OR2_X1    g516(.A1(new_n702), .A2(KEYINPUT103), .ZN(new_n703));
  INV_X1    g517(.A(new_n578), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n702), .A2(KEYINPUT103), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n703), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n678), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n699), .A2(new_n700), .A3(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(KEYINPUT104), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(new_n219), .ZN(G30));
  OR2_X1    g525(.A1(new_n309), .A2(KEYINPUT38), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n309), .A2(KEYINPUT38), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(new_n373), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n353), .B1(new_n338), .B2(new_n386), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n286), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(G472), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n381), .A2(new_n696), .A3(new_n718), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n513), .A2(new_n576), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n714), .A2(new_n310), .A3(new_n719), .A4(new_n720), .ZN(new_n721));
  XOR2_X1   g535(.A(new_n706), .B(KEYINPUT39), .Z(new_n722));
  NOR2_X1   g536(.A1(new_n644), .A2(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT40), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NOR3_X1   g539(.A1(new_n644), .A2(KEYINPUT40), .A3(new_n722), .ZN(new_n726));
  NOR4_X1   g540(.A1(new_n721), .A2(new_n725), .A3(new_n686), .A4(new_n726), .ZN(new_n727));
  XOR2_X1   g541(.A(new_n727), .B(KEYINPUT105), .Z(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G143), .ZN(G45));
  NAND4_X1  g543(.A1(new_n699), .A2(new_n672), .A3(new_n700), .A4(new_n706), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G146), .ZN(G48));
  NAND2_X1  g545(.A1(new_n630), .A2(new_n395), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(G469), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n733), .A2(new_n643), .A3(new_n632), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(KEYINPUT106), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT106), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n733), .A2(new_n736), .A3(new_n643), .A4(new_n632), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n738), .A2(new_n460), .A3(new_n672), .A4(new_n657), .ZN(new_n739));
  XNOR2_X1  g553(.A(KEYINPUT41), .B(G113), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n739), .B(new_n740), .ZN(G15));
  NAND3_X1  g555(.A1(new_n679), .A2(new_n738), .A3(new_n460), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G116), .ZN(G18));
  NOR2_X1   g557(.A1(new_n584), .A2(new_n698), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n656), .A2(new_n734), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G119), .ZN(G21));
  NOR2_X1   g561(.A1(new_n450), .A2(new_n454), .ZN(new_n748));
  OAI22_X1  g562(.A1(new_n363), .A2(new_n368), .B1(new_n353), .B2(new_n387), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(new_n370), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n688), .A2(new_n748), .A3(new_n750), .ZN(new_n751));
  NOR3_X1   g565(.A1(new_n751), .A2(new_n513), .A3(new_n576), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n738), .A2(new_n657), .A3(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G122), .ZN(G24));
  NAND3_X1  g568(.A1(new_n688), .A2(new_n686), .A3(new_n750), .ZN(new_n755));
  INV_X1    g569(.A(new_n755), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n745), .A2(new_n672), .A3(new_n706), .A4(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G125), .ZN(G27));
  INV_X1    g572(.A(KEYINPUT109), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT42), .ZN(new_n760));
  AND3_X1   g574(.A1(new_n572), .A2(new_n565), .A3(new_n659), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n659), .B1(new_n572), .B2(new_n565), .ZN(new_n762));
  INV_X1    g576(.A(new_n663), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n761), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  AOI21_X1  g578(.A(KEYINPUT100), .B1(new_n567), .B2(new_n514), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n669), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(KEYINPUT101), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n676), .A2(new_n677), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n767), .A2(new_n768), .A3(new_n769), .A4(new_n706), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT108), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n771), .B1(new_n392), .B2(KEYINPUT32), .ZN(new_n772));
  OAI211_X1 g586(.A(KEYINPUT108), .B(new_n380), .C1(new_n376), .C2(new_n377), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n772), .A2(new_n393), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(new_n748), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n770), .A2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(new_n643), .ZN(new_n777));
  INV_X1    g591(.A(new_n310), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  OAI211_X1 g593(.A(new_n303), .B(new_n779), .C1(new_n307), .C2(new_n308), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n642), .A2(KEYINPUT107), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT107), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n632), .A2(new_n640), .A3(new_n782), .A4(new_n641), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n780), .B1(new_n781), .B2(new_n783), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n760), .B1(new_n776), .B2(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n672), .A2(new_n760), .A3(new_n706), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n781), .A2(new_n783), .ZN(new_n787));
  INV_X1    g601(.A(new_n780), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n787), .A2(new_n460), .A3(new_n788), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n786), .A2(new_n789), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n759), .B1(new_n785), .B2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(new_n775), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n792), .A2(new_n672), .A3(new_n706), .ZN(new_n793));
  INV_X1    g607(.A(new_n784), .ZN(new_n794));
  OAI21_X1  g608(.A(KEYINPUT42), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(new_n770), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n796), .A2(new_n760), .A3(new_n784), .A4(new_n460), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n795), .A2(KEYINPUT109), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n791), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G131), .ZN(G33));
  NAND3_X1  g614(.A1(new_n784), .A2(new_n460), .A3(new_n708), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G134), .ZN(G36));
  NOR2_X1   g616(.A1(new_n309), .A2(new_n778), .ZN(new_n803));
  INV_X1    g617(.A(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n686), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n670), .A2(new_n671), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(new_n513), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT43), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n806), .A2(KEYINPUT43), .A3(new_n513), .ZN(new_n810));
  AOI211_X1 g624(.A(new_n651), .B(new_n805), .C1(new_n809), .C2(new_n810), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n804), .B1(new_n811), .B2(KEYINPUT44), .ZN(new_n812));
  OR3_X1    g626(.A1(new_n637), .A2(KEYINPUT45), .A3(new_n639), .ZN(new_n813));
  OAI21_X1  g627(.A(KEYINPUT45), .B1(new_n637), .B2(new_n639), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n813), .A2(G469), .A3(new_n814), .ZN(new_n815));
  AOI21_X1  g629(.A(KEYINPUT46), .B1(new_n815), .B2(new_n641), .ZN(new_n816));
  INV_X1    g630(.A(new_n632), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n815), .A2(KEYINPUT46), .A3(new_n641), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(new_n643), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n821), .A2(new_n722), .ZN(new_n822));
  OAI211_X1 g636(.A(new_n812), .B(new_n822), .C1(KEYINPUT44), .C2(new_n811), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(G137), .ZN(G39));
  NOR2_X1   g638(.A1(new_n821), .A2(KEYINPUT47), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT47), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n826), .B1(new_n820), .B2(new_n643), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  NOR4_X1   g642(.A1(new_n770), .A2(new_n649), .A3(new_n694), .A4(new_n697), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n828), .A2(new_n803), .A3(new_n829), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n830), .B(G140), .ZN(G42));
  OR2_X1    g645(.A1(new_n719), .A2(new_n704), .ZN(new_n832));
  INV_X1    g646(.A(new_n734), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n833), .A2(new_n803), .A3(new_n649), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n767), .A2(new_n768), .A3(new_n769), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n832), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n809), .A2(new_n810), .ZN(new_n837));
  AND4_X1   g651(.A1(new_n578), .A2(new_n837), .A3(new_n833), .A4(new_n803), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(new_n792), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n839), .B(KEYINPUT48), .ZN(new_n840));
  INV_X1    g654(.A(G952), .ZN(new_n841));
  AOI211_X1 g655(.A(new_n704), .B(new_n751), .C1(new_n809), .C2(new_n810), .ZN(new_n842));
  AOI211_X1 g656(.A(new_n841), .B(G953), .C1(new_n842), .C2(new_n745), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n733), .A2(new_n632), .ZN(new_n845));
  OAI22_X1  g659(.A1(new_n825), .A2(new_n827), .B1(new_n643), .B2(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n846), .A2(new_n803), .A3(new_n842), .ZN(new_n847));
  NOR4_X1   g661(.A1(new_n832), .A2(new_n834), .A3(new_n768), .A4(new_n806), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n712), .A2(new_n833), .A3(new_n778), .A4(new_n713), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n849), .B(KEYINPUT113), .ZN(new_n850));
  INV_X1    g664(.A(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT114), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT50), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n851), .A2(new_n842), .A3(new_n854), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n852), .A2(new_n853), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n848), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n838), .A2(new_n756), .ZN(new_n858));
  INV_X1    g672(.A(new_n856), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n851), .A2(new_n842), .A3(new_n859), .A4(new_n854), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n847), .A2(new_n857), .A3(new_n858), .A4(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT115), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT51), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n861), .A2(new_n862), .A3(new_n868), .ZN(new_n869));
  AOI211_X1 g683(.A(new_n836), .B(new_n844), .C1(new_n865), .C2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT112), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT54), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT52), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n730), .A2(new_n757), .A3(new_n709), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n656), .A2(new_n576), .A3(new_n513), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(new_n787), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n719), .A2(new_n643), .A3(new_n805), .A4(new_n706), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n873), .B1(new_n874), .B2(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n770), .A2(new_n755), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n698), .A2(new_n656), .A3(new_n644), .ZN(new_n881));
  AOI22_X1  g695(.A1(new_n745), .A2(new_n880), .B1(new_n881), .B2(new_n708), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n719), .A2(new_n805), .A3(new_n706), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n883), .A2(new_n643), .A3(new_n787), .A4(new_n875), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n882), .A2(KEYINPUT52), .A3(new_n730), .A4(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n879), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n835), .A2(new_n678), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n315), .A2(new_n887), .A3(new_n583), .A4(new_n652), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n888), .A2(new_n691), .A3(new_n739), .A4(new_n742), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n646), .A2(new_n746), .A3(new_n753), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n768), .A2(new_n575), .A3(new_n707), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n699), .A2(new_n803), .A3(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n672), .A2(new_n706), .A3(new_n756), .ZN(new_n893));
  OAI211_X1 g707(.A(new_n801), .B(new_n892), .C1(new_n893), .C2(new_n794), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n889), .A2(new_n890), .A3(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n785), .A2(new_n790), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n886), .A2(new_n895), .A3(KEYINPUT53), .A4(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n886), .A2(new_n895), .A3(new_n799), .ZN(new_n898));
  XNOR2_X1  g712(.A(KEYINPUT110), .B(KEYINPUT53), .ZN(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  AND3_X1   g714(.A1(new_n898), .A2(KEYINPUT111), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(KEYINPUT111), .B1(new_n898), .B2(new_n900), .ZN(new_n902));
  OAI211_X1 g716(.A(new_n872), .B(new_n897), .C1(new_n901), .C2(new_n902), .ZN(new_n903));
  OR2_X1    g717(.A1(new_n898), .A2(new_n899), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n898), .A2(KEYINPUT53), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n904), .A2(KEYINPUT54), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n871), .B1(new_n903), .B2(new_n906), .ZN(new_n907));
  AND3_X1   g721(.A1(new_n903), .A2(new_n871), .A3(new_n906), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n870), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT116), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n841), .A2(new_n199), .ZN(new_n912));
  OAI211_X1 g726(.A(new_n870), .B(KEYINPUT116), .C1(new_n907), .C2(new_n908), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  OR2_X1    g728(.A1(new_n845), .A2(KEYINPUT49), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n845), .A2(KEYINPUT49), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n915), .A2(new_n748), .A3(new_n779), .A4(new_n916), .ZN(new_n917));
  OR4_X1    g731(.A1(new_n719), .A2(new_n917), .A3(new_n714), .A4(new_n807), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n914), .A2(new_n918), .ZN(G75));
  NOR2_X1   g733(.A1(new_n296), .A2(new_n298), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n920), .A2(new_n306), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT117), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT55), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n898), .A2(new_n900), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT111), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n898), .A2(KEYINPUT111), .A3(new_n900), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n395), .B1(new_n928), .B2(new_n897), .ZN(new_n929));
  INV_X1    g743(.A(new_n300), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT56), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n923), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n199), .A2(G952), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n923), .A2(new_n932), .ZN(new_n935));
  INV_X1    g749(.A(new_n308), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n935), .B1(new_n929), .B2(new_n936), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n933), .A2(new_n934), .A3(new_n937), .ZN(G51));
  INV_X1    g752(.A(new_n815), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n929), .A2(new_n939), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(KEYINPUT119), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n630), .B(KEYINPUT118), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n897), .B1(new_n901), .B2(new_n902), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(KEYINPUT54), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(new_n903), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n641), .B(KEYINPUT57), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n942), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n934), .B1(new_n941), .B2(new_n948), .ZN(G54));
  NAND3_X1  g763(.A1(new_n929), .A2(KEYINPUT58), .A3(G475), .ZN(new_n950));
  INV_X1    g764(.A(new_n507), .ZN(new_n951));
  AND3_X1   g765(.A1(new_n950), .A2(KEYINPUT120), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(KEYINPUT120), .B1(new_n950), .B2(new_n951), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n950), .A2(new_n951), .ZN(new_n954));
  NOR4_X1   g768(.A1(new_n952), .A2(new_n953), .A3(new_n954), .A4(new_n934), .ZN(G60));
  INV_X1    g769(.A(KEYINPUT122), .ZN(new_n956));
  INV_X1    g770(.A(new_n934), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT121), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n761), .A2(new_n762), .ZN(new_n959));
  NAND2_X1  g773(.A1(G478), .A2(G902), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(KEYINPUT59), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n958), .B1(new_n945), .B2(new_n963), .ZN(new_n964));
  AOI211_X1 g778(.A(KEYINPUT121), .B(new_n962), .C1(new_n944), .C2(new_n903), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n957), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n908), .A2(new_n907), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n959), .B1(new_n967), .B2(new_n961), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n956), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n903), .A2(new_n906), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(KEYINPUT112), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n903), .A2(new_n871), .A3(new_n906), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n971), .A2(new_n972), .A3(new_n961), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n973), .B1(new_n762), .B2(new_n761), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n872), .B1(new_n928), .B2(new_n897), .ZN(new_n975));
  INV_X1    g789(.A(new_n903), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n963), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(KEYINPUT121), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n945), .A2(new_n958), .A3(new_n963), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND4_X1  g794(.A1(new_n974), .A2(new_n980), .A3(KEYINPUT122), .A4(new_n957), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n969), .A2(new_n981), .ZN(G63));
  NAND2_X1  g796(.A1(G217), .A2(G902), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n983), .B(KEYINPUT60), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n984), .B1(new_n928), .B2(new_n897), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n985), .A2(new_n684), .ZN(new_n986));
  OAI211_X1 g800(.A(new_n986), .B(new_n957), .C1(new_n451), .C2(new_n985), .ZN(new_n987));
  XNOR2_X1  g801(.A(KEYINPUT123), .B(KEYINPUT61), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT124), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n987), .A2(KEYINPUT124), .A3(new_n988), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT61), .ZN(new_n993));
  OAI211_X1 g807(.A(new_n991), .B(new_n992), .C1(new_n993), .C2(new_n987), .ZN(G66));
  AOI21_X1  g808(.A(new_n199), .B1(new_n580), .B2(G224), .ZN(new_n995));
  OR2_X1    g809(.A1(new_n889), .A2(new_n890), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n995), .B1(new_n996), .B2(new_n199), .ZN(new_n997));
  OAI211_X1 g811(.A(new_n292), .B(new_n295), .C1(G898), .C2(new_n199), .ZN(new_n998));
  XOR2_X1   g812(.A(new_n997), .B(new_n998), .Z(G69));
  AOI21_X1  g813(.A(new_n199), .B1(G227), .B2(G900), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n1000), .A2(KEYINPUT127), .ZN(new_n1001));
  INV_X1    g815(.A(new_n1000), .ZN(new_n1002));
  INV_X1    g816(.A(KEYINPUT127), .ZN(new_n1003));
  NOR2_X1   g817(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n498), .A2(new_n500), .ZN(new_n1005));
  XOR2_X1   g819(.A(new_n1005), .B(KEYINPUT125), .Z(new_n1006));
  XNOR2_X1  g820(.A(new_n361), .B(new_n1006), .ZN(new_n1007));
  INV_X1    g821(.A(new_n1007), .ZN(new_n1008));
  INV_X1    g822(.A(new_n460), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n835), .A2(KEYINPUT126), .A3(new_n678), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n1010), .A2(new_n723), .A3(new_n803), .ZN(new_n1011));
  INV_X1    g825(.A(KEYINPUT126), .ZN(new_n1012));
  AOI211_X1 g826(.A(new_n1009), .B(new_n1011), .C1(new_n1012), .C2(new_n887), .ZN(new_n1013));
  INV_X1    g827(.A(KEYINPUT62), .ZN(new_n1014));
  INV_X1    g828(.A(new_n728), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n1014), .B1(new_n1015), .B2(new_n874), .ZN(new_n1016));
  INV_X1    g830(.A(new_n874), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n728), .A2(KEYINPUT62), .A3(new_n1017), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1013), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1019));
  AND2_X1   g833(.A1(new_n823), .A2(new_n830), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n1008), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n822), .A2(new_n792), .A3(new_n875), .ZN(new_n1022));
  AND3_X1   g836(.A1(new_n1022), .A2(new_n801), .A3(new_n1017), .ZN(new_n1023));
  NAND3_X1  g837(.A1(new_n1020), .A2(new_n799), .A3(new_n1023), .ZN(new_n1024));
  AOI21_X1  g838(.A(new_n1007), .B1(new_n1024), .B2(new_n199), .ZN(new_n1025));
  OAI21_X1  g839(.A(new_n199), .B1(new_n1021), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1025), .A2(G900), .ZN(new_n1027));
  AOI211_X1 g841(.A(new_n1001), .B(new_n1004), .C1(new_n1026), .C2(new_n1027), .ZN(new_n1028));
  AND4_X1   g842(.A1(new_n1003), .A2(new_n1026), .A3(new_n1002), .A4(new_n1027), .ZN(new_n1029));
  NOR2_X1   g843(.A1(new_n1028), .A2(new_n1029), .ZN(G72));
  NAND2_X1  g844(.A1(G472), .A2(G902), .ZN(new_n1031));
  XOR2_X1   g845(.A(new_n1031), .B(KEYINPUT63), .Z(new_n1032));
  NAND2_X1  g846(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1033));
  OAI211_X1 g847(.A(new_n353), .B(new_n1032), .C1(new_n1033), .C2(new_n996), .ZN(new_n1034));
  NOR2_X1   g848(.A1(new_n362), .A2(new_n353), .ZN(new_n1035));
  NOR2_X1   g849(.A1(new_n1035), .A2(new_n715), .ZN(new_n1036));
  OAI211_X1 g850(.A(new_n354), .B(new_n1032), .C1(new_n1024), .C2(new_n996), .ZN(new_n1037));
  NAND3_X1  g851(.A1(new_n1034), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g852(.A(new_n1036), .ZN(new_n1039));
  NAND4_X1  g853(.A1(new_n904), .A2(new_n905), .A3(new_n1032), .A4(new_n1039), .ZN(new_n1040));
  AND3_X1   g854(.A1(new_n1038), .A2(new_n957), .A3(new_n1040), .ZN(G57));
endmodule


