

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759;

  NOR2_X1 U381 ( .A1(G953), .A2(G237), .ZN(n472) );
  XNOR2_X2 U382 ( .A(n407), .B(G469), .ZN(n542) );
  OR2_X2 U383 ( .A1(n626), .A2(G902), .ZN(n446) );
  NOR2_X1 U384 ( .A1(n663), .A2(n368), .ZN(n565) );
  INV_X1 U385 ( .A(n516), .ZN(n549) );
  XNOR2_X1 U386 ( .A(n369), .B(n359), .ZN(n516) );
  XNOR2_X1 U387 ( .A(n494), .B(n367), .ZN(n451) );
  XNOR2_X1 U388 ( .A(KEYINPUT70), .B(KEYINPUT4), .ZN(n367) );
  INV_X2 U389 ( .A(G953), .ZN(n747) );
  NOR2_X1 U390 ( .A1(n756), .A2(n759), .ZN(n373) );
  NOR2_X1 U391 ( .A1(n598), .A2(n597), .ZN(n606) );
  XNOR2_X1 U392 ( .A(n373), .B(n372), .ZN(n371) );
  NOR2_X1 U393 ( .A1(n504), .A2(KEYINPUT76), .ZN(n391) );
  NAND2_X1 U394 ( .A1(n618), .A2(n611), .ZN(n369) );
  XNOR2_X1 U395 ( .A(n417), .B(n416), .ZN(n422) );
  XOR2_X1 U396 ( .A(KEYINPUT24), .B(G110), .Z(n419) );
  INV_X1 U397 ( .A(G146), .ZN(n423) );
  XNOR2_X1 U398 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n454) );
  XNOR2_X1 U399 ( .A(KEYINPUT73), .B(G110), .ZN(n396) );
  NOR2_X1 U400 ( .A1(n693), .A2(n695), .ZN(n509) );
  INV_X1 U401 ( .A(KEYINPUT39), .ZN(n468) );
  NOR2_X1 U402 ( .A1(n657), .A2(n537), .ZN(n539) );
  AND2_X1 U403 ( .A1(n574), .A2(n360), .ZN(n393) );
  XNOR2_X1 U404 ( .A(n508), .B(KEYINPUT105), .ZN(n520) );
  BUF_X1 U405 ( .A(n555), .Z(n674) );
  AND2_X1 U406 ( .A1(n581), .A2(n575), .ZN(n595) );
  NOR2_X1 U407 ( .A1(n669), .A2(n668), .ZN(n670) );
  INV_X1 U408 ( .A(KEYINPUT46), .ZN(n372) );
  XNOR2_X1 U409 ( .A(n410), .B(n409), .ZN(n425) );
  XNOR2_X1 U410 ( .A(KEYINPUT20), .B(KEYINPUT90), .ZN(n409) );
  XNOR2_X1 U411 ( .A(G113), .B(G116), .ZN(n437) );
  XNOR2_X1 U412 ( .A(G143), .B(G140), .ZN(n470) );
  XNOR2_X1 U413 ( .A(n479), .B(n478), .ZN(n480) );
  INV_X1 U414 ( .A(G122), .ZN(n478) );
  XNOR2_X1 U415 ( .A(n395), .B(G101), .ZN(n441) );
  INV_X1 U416 ( .A(KEYINPUT68), .ZN(n395) );
  XOR2_X1 U417 ( .A(G113), .B(G104), .Z(n477) );
  XOR2_X1 U418 ( .A(KEYINPUT3), .B(G119), .Z(n461) );
  XNOR2_X1 U419 ( .A(G116), .B(G107), .ZN(n459) );
  XNOR2_X1 U420 ( .A(n549), .B(KEYINPUT38), .ZN(n690) );
  NOR2_X1 U421 ( .A1(n676), .A2(n504), .ZN(n380) );
  AND2_X1 U422 ( .A1(n502), .A2(n360), .ZN(n506) );
  INV_X1 U423 ( .A(KEYINPUT72), .ZN(n405) );
  XNOR2_X1 U424 ( .A(n502), .B(n538), .ZN(n574) );
  XNOR2_X1 U425 ( .A(KEYINPUT71), .B(KEYINPUT8), .ZN(n413) );
  XOR2_X1 U426 ( .A(G137), .B(G140), .Z(n401) );
  NAND2_X1 U427 ( .A1(n504), .A2(KEYINPUT76), .ZN(n387) );
  XNOR2_X1 U428 ( .A(n486), .B(n485), .ZN(n525) );
  XNOR2_X1 U429 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U430 ( .A(n564), .B(KEYINPUT0), .ZN(n590) );
  NOR2_X1 U431 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U432 ( .A(n376), .B(n375), .ZN(n724) );
  INV_X1 U433 ( .A(n424), .ZN(n375) );
  NAND2_X1 U434 ( .A1(n384), .A2(n365), .ZN(n383) );
  XNOR2_X1 U435 ( .A(n464), .B(n732), .ZN(n618) );
  XNOR2_X1 U436 ( .A(n512), .B(n511), .ZN(n756) );
  XNOR2_X1 U437 ( .A(n544), .B(KEYINPUT108), .ZN(n757) );
  NOR2_X1 U438 ( .A1(n546), .A2(n549), .ZN(n540) );
  XNOR2_X1 U439 ( .A(n370), .B(n364), .ZN(n583) );
  NOR2_X1 U440 ( .A1(n709), .A2(n708), .ZN(n710) );
  AND2_X2 U441 ( .A1(n383), .A2(n382), .ZN(n711) );
  XOR2_X1 U442 ( .A(n467), .B(KEYINPUT86), .Z(n359) );
  AND2_X1 U443 ( .A1(n503), .A2(n380), .ZN(n360) );
  NOR2_X1 U444 ( .A1(n389), .A2(n386), .ZN(n523) );
  XOR2_X1 U445 ( .A(n450), .B(n449), .Z(n361) );
  XOR2_X1 U446 ( .A(KEYINPUT83), .B(n757), .Z(n362) );
  AND2_X1 U447 ( .A1(n640), .A2(n662), .ZN(n363) );
  XOR2_X1 U448 ( .A(KEYINPUT65), .B(KEYINPUT32), .Z(n364) );
  XNOR2_X1 U449 ( .A(n408), .B(n497), .ZN(n611) );
  NAND2_X1 U450 ( .A1(n613), .A2(KEYINPUT67), .ZN(n365) );
  XOR2_X1 U451 ( .A(n633), .B(n632), .Z(n366) );
  AND2_X1 U452 ( .A1(n551), .A2(n640), .ZN(n381) );
  INV_X1 U453 ( .A(n668), .ZN(n382) );
  NOR2_X2 U454 ( .A1(n635), .A2(n726), .ZN(n636) );
  XNOR2_X2 U455 ( .A(n446), .B(G472), .ZN(n502) );
  XNOR2_X2 U456 ( .A(G143), .B(G128), .ZN(n494) );
  NOR2_X1 U457 ( .A1(n684), .A2(n368), .ZN(n587) );
  INV_X1 U458 ( .A(n590), .ZN(n368) );
  INV_X1 U459 ( .A(n583), .ZN(n643) );
  NAND2_X1 U460 ( .A1(n595), .A2(n577), .ZN(n370) );
  NOR2_X2 U461 ( .A1(n374), .A2(n371), .ZN(n545) );
  NAND2_X1 U462 ( .A1(n362), .A2(n536), .ZN(n374) );
  NAND2_X1 U463 ( .A1(n378), .A2(n377), .ZN(n376) );
  NAND2_X1 U464 ( .A1(n422), .A2(n421), .ZN(n377) );
  NAND2_X1 U465 ( .A1(n379), .A2(n420), .ZN(n378) );
  INV_X1 U466 ( .A(n422), .ZN(n379) );
  INV_X1 U467 ( .A(n503), .ZN(n576) );
  AND2_X1 U468 ( .A1(n551), .A2(n363), .ZN(n745) );
  NAND2_X1 U469 ( .A1(n381), .A2(n615), .ZN(n616) );
  NAND2_X1 U470 ( .A1(n385), .A2(n612), .ZN(n384) );
  OR2_X2 U471 ( .A1(n665), .A2(n610), .ZN(n385) );
  NAND2_X1 U472 ( .A1(n388), .A2(n387), .ZN(n386) );
  NAND2_X1 U473 ( .A1(n588), .A2(KEYINPUT76), .ZN(n388) );
  NAND2_X1 U474 ( .A1(n361), .A2(n390), .ZN(n389) );
  NAND2_X1 U475 ( .A1(n392), .A2(n391), .ZN(n390) );
  INV_X1 U476 ( .A(n588), .ZN(n392) );
  NAND2_X1 U477 ( .A1(n554), .A2(n542), .ZN(n588) );
  NAND2_X1 U478 ( .A1(n711), .A2(G478), .ZN(n721) );
  XNOR2_X1 U479 ( .A(n634), .B(n366), .ZN(n635) );
  NAND2_X1 U480 ( .A1(n711), .A2(G475), .ZN(n634) );
  XNOR2_X1 U481 ( .A(n469), .B(n468), .ZN(n553) );
  NOR2_X2 U482 ( .A1(n623), .A2(n726), .ZN(n624) );
  XOR2_X1 U483 ( .A(n626), .B(n625), .Z(n394) );
  NAND2_X1 U484 ( .A1(n552), .A2(n657), .ZN(n530) );
  INV_X1 U485 ( .A(n689), .ZN(n537) );
  XNOR2_X1 U486 ( .A(n480), .B(n424), .ZN(n481) );
  XNOR2_X1 U487 ( .A(KEYINPUT85), .B(KEYINPUT15), .ZN(n408) );
  INV_X1 U488 ( .A(KEYINPUT101), .ZN(n514) );
  INV_X1 U489 ( .A(n726), .ZN(n628) );
  INV_X1 U490 ( .A(n719), .ZN(n720) );
  XNOR2_X1 U491 ( .A(n660), .B(n514), .ZN(n552) );
  XNOR2_X1 U492 ( .A(n721), .B(n720), .ZN(n722) );
  INV_X1 U493 ( .A(n441), .ZN(n397) );
  XNOR2_X2 U494 ( .A(n397), .B(n396), .ZN(n452) );
  XOR2_X1 U495 ( .A(G104), .B(G107), .Z(n399) );
  NAND2_X1 U496 ( .A1(G227), .A2(n747), .ZN(n398) );
  XOR2_X1 U497 ( .A(n399), .B(n398), .Z(n400) );
  XNOR2_X1 U498 ( .A(n452), .B(n400), .ZN(n402) );
  XNOR2_X1 U499 ( .A(KEYINPUT89), .B(n401), .ZN(n739) );
  XNOR2_X1 U500 ( .A(n402), .B(n739), .ZN(n404) );
  XNOR2_X1 U501 ( .A(G131), .B(G134), .ZN(n403) );
  XNOR2_X1 U502 ( .A(n451), .B(n403), .ZN(n742) );
  XNOR2_X1 U503 ( .A(n742), .B(G146), .ZN(n444) );
  XNOR2_X1 U504 ( .A(n404), .B(n444), .ZN(n715) );
  NOR2_X1 U505 ( .A1(n715), .A2(G902), .ZN(n406) );
  XNOR2_X1 U506 ( .A(n406), .B(n405), .ZN(n407) );
  INV_X1 U507 ( .A(G902), .ZN(n497) );
  NAND2_X1 U508 ( .A1(n611), .A2(G234), .ZN(n410) );
  AND2_X1 U509 ( .A1(n425), .A2(G221), .ZN(n412) );
  INV_X1 U510 ( .A(KEYINPUT21), .ZN(n411) );
  XNOR2_X1 U511 ( .A(n412), .B(n411), .ZN(n676) );
  NAND2_X1 U512 ( .A1(n747), .A2(G234), .ZN(n414) );
  XNOR2_X1 U513 ( .A(n414), .B(n413), .ZN(n491) );
  NAND2_X1 U514 ( .A1(G221), .A2(n491), .ZN(n417) );
  XNOR2_X1 U515 ( .A(G137), .B(G140), .ZN(n415) );
  XNOR2_X1 U516 ( .A(n415), .B(KEYINPUT23), .ZN(n416) );
  XNOR2_X1 U517 ( .A(G128), .B(G119), .ZN(n418) );
  XNOR2_X1 U518 ( .A(n419), .B(n418), .ZN(n421) );
  INV_X1 U519 ( .A(n421), .ZN(n420) );
  XNOR2_X1 U520 ( .A(n423), .B(G125), .ZN(n456) );
  XOR2_X1 U521 ( .A(n456), .B(KEYINPUT10), .Z(n424) );
  NOR2_X1 U522 ( .A1(n724), .A2(G902), .ZN(n429) );
  XNOR2_X1 U523 ( .A(KEYINPUT91), .B(KEYINPUT25), .ZN(n427) );
  NAND2_X1 U524 ( .A1(G217), .A2(n425), .ZN(n426) );
  XNOR2_X1 U525 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U526 ( .A(n429), .B(n428), .ZN(n503) );
  NOR2_X1 U527 ( .A1(n676), .A2(n503), .ZN(n554) );
  XOR2_X1 U528 ( .A(KEYINPUT14), .B(KEYINPUT87), .Z(n431) );
  NAND2_X1 U529 ( .A1(G234), .A2(G237), .ZN(n430) );
  XNOR2_X1 U530 ( .A(n431), .B(n430), .ZN(n432) );
  NAND2_X1 U531 ( .A1(G952), .A2(n432), .ZN(n706) );
  NOR2_X1 U532 ( .A1(n706), .A2(G953), .ZN(n561) );
  NAND2_X1 U533 ( .A1(G902), .A2(n432), .ZN(n559) );
  OR2_X1 U534 ( .A1(n747), .A2(n559), .ZN(n433) );
  NOR2_X1 U535 ( .A1(G900), .A2(n433), .ZN(n434) );
  NOR2_X1 U536 ( .A1(n561), .A2(n434), .ZN(n504) );
  XOR2_X1 U537 ( .A(KEYINPUT30), .B(KEYINPUT103), .Z(n450) );
  XOR2_X1 U538 ( .A(KEYINPUT92), .B(KEYINPUT75), .Z(n436) );
  NAND2_X1 U539 ( .A1(n472), .A2(G210), .ZN(n435) );
  XNOR2_X1 U540 ( .A(n436), .B(n435), .ZN(n440) );
  XOR2_X1 U541 ( .A(G137), .B(KEYINPUT5), .Z(n438) );
  XNOR2_X1 U542 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U543 ( .A(n440), .B(n439), .Z(n443) );
  XNOR2_X1 U544 ( .A(n441), .B(n461), .ZN(n442) );
  XNOR2_X1 U545 ( .A(n443), .B(n442), .ZN(n445) );
  XNOR2_X1 U546 ( .A(n445), .B(n444), .ZN(n626) );
  NOR2_X1 U547 ( .A1(G237), .A2(G902), .ZN(n447) );
  XNOR2_X1 U548 ( .A(n447), .B(KEYINPUT74), .ZN(n466) );
  INV_X1 U549 ( .A(G214), .ZN(n448) );
  OR2_X1 U550 ( .A1(n466), .A2(n448), .ZN(n689) );
  NAND2_X1 U551 ( .A1(n502), .A2(n689), .ZN(n449) );
  XNOR2_X1 U552 ( .A(n452), .B(n451), .ZN(n458) );
  NAND2_X1 U553 ( .A1(n747), .A2(G224), .ZN(n453) );
  XNOR2_X1 U554 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U555 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U556 ( .A(n458), .B(n457), .ZN(n464) );
  XNOR2_X1 U557 ( .A(n459), .B(G122), .ZN(n490) );
  XNOR2_X1 U558 ( .A(n490), .B(n477), .ZN(n463) );
  INV_X1 U559 ( .A(KEYINPUT16), .ZN(n460) );
  XNOR2_X1 U560 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U561 ( .A(n463), .B(n462), .ZN(n732) );
  INV_X1 U562 ( .A(G210), .ZN(n465) );
  OR2_X1 U563 ( .A1(n466), .A2(n465), .ZN(n467) );
  NAND2_X1 U564 ( .A1(n523), .A2(n690), .ZN(n469) );
  XOR2_X1 U565 ( .A(KEYINPUT95), .B(KEYINPUT11), .Z(n471) );
  XNOR2_X1 U566 ( .A(n471), .B(n470), .ZN(n476) );
  XOR2_X1 U567 ( .A(KEYINPUT94), .B(KEYINPUT12), .Z(n474) );
  NAND2_X1 U568 ( .A1(G214), .A2(n472), .ZN(n473) );
  XNOR2_X1 U569 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U570 ( .A(n476), .B(n475), .ZN(n482) );
  XNOR2_X1 U571 ( .A(G131), .B(n477), .ZN(n479) );
  XNOR2_X1 U572 ( .A(n482), .B(n481), .ZN(n631) );
  NOR2_X1 U573 ( .A1(G902), .A2(n631), .ZN(n486) );
  XNOR2_X1 U574 ( .A(KEYINPUT96), .B(KEYINPUT13), .ZN(n484) );
  INV_X1 U575 ( .A(G475), .ZN(n483) );
  XOR2_X1 U576 ( .A(KEYINPUT9), .B(KEYINPUT97), .Z(n488) );
  XNOR2_X1 U577 ( .A(G134), .B(KEYINPUT98), .ZN(n487) );
  XNOR2_X1 U578 ( .A(n488), .B(n487), .ZN(n489) );
  XOR2_X1 U579 ( .A(n490), .B(n489), .Z(n493) );
  NAND2_X1 U580 ( .A1(G217), .A2(n491), .ZN(n492) );
  XNOR2_X1 U581 ( .A(n493), .B(n492), .ZN(n496) );
  XNOR2_X1 U582 ( .A(n494), .B(KEYINPUT7), .ZN(n495) );
  XNOR2_X1 U583 ( .A(n496), .B(n495), .ZN(n719) );
  NAND2_X1 U584 ( .A1(n719), .A2(n497), .ZN(n500) );
  XOR2_X1 U585 ( .A(G478), .B(KEYINPUT100), .Z(n498) );
  XOR2_X1 U586 ( .A(KEYINPUT99), .B(n498), .Z(n499) );
  XNOR2_X1 U587 ( .A(n500), .B(n499), .ZN(n524) );
  INV_X1 U588 ( .A(n524), .ZN(n513) );
  OR2_X1 U589 ( .A1(n525), .A2(n513), .ZN(n657) );
  NOR2_X1 U590 ( .A1(n553), .A2(n657), .ZN(n501) );
  XNOR2_X1 U591 ( .A(n501), .B(KEYINPUT40), .ZN(n759) );
  XNOR2_X1 U592 ( .A(KEYINPUT28), .B(KEYINPUT104), .ZN(n505) );
  XNOR2_X1 U593 ( .A(n506), .B(n505), .ZN(n507) );
  NAND2_X1 U594 ( .A1(n542), .A2(n507), .ZN(n508) );
  NAND2_X1 U595 ( .A1(n525), .A2(n524), .ZN(n693) );
  NAND2_X1 U596 ( .A1(n690), .A2(n689), .ZN(n695) );
  XOR2_X1 U597 ( .A(KEYINPUT41), .B(n509), .Z(n688) );
  NAND2_X1 U598 ( .A1(n520), .A2(n688), .ZN(n512) );
  XNOR2_X1 U599 ( .A(KEYINPUT106), .B(KEYINPUT42), .ZN(n510) );
  XNOR2_X1 U600 ( .A(n510), .B(KEYINPUT107), .ZN(n511) );
  NAND2_X1 U601 ( .A1(n525), .A2(n513), .ZN(n660) );
  INV_X1 U602 ( .A(n530), .ZN(n696) );
  NAND2_X1 U603 ( .A1(KEYINPUT47), .A2(n696), .ZN(n515) );
  NAND2_X1 U604 ( .A1(n515), .A2(KEYINPUT79), .ZN(n529) );
  NAND2_X1 U605 ( .A1(n516), .A2(n689), .ZN(n518) );
  INV_X1 U606 ( .A(KEYINPUT19), .ZN(n517) );
  XNOR2_X1 U607 ( .A(n518), .B(n517), .ZN(n563) );
  INV_X1 U608 ( .A(n563), .ZN(n519) );
  NAND2_X1 U609 ( .A1(n520), .A2(n519), .ZN(n655) );
  XNOR2_X1 U610 ( .A(KEYINPUT47), .B(KEYINPUT69), .ZN(n521) );
  XNOR2_X1 U611 ( .A(KEYINPUT80), .B(n530), .ZN(n591) );
  NAND2_X1 U612 ( .A1(n521), .A2(n591), .ZN(n522) );
  NOR2_X1 U613 ( .A1(n655), .A2(n522), .ZN(n527) );
  NOR2_X1 U614 ( .A1(n525), .A2(n524), .ZN(n566) );
  NAND2_X1 U615 ( .A1(n523), .A2(n566), .ZN(n526) );
  NOR2_X1 U616 ( .A1(n549), .A2(n526), .ZN(n653) );
  NOR2_X1 U617 ( .A1(n527), .A2(n653), .ZN(n528) );
  NAND2_X1 U618 ( .A1(n529), .A2(n528), .ZN(n535) );
  INV_X1 U619 ( .A(KEYINPUT47), .ZN(n533) );
  NOR2_X1 U620 ( .A1(KEYINPUT79), .A2(n530), .ZN(n531) );
  NOR2_X1 U621 ( .A1(n655), .A2(n531), .ZN(n532) );
  NOR2_X1 U622 ( .A1(n533), .A2(n532), .ZN(n534) );
  NOR2_X1 U623 ( .A1(n535), .A2(n534), .ZN(n536) );
  INV_X1 U624 ( .A(KEYINPUT6), .ZN(n538) );
  NAND2_X1 U625 ( .A1(n539), .A2(n393), .ZN(n546) );
  XNOR2_X1 U626 ( .A(n540), .B(KEYINPUT36), .ZN(n543) );
  INV_X1 U627 ( .A(KEYINPUT1), .ZN(n541) );
  XNOR2_X1 U628 ( .A(n542), .B(n541), .ZN(n555) );
  INV_X1 U629 ( .A(n674), .ZN(n593) );
  NAND2_X1 U630 ( .A1(n543), .A2(n593), .ZN(n544) );
  XNOR2_X1 U631 ( .A(n545), .B(KEYINPUT48), .ZN(n551) );
  XOR2_X1 U632 ( .A(n546), .B(KEYINPUT102), .Z(n547) );
  NAND2_X1 U633 ( .A1(n547), .A2(n674), .ZN(n548) );
  XNOR2_X1 U634 ( .A(KEYINPUT43), .B(n548), .ZN(n550) );
  NAND2_X1 U635 ( .A1(n550), .A2(n549), .ZN(n640) );
  OR2_X1 U636 ( .A1(n553), .A2(n552), .ZN(n662) );
  INV_X1 U637 ( .A(n554), .ZN(n673) );
  NOR2_X1 U638 ( .A1(n555), .A2(n673), .ZN(n585) );
  NAND2_X1 U639 ( .A1(n585), .A2(n574), .ZN(n557) );
  XOR2_X1 U640 ( .A(KEYINPUT84), .B(KEYINPUT33), .Z(n556) );
  XNOR2_X1 U641 ( .A(n557), .B(n556), .ZN(n663) );
  NOR2_X1 U642 ( .A1(G898), .A2(n747), .ZN(n558) );
  XOR2_X1 U643 ( .A(KEYINPUT88), .B(n558), .Z(n736) );
  NOR2_X1 U644 ( .A1(n736), .A2(n559), .ZN(n560) );
  NOR2_X1 U645 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U646 ( .A(n565), .B(KEYINPUT34), .ZN(n567) );
  NAND2_X1 U647 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X2 U648 ( .A(n568), .B(KEYINPUT35), .ZN(n755) );
  NOR2_X1 U649 ( .A1(n755), .A2(KEYINPUT44), .ZN(n570) );
  INV_X1 U650 ( .A(KEYINPUT64), .ZN(n569) );
  NOR2_X1 U651 ( .A1(n570), .A2(n569), .ZN(n584) );
  NOR2_X1 U652 ( .A1(n693), .A2(n676), .ZN(n571) );
  NAND2_X1 U653 ( .A1(n590), .A2(n571), .ZN(n573) );
  INV_X1 U654 ( .A(KEYINPUT22), .ZN(n572) );
  XNOR2_X1 U655 ( .A(n573), .B(n572), .ZN(n581) );
  INV_X1 U656 ( .A(n574), .ZN(n575) );
  NOR2_X1 U657 ( .A1(n674), .A2(n576), .ZN(n577) );
  INV_X1 U658 ( .A(n502), .ZN(n578) );
  INV_X1 U659 ( .A(n576), .ZN(n677) );
  AND2_X1 U660 ( .A1(n578), .A2(n677), .ZN(n579) );
  AND2_X1 U661 ( .A1(n674), .A2(n579), .ZN(n580) );
  AND2_X1 U662 ( .A1(n581), .A2(n580), .ZN(n638) );
  INV_X1 U663 ( .A(n638), .ZN(n582) );
  NAND2_X1 U664 ( .A1(n583), .A2(n582), .ZN(n599) );
  NOR2_X1 U665 ( .A1(n584), .A2(n599), .ZN(n598) );
  AND2_X1 U666 ( .A1(n502), .A2(n585), .ZN(n586) );
  XNOR2_X1 U667 ( .A(KEYINPUT93), .B(n586), .ZN(n684) );
  XNOR2_X1 U668 ( .A(n587), .B(KEYINPUT31), .ZN(n659) );
  NOR2_X1 U669 ( .A1(n588), .A2(n502), .ZN(n589) );
  NAND2_X1 U670 ( .A1(n590), .A2(n589), .ZN(n645) );
  NAND2_X1 U671 ( .A1(n659), .A2(n645), .ZN(n592) );
  NAND2_X1 U672 ( .A1(n592), .A2(n591), .ZN(n596) );
  NOR2_X1 U673 ( .A1(n593), .A2(n677), .ZN(n594) );
  NAND2_X1 U674 ( .A1(n595), .A2(n594), .ZN(n641) );
  NAND2_X1 U675 ( .A1(n596), .A2(n641), .ZN(n597) );
  NAND2_X1 U676 ( .A1(n599), .A2(KEYINPUT64), .ZN(n601) );
  INV_X1 U677 ( .A(KEYINPUT44), .ZN(n602) );
  NOR2_X1 U678 ( .A1(n755), .A2(n602), .ZN(n600) );
  NAND2_X1 U679 ( .A1(n601), .A2(n600), .ZN(n604) );
  NAND2_X1 U680 ( .A1(n602), .A2(KEYINPUT64), .ZN(n603) );
  NAND2_X1 U681 ( .A1(n604), .A2(n603), .ZN(n605) );
  NAND2_X1 U682 ( .A1(n606), .A2(n605), .ZN(n608) );
  XNOR2_X1 U683 ( .A(KEYINPUT82), .B(KEYINPUT45), .ZN(n607) );
  XNOR2_X2 U684 ( .A(n608), .B(n607), .ZN(n727) );
  AND2_X2 U685 ( .A1(n745), .A2(n727), .ZN(n665) );
  INV_X1 U686 ( .A(KEYINPUT2), .ZN(n609) );
  NOR2_X1 U687 ( .A1(n609), .A2(KEYINPUT67), .ZN(n610) );
  INV_X1 U688 ( .A(n611), .ZN(n612) );
  NAND2_X1 U689 ( .A1(n612), .A2(KEYINPUT2), .ZN(n613) );
  INV_X1 U690 ( .A(n727), .ZN(n617) );
  NAND2_X1 U691 ( .A1(KEYINPUT2), .A2(n662), .ZN(n614) );
  XNOR2_X1 U692 ( .A(n614), .B(KEYINPUT77), .ZN(n615) );
  NOR2_X1 U693 ( .A1(n617), .A2(n616), .ZN(n668) );
  NAND2_X1 U694 ( .A1(n711), .A2(G210), .ZN(n621) );
  XOR2_X1 U695 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n619) );
  XOR2_X1 U696 ( .A(n619), .B(n618), .Z(n620) );
  XNOR2_X1 U697 ( .A(n621), .B(n620), .ZN(n623) );
  INV_X1 U698 ( .A(G952), .ZN(n622) );
  AND2_X1 U699 ( .A1(n622), .A2(G953), .ZN(n726) );
  XNOR2_X1 U700 ( .A(n624), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U701 ( .A1(n711), .A2(G472), .ZN(n627) );
  XOR2_X1 U702 ( .A(KEYINPUT109), .B(KEYINPUT62), .Z(n625) );
  XNOR2_X1 U703 ( .A(n627), .B(n394), .ZN(n629) );
  NAND2_X1 U704 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U705 ( .A(n630), .B(KEYINPUT63), .ZN(G57) );
  XOR2_X1 U706 ( .A(KEYINPUT59), .B(KEYINPUT123), .Z(n633) );
  XNOR2_X1 U707 ( .A(n631), .B(KEYINPUT66), .ZN(n632) );
  XNOR2_X1 U708 ( .A(n636), .B(KEYINPUT60), .ZN(G60) );
  XOR2_X1 U709 ( .A(G110), .B(KEYINPUT110), .Z(n637) );
  XNOR2_X1 U710 ( .A(n638), .B(n637), .ZN(G12) );
  XNOR2_X1 U711 ( .A(G140), .B(KEYINPUT114), .ZN(n639) );
  XNOR2_X1 U712 ( .A(n640), .B(n639), .ZN(G42) );
  XNOR2_X1 U713 ( .A(n641), .B(G101), .ZN(G3) );
  XNOR2_X1 U714 ( .A(G119), .B(KEYINPUT127), .ZN(n642) );
  XNOR2_X1 U715 ( .A(n643), .B(n642), .ZN(G21) );
  NOR2_X1 U716 ( .A1(n657), .A2(n645), .ZN(n644) );
  XOR2_X1 U717 ( .A(G104), .B(n644), .Z(G6) );
  NOR2_X1 U718 ( .A1(n660), .A2(n645), .ZN(n647) );
  XNOR2_X1 U719 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n646) );
  XNOR2_X1 U720 ( .A(n647), .B(n646), .ZN(n648) );
  XNOR2_X1 U721 ( .A(G107), .B(n648), .ZN(G9) );
  NOR2_X1 U722 ( .A1(n655), .A2(n660), .ZN(n652) );
  XOR2_X1 U723 ( .A(KEYINPUT111), .B(KEYINPUT29), .Z(n650) );
  XNOR2_X1 U724 ( .A(G128), .B(KEYINPUT112), .ZN(n649) );
  XNOR2_X1 U725 ( .A(n650), .B(n649), .ZN(n651) );
  XNOR2_X1 U726 ( .A(n652), .B(n651), .ZN(G30) );
  XNOR2_X1 U727 ( .A(n653), .B(G143), .ZN(n654) );
  XNOR2_X1 U728 ( .A(n654), .B(KEYINPUT113), .ZN(G45) );
  NOR2_X1 U729 ( .A1(n655), .A2(n657), .ZN(n656) );
  XOR2_X1 U730 ( .A(G146), .B(n656), .Z(G48) );
  NOR2_X1 U731 ( .A1(n657), .A2(n659), .ZN(n658) );
  XOR2_X1 U732 ( .A(G113), .B(n658), .Z(G15) );
  NOR2_X1 U733 ( .A1(n660), .A2(n659), .ZN(n661) );
  XOR2_X1 U734 ( .A(G116), .B(n661), .Z(G18) );
  XNOR2_X1 U735 ( .A(G134), .B(n662), .ZN(G36) );
  INV_X1 U736 ( .A(n663), .ZN(n700) );
  AND2_X1 U737 ( .A1(n700), .A2(n688), .ZN(n664) );
  NOR2_X1 U738 ( .A1(G953), .A2(n664), .ZN(n672) );
  INV_X1 U739 ( .A(n665), .ZN(n667) );
  XOR2_X1 U740 ( .A(KEYINPUT2), .B(KEYINPUT78), .Z(n666) );
  AND2_X1 U741 ( .A1(n667), .A2(n666), .ZN(n669) );
  XNOR2_X1 U742 ( .A(n670), .B(KEYINPUT81), .ZN(n671) );
  NAND2_X1 U743 ( .A1(n672), .A2(n671), .ZN(n709) );
  NAND2_X1 U744 ( .A1(n674), .A2(n673), .ZN(n675) );
  XNOR2_X1 U745 ( .A(KEYINPUT50), .B(n675), .ZN(n682) );
  XOR2_X1 U746 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n679) );
  NAND2_X1 U747 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U748 ( .A(n679), .B(n678), .ZN(n680) );
  NOR2_X1 U749 ( .A1(n680), .A2(n502), .ZN(n681) );
  NAND2_X1 U750 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U751 ( .A1(n684), .A2(n683), .ZN(n686) );
  XOR2_X1 U752 ( .A(KEYINPUT116), .B(KEYINPUT51), .Z(n685) );
  XNOR2_X1 U753 ( .A(n686), .B(n685), .ZN(n687) );
  NAND2_X1 U754 ( .A1(n688), .A2(n687), .ZN(n703) );
  NOR2_X1 U755 ( .A1(n690), .A2(n689), .ZN(n691) );
  XOR2_X1 U756 ( .A(KEYINPUT117), .B(n691), .Z(n692) );
  NOR2_X1 U757 ( .A1(n693), .A2(n692), .ZN(n694) );
  XOR2_X1 U758 ( .A(KEYINPUT118), .B(n694), .Z(n699) );
  NOR2_X1 U759 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U760 ( .A(KEYINPUT119), .B(n697), .ZN(n698) );
  NAND2_X1 U761 ( .A1(n699), .A2(n698), .ZN(n701) );
  NAND2_X1 U762 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U763 ( .A1(n703), .A2(n702), .ZN(n705) );
  XOR2_X1 U764 ( .A(KEYINPUT52), .B(KEYINPUT120), .Z(n704) );
  XNOR2_X1 U765 ( .A(n705), .B(n704), .ZN(n707) );
  NOR2_X1 U766 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U767 ( .A(KEYINPUT53), .B(n710), .ZN(G75) );
  NAND2_X1 U768 ( .A1(n711), .A2(G469), .ZN(n717) );
  XOR2_X1 U769 ( .A(KEYINPUT122), .B(KEYINPUT121), .Z(n713) );
  XNOR2_X1 U770 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n712) );
  XNOR2_X1 U771 ( .A(n713), .B(n712), .ZN(n714) );
  XOR2_X1 U772 ( .A(n715), .B(n714), .Z(n716) );
  XNOR2_X1 U773 ( .A(n717), .B(n716), .ZN(n718) );
  NOR2_X1 U774 ( .A1(n726), .A2(n718), .ZN(G54) );
  NOR2_X1 U775 ( .A1(n726), .A2(n722), .ZN(G63) );
  NAND2_X1 U776 ( .A1(n711), .A2(G217), .ZN(n723) );
  XNOR2_X1 U777 ( .A(n724), .B(n723), .ZN(n725) );
  NOR2_X1 U778 ( .A1(n726), .A2(n725), .ZN(G66) );
  NAND2_X1 U779 ( .A1(n727), .A2(n747), .ZN(n731) );
  NAND2_X1 U780 ( .A1(G953), .A2(G224), .ZN(n728) );
  XNOR2_X1 U781 ( .A(KEYINPUT61), .B(n728), .ZN(n729) );
  NAND2_X1 U782 ( .A1(n729), .A2(G898), .ZN(n730) );
  NAND2_X1 U783 ( .A1(n731), .A2(n730), .ZN(n738) );
  XNOR2_X1 U784 ( .A(n732), .B(G110), .ZN(n733) );
  XNOR2_X1 U785 ( .A(n733), .B(KEYINPUT124), .ZN(n734) );
  XNOR2_X1 U786 ( .A(G101), .B(n734), .ZN(n735) );
  NAND2_X1 U787 ( .A1(n736), .A2(n735), .ZN(n737) );
  XOR2_X1 U788 ( .A(n738), .B(n737), .Z(G69) );
  XNOR2_X1 U789 ( .A(KEYINPUT125), .B(KEYINPUT126), .ZN(n741) );
  XNOR2_X1 U790 ( .A(n739), .B(n424), .ZN(n740) );
  XNOR2_X1 U791 ( .A(n741), .B(n740), .ZN(n744) );
  INV_X1 U792 ( .A(n742), .ZN(n743) );
  XNOR2_X1 U793 ( .A(n744), .B(n743), .ZN(n749) );
  BUF_X1 U794 ( .A(n745), .Z(n746) );
  XNOR2_X1 U795 ( .A(n749), .B(n746), .ZN(n748) );
  NAND2_X1 U796 ( .A1(n748), .A2(n747), .ZN(n754) );
  INV_X1 U797 ( .A(n749), .ZN(n750) );
  XNOR2_X1 U798 ( .A(G227), .B(n750), .ZN(n751) );
  NAND2_X1 U799 ( .A1(n751), .A2(G900), .ZN(n752) );
  NAND2_X1 U800 ( .A1(n752), .A2(G953), .ZN(n753) );
  NAND2_X1 U801 ( .A1(n754), .A2(n753), .ZN(G72) );
  XOR2_X1 U802 ( .A(G122), .B(n755), .Z(G24) );
  XOR2_X1 U803 ( .A(n756), .B(G137), .Z(G39) );
  XOR2_X1 U804 ( .A(G125), .B(n757), .Z(n758) );
  XNOR2_X1 U805 ( .A(KEYINPUT37), .B(n758), .ZN(G27) );
  XOR2_X1 U806 ( .A(n759), .B(G131), .Z(G33) );
endmodule

