//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 1 1 1 0 1 1 1 1 1 1 0 1 0 1 1 0 1 1 0 1 1 1 0 1 1 1 1 0 1 1 0 0 0 0 1 1 1 0 0 0 1 0 1 0 1 0 0 0 0 1 1 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n764, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n859, new_n860, new_n861, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n905, new_n906, new_n907, new_n908, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n930, new_n931, new_n932, new_n933, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n949, new_n950, new_n951, new_n952,
    new_n954, new_n955;
  NAND2_X1  g000(.A1(G225gat), .A2(G233gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT80), .ZN(new_n203));
  XNOR2_X1  g002(.A(G141gat), .B(G148gat), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206));
  INV_X1    g005(.A(G155gat), .ZN(new_n207));
  INV_X1    g006(.A(G162gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n206), .B1(new_n209), .B2(KEYINPUT2), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n205), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(KEYINPUT77), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n209), .A2(KEYINPUT77), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n206), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AND3_X1   g014(.A1(new_n206), .A2(KEYINPUT78), .A3(KEYINPUT2), .ZN(new_n216));
  AOI21_X1  g015(.A(KEYINPUT78), .B1(new_n206), .B2(KEYINPUT2), .ZN(new_n217));
  NOR3_X1   g016(.A1(new_n216), .A2(new_n204), .A3(new_n217), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n211), .B1(new_n215), .B2(new_n218), .ZN(new_n219));
  OR3_X1    g018(.A1(new_n219), .A2(KEYINPUT79), .A3(KEYINPUT3), .ZN(new_n220));
  OAI21_X1  g019(.A(KEYINPUT79), .B1(new_n219), .B2(KEYINPUT3), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  XOR2_X1   g021(.A(G113gat), .B(G120gat), .Z(new_n223));
  INV_X1    g022(.A(KEYINPUT1), .ZN(new_n224));
  XNOR2_X1  g023(.A(G127gat), .B(G134gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT69), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n226), .B(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n223), .A2(new_n224), .ZN(new_n229));
  INV_X1    g028(.A(G127gat), .ZN(new_n230));
  INV_X1    g029(.A(G134gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  XOR2_X1   g031(.A(KEYINPUT68), .B(G134gat), .Z(new_n233));
  OAI211_X1 g032(.A(new_n229), .B(new_n232), .C1(new_n230), .C2(new_n233), .ZN(new_n234));
  AOI22_X1  g033(.A1(new_n228), .A2(new_n234), .B1(new_n219), .B2(KEYINPUT3), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n203), .B1(new_n222), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(new_n219), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n237), .A2(new_n228), .A3(new_n234), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(KEYINPUT4), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT4), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n237), .A2(new_n228), .A3(new_n240), .A4(new_n234), .ZN(new_n241));
  AOI21_X1  g040(.A(KEYINPUT5), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n236), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT81), .ZN(new_n244));
  OR2_X1    g043(.A1(new_n241), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n241), .A2(new_n244), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n245), .A2(new_n246), .A3(new_n239), .ZN(new_n247));
  AND2_X1   g046(.A1(new_n247), .A2(new_n236), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n228), .A2(new_n234), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(new_n219), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(new_n238), .ZN(new_n251));
  AOI21_X1  g050(.A(KEYINPUT82), .B1(new_n251), .B2(new_n203), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT82), .ZN(new_n253));
  INV_X1    g052(.A(new_n203), .ZN(new_n254));
  AOI211_X1 g053(.A(new_n253), .B(new_n254), .C1(new_n250), .C2(new_n238), .ZN(new_n255));
  OAI21_X1  g054(.A(KEYINPUT5), .B1(new_n252), .B2(new_n255), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n243), .B1(new_n248), .B2(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(G1gat), .B(G29gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n258), .B(KEYINPUT0), .ZN(new_n259));
  XNOR2_X1  g058(.A(G57gat), .B(G85gat), .ZN(new_n260));
  XOR2_X1   g059(.A(new_n259), .B(new_n260), .Z(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n257), .A2(KEYINPUT6), .A3(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT6), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n264), .B1(new_n257), .B2(new_n262), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT5), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n249), .A2(new_n219), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n237), .B1(new_n228), .B2(new_n234), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n203), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(new_n253), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n251), .A2(KEYINPUT82), .A3(new_n203), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n266), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n247), .A2(new_n236), .ZN(new_n273));
  AOI22_X1  g072(.A1(new_n272), .A2(new_n273), .B1(new_n236), .B2(new_n242), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n274), .A2(new_n261), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n263), .B1(new_n265), .B2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT103), .ZN(new_n278));
  NOR2_X1   g077(.A1(G169gat), .A2(G176gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(KEYINPUT23), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT23), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n281), .B1(G169gat), .B2(G176gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(G169gat), .A2(G176gat), .ZN(new_n283));
  AND3_X1   g082(.A1(new_n280), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  OAI21_X1  g083(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(G183gat), .A2(G190gat), .ZN(new_n286));
  AND2_X1   g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  AND3_X1   g086(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n288));
  OAI211_X1 g087(.A(new_n284), .B(KEYINPUT25), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(KEYINPUT65), .ZN(new_n290));
  OR2_X1    g089(.A1(new_n287), .A2(new_n288), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT65), .ZN(new_n292));
  NAND4_X1  g091(.A1(new_n291), .A2(new_n284), .A3(new_n292), .A4(KEYINPUT25), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n280), .A2(new_n283), .A3(new_n282), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n288), .A2(KEYINPUT64), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n287), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n288), .A2(KEYINPUT64), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n294), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  OAI211_X1 g097(.A(new_n290), .B(new_n293), .C1(KEYINPUT25), .C2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n279), .A2(KEYINPUT26), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(new_n286), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n279), .A2(KEYINPUT26), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n301), .B1(new_n283), .B2(new_n302), .ZN(new_n303));
  XOR2_X1   g102(.A(KEYINPUT67), .B(KEYINPUT28), .Z(new_n304));
  XOR2_X1   g103(.A(KEYINPUT27), .B(G183gat), .Z(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(KEYINPUT66), .ZN(new_n306));
  INV_X1    g105(.A(G183gat), .ZN(new_n307));
  OR2_X1    g106(.A1(new_n307), .A2(KEYINPUT27), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT66), .ZN(new_n309));
  AOI21_X1  g108(.A(G190gat), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n304), .B1(new_n306), .B2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT28), .ZN(new_n312));
  NOR3_X1   g111(.A1(new_n305), .A2(new_n312), .A3(G190gat), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n303), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n299), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n315), .A2(new_n228), .A3(new_n234), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n299), .A2(new_n249), .A3(new_n314), .ZN(new_n317));
  AND2_X1   g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AND2_X1   g117(.A1(G227gat), .A2(G233gat), .ZN(new_n319));
  AND2_X1   g118(.A1(KEYINPUT72), .A2(KEYINPUT34), .ZN(new_n320));
  OR3_X1    g119(.A1(new_n318), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n318), .A2(new_n319), .ZN(new_n322));
  NOR2_X1   g121(.A1(KEYINPUT72), .A2(KEYINPUT34), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n320), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n321), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n316), .A2(new_n319), .A3(new_n317), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT33), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n326), .A2(KEYINPUT32), .ZN(new_n329));
  XOR2_X1   g128(.A(G15gat), .B(G43gat), .Z(new_n330));
  XNOR2_X1  g129(.A(new_n330), .B(KEYINPUT70), .ZN(new_n331));
  XNOR2_X1  g130(.A(G71gat), .B(G99gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n331), .B(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n328), .A2(new_n329), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(KEYINPUT33), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n326), .A2(KEYINPUT32), .A3(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n334), .A2(KEYINPUT71), .A3(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT71), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n328), .A2(new_n329), .A3(new_n338), .A4(new_n333), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n325), .A2(new_n337), .A3(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n325), .B1(new_n337), .B2(new_n339), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT85), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT22), .ZN(new_n346));
  XNOR2_X1  g145(.A(KEYINPUT73), .B(G218gat), .ZN(new_n347));
  INV_X1    g146(.A(G211gat), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n346), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(G197gat), .B(G204gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  XNOR2_X1  g150(.A(G211gat), .B(G218gat), .ZN(new_n352));
  XOR2_X1   g151(.A(new_n351), .B(new_n352), .Z(new_n353));
  XOR2_X1   g152(.A(KEYINPUT74), .B(KEYINPUT29), .Z(new_n354));
  AOI21_X1  g153(.A(new_n353), .B1(new_n222), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(G228gat), .A2(G233gat), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT29), .ZN(new_n358));
  INV_X1    g157(.A(new_n351), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(new_n352), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n359), .A2(new_n352), .ZN(new_n362));
  OAI211_X1 g161(.A(KEYINPUT83), .B(new_n358), .C1(new_n361), .C2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT3), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(KEYINPUT83), .B1(new_n353), .B2(new_n358), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n219), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n357), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n354), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n237), .B1(new_n369), .B2(new_n364), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n356), .B1(new_n355), .B2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(G22gat), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n368), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(G78gat), .B(G106gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(KEYINPUT31), .B(G50gat), .ZN(new_n375));
  XOR2_X1   g174(.A(new_n374), .B(new_n375), .Z(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n373), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n372), .B1(new_n368), .B2(new_n371), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n345), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n379), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n381), .A2(KEYINPUT85), .A3(new_n377), .A4(new_n373), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT84), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n373), .A2(new_n383), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n368), .A2(new_n371), .A3(KEYINPUT84), .A4(new_n372), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n384), .A2(new_n381), .A3(new_n385), .ZN(new_n386));
  AOI22_X1  g185(.A1(new_n380), .A2(new_n382), .B1(new_n386), .B2(new_n376), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n344), .A2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n353), .ZN(new_n389));
  INV_X1    g188(.A(G226gat), .ZN(new_n390));
  INV_X1    g189(.A(G233gat), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n392), .B1(new_n315), .B2(new_n354), .ZN(new_n393));
  AOI211_X1 g192(.A(new_n390), .B(new_n391), .C1(new_n299), .C2(new_n314), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n389), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n315), .A2(new_n392), .ZN(new_n396));
  AOI21_X1  g195(.A(KEYINPUT29), .B1(new_n299), .B2(new_n314), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n396), .B(new_n353), .C1(new_n392), .C2(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n395), .A2(KEYINPUT75), .A3(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT75), .ZN(new_n400));
  OAI211_X1 g199(.A(new_n400), .B(new_n389), .C1(new_n393), .C2(new_n394), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(G8gat), .B(G36gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(G64gat), .B(G92gat), .ZN(new_n404));
  XOR2_X1   g203(.A(new_n403), .B(new_n404), .Z(new_n405));
  NAND2_X1  g204(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT76), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT30), .ZN(new_n409));
  INV_X1    g208(.A(new_n405), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n410), .B1(new_n399), .B2(new_n401), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(KEYINPUT76), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n408), .A2(new_n409), .A3(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n399), .A2(new_n410), .A3(new_n401), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n415), .B1(KEYINPUT30), .B2(new_n411), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n263), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n274), .A2(KEYINPUT87), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT87), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n257), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n419), .A2(new_n421), .A3(new_n262), .ZN(new_n422));
  AOI21_X1  g221(.A(KEYINPUT6), .B1(new_n274), .B2(new_n261), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n418), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NOR3_X1   g223(.A1(new_n417), .A2(new_n424), .A3(KEYINPUT35), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n380), .A2(new_n382), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n386), .A2(new_n376), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n414), .B1(new_n406), .B2(new_n409), .ZN(new_n429));
  AOI21_X1  g228(.A(KEYINPUT76), .B1(new_n402), .B2(new_n405), .ZN(new_n430));
  AOI211_X1 g229(.A(new_n407), .B(new_n410), .C1(new_n399), .C2(new_n401), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n429), .B1(new_n432), .B2(new_n409), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n428), .A2(new_n433), .A3(new_n343), .A4(new_n276), .ZN(new_n434));
  AOI22_X1  g233(.A1(new_n388), .A2(new_n425), .B1(new_n434), .B2(KEYINPUT35), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT36), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n436), .B1(new_n341), .B2(new_n342), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n337), .A2(new_n339), .ZN(new_n438));
  INV_X1    g237(.A(new_n325), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n440), .A2(KEYINPUT36), .A3(new_n340), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n437), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n413), .A2(new_n276), .A3(new_n416), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(new_n387), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT37), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n405), .B1(new_n402), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n399), .A2(KEYINPUT37), .A3(new_n401), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(KEYINPUT38), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n397), .A2(new_n392), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n451), .A2(new_n394), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n446), .B1(new_n452), .B2(new_n389), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n353), .B1(new_n393), .B2(new_n394), .ZN(new_n454));
  AOI21_X1  g253(.A(KEYINPUT38), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n447), .A2(new_n455), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n424), .A2(new_n450), .A3(new_n432), .A4(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n222), .A2(new_n235), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n239), .A2(new_n241), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n254), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT39), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n262), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n250), .A2(new_n254), .A3(new_n238), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(KEYINPUT39), .ZN(new_n464));
  XNOR2_X1  g263(.A(new_n464), .B(KEYINPUT86), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n462), .B1(new_n465), .B2(new_n460), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n466), .B(KEYINPUT40), .ZN(new_n467));
  NOR3_X1   g266(.A1(new_n430), .A2(new_n431), .A3(KEYINPUT30), .ZN(new_n468));
  OAI211_X1 g267(.A(new_n422), .B(new_n467), .C1(new_n468), .C2(new_n429), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n457), .A2(new_n469), .A3(new_n428), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n445), .B1(KEYINPUT88), .B2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT88), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n457), .A2(new_n469), .A3(new_n472), .A4(new_n428), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n435), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  XNOR2_X1  g273(.A(G15gat), .B(G22gat), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT16), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n475), .B1(new_n476), .B2(G1gat), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n477), .B1(G1gat), .B2(new_n475), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(G8gat), .ZN(new_n479));
  INV_X1    g278(.A(G8gat), .ZN(new_n480));
  OAI211_X1 g279(.A(new_n477), .B(new_n480), .C1(G1gat), .C2(new_n475), .ZN(new_n481));
  NOR2_X1   g280(.A1(G29gat), .A2(G36gat), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT14), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT14), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n484), .B1(G29gat), .B2(G36gat), .ZN(new_n485));
  NAND2_X1  g284(.A1(G29gat), .A2(G36gat), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n483), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT15), .ZN(new_n488));
  INV_X1    g287(.A(G43gat), .ZN(new_n489));
  INV_X1    g288(.A(G50gat), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(G43gat), .A2(G50gat), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n488), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n487), .A2(new_n493), .ZN(new_n494));
  AND2_X1   g293(.A1(G29gat), .A2(G36gat), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n495), .B1(KEYINPUT14), .B2(new_n482), .ZN(new_n496));
  AND2_X1   g295(.A1(G43gat), .A2(G50gat), .ZN(new_n497));
  NOR2_X1   g296(.A1(G43gat), .A2(G50gat), .ZN(new_n498));
  OAI21_X1  g297(.A(KEYINPUT15), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n491), .A2(new_n488), .A3(new_n492), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n496), .A2(new_n499), .A3(new_n500), .A4(new_n485), .ZN(new_n501));
  AOI22_X1  g300(.A1(new_n479), .A2(new_n481), .B1(new_n494), .B2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(G229gat), .A2(G233gat), .ZN(new_n504));
  XNOR2_X1  g303(.A(new_n504), .B(KEYINPUT91), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT90), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n501), .A2(new_n494), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT17), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  AOI211_X1 g308(.A(KEYINPUT90), .B(KEYINPUT17), .C1(new_n501), .C2(new_n494), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n501), .A2(KEYINPUT17), .A3(new_n494), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n479), .A2(new_n481), .A3(new_n512), .ZN(new_n513));
  OAI211_X1 g312(.A(new_n503), .B(new_n505), .C1(new_n511), .C2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT92), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT18), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT18), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n514), .A2(new_n515), .A3(new_n518), .ZN(new_n519));
  XOR2_X1   g318(.A(new_n505), .B(KEYINPUT13), .Z(new_n520));
  NAND2_X1  g319(.A1(new_n479), .A2(new_n481), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n521), .A2(new_n507), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n520), .B1(new_n522), .B2(new_n502), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n517), .A2(new_n519), .A3(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(G113gat), .B(G141gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n525), .B(new_n526), .ZN(new_n527));
  XNOR2_X1  g326(.A(G169gat), .B(G197gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n527), .B(new_n528), .ZN(new_n529));
  XOR2_X1   g328(.A(new_n529), .B(KEYINPUT12), .Z(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n524), .A2(new_n531), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n517), .A2(new_n519), .A3(new_n523), .A4(new_n530), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n532), .A2(KEYINPUT93), .A3(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT93), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n524), .A2(new_n535), .A3(new_n531), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n474), .A2(new_n537), .ZN(new_n538));
  AND2_X1   g337(.A1(G71gat), .A2(G78gat), .ZN(new_n539));
  NOR2_X1   g338(.A1(G71gat), .A2(G78gat), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  OR2_X1    g341(.A1(new_n539), .A2(KEYINPUT9), .ZN(new_n543));
  INV_X1    g342(.A(G64gat), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT95), .ZN(new_n545));
  INV_X1    g344(.A(G57gat), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(KEYINPUT95), .A2(G57gat), .A3(G64gat), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n542), .A2(new_n543), .A3(new_n547), .A4(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n546), .A2(new_n544), .ZN(new_n550));
  NAND2_X1  g349(.A1(G57gat), .A2(G64gat), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n550), .A2(KEYINPUT9), .A3(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT94), .ZN(new_n553));
  AND3_X1   g352(.A1(new_n552), .A2(new_n553), .A3(new_n541), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n553), .B1(new_n552), .B2(new_n541), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n549), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n557), .A2(KEYINPUT21), .ZN(new_n558));
  NAND2_X1  g357(.A1(G231gat), .A2(G233gat), .ZN(new_n559));
  XOR2_X1   g358(.A(new_n558), .B(new_n559), .Z(new_n560));
  XNOR2_X1  g359(.A(new_n560), .B(G127gat), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n521), .B1(new_n557), .B2(KEYINPUT21), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n561), .B(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(KEYINPUT96), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n566), .B(G155gat), .ZN(new_n567));
  XOR2_X1   g366(.A(G183gat), .B(G211gat), .Z(new_n568));
  XNOR2_X1  g367(.A(new_n567), .B(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n564), .B(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(G232gat), .A2(G233gat), .ZN(new_n571));
  XOR2_X1   g370(.A(new_n571), .B(KEYINPUT97), .Z(new_n572));
  INV_X1    g371(.A(KEYINPUT41), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(new_n231), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(new_n208), .ZN(new_n576));
  XOR2_X1   g375(.A(G190gat), .B(G218gat), .Z(new_n577));
  NAND2_X1  g376(.A1(G99gat), .A2(G106gat), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(KEYINPUT8), .ZN(new_n579));
  NAND2_X1  g378(.A1(G85gat), .A2(G92gat), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT7), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(G85gat), .ZN(new_n583));
  INV_X1    g382(.A(G92gat), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n586));
  NAND4_X1  g385(.A1(new_n579), .A2(new_n582), .A3(new_n585), .A4(new_n586), .ZN(new_n587));
  AND2_X1   g386(.A1(G99gat), .A2(G106gat), .ZN(new_n588));
  NOR2_X1   g387(.A1(G99gat), .A2(G106gat), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  AND3_X1   g391(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n593));
  AOI21_X1  g392(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AOI22_X1  g394(.A1(KEYINPUT8), .A2(new_n578), .B1(new_n583), .B2(new_n584), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n590), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n592), .A2(new_n597), .ZN(new_n598));
  AND2_X1   g397(.A1(new_n598), .A2(new_n512), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n599), .B1(new_n509), .B2(new_n510), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n572), .A2(new_n573), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n587), .A2(new_n591), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n595), .A2(new_n590), .A3(new_n596), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n601), .B1(new_n507), .B2(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n577), .B1(new_n600), .B2(new_n605), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n576), .B1(new_n606), .B2(KEYINPUT98), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(KEYINPUT99), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n600), .A2(new_n605), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(new_n577), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT99), .ZN(new_n611));
  OAI211_X1 g410(.A(new_n611), .B(new_n576), .C1(new_n606), .C2(KEYINPUT98), .ZN(new_n612));
  AND3_X1   g411(.A1(new_n608), .A2(new_n610), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n610), .B1(new_n608), .B2(new_n612), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n570), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n557), .A2(KEYINPUT10), .A3(new_n604), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n552), .A2(new_n541), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n619), .A2(KEYINPUT94), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n552), .A2(new_n553), .A3(new_n541), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT100), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n587), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(new_n590), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n587), .A2(new_n591), .A3(new_n623), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n622), .A2(new_n549), .A3(new_n625), .A4(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n556), .A2(new_n604), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT10), .ZN(new_n630));
  AOI21_X1  g429(.A(KEYINPUT101), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT101), .ZN(new_n632));
  AOI211_X1 g431(.A(new_n632), .B(KEYINPUT10), .C1(new_n627), .C2(new_n628), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n618), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(G230gat), .A2(G233gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(KEYINPUT102), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n634), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n627), .A2(new_n628), .A3(new_n636), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(G120gat), .B(G148gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(G176gat), .B(G204gat), .ZN(new_n642));
  XOR2_X1   g441(.A(new_n641), .B(new_n642), .Z(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n640), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n638), .A2(new_n639), .A3(new_n643), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n617), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n278), .B1(new_n538), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n467), .A2(new_n422), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n428), .B1(new_n433), .B2(new_n650), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n262), .B1(new_n274), .B2(KEYINPUT87), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n257), .A2(new_n420), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n423), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND4_X1  g453(.A1(new_n654), .A2(new_n432), .A3(new_n263), .A4(new_n456), .ZN(new_n655));
  INV_X1    g454(.A(new_n450), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g456(.A(KEYINPUT88), .B1(new_n651), .B2(new_n657), .ZN(new_n658));
  AND2_X1   g457(.A1(new_n442), .A2(new_n444), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n658), .A2(new_n473), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n388), .A2(new_n425), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n434), .A2(KEYINPUT35), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n537), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n648), .ZN(new_n667));
  NOR3_X1   g466(.A1(new_n666), .A2(KEYINPUT103), .A3(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n277), .B1(new_n649), .B2(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(KEYINPUT104), .B(G1gat), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(G1324gat));
  XOR2_X1   g470(.A(KEYINPUT16), .B(G8gat), .Z(new_n672));
  OAI211_X1 g471(.A(new_n417), .B(new_n672), .C1(new_n649), .C2(new_n668), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n538), .A2(new_n278), .A3(new_n648), .ZN(new_n674));
  OAI21_X1  g473(.A(KEYINPUT103), .B1(new_n666), .B2(new_n667), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n433), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n673), .B1(new_n480), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(KEYINPUT42), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT42), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n673), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n678), .A2(new_n680), .ZN(G1325gat));
  INV_X1    g480(.A(new_n442), .ZN(new_n682));
  OAI211_X1 g481(.A(G15gat), .B(new_n682), .C1(new_n649), .C2(new_n668), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n344), .B1(new_n674), .B2(new_n675), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n683), .B1(G15gat), .B2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT105), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  OAI211_X1 g486(.A(new_n683), .B(KEYINPUT105), .C1(G15gat), .C2(new_n684), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(G1326gat));
  AOI21_X1  g488(.A(new_n428), .B1(new_n674), .B2(new_n675), .ZN(new_n690));
  XOR2_X1   g489(.A(KEYINPUT43), .B(G22gat), .Z(new_n691));
  XNOR2_X1  g490(.A(new_n690), .B(new_n691), .ZN(G1327gat));
  AOI21_X1  g491(.A(new_n616), .B1(new_n660), .B2(new_n663), .ZN(new_n693));
  INV_X1    g492(.A(G29gat), .ZN(new_n694));
  INV_X1    g493(.A(new_n570), .ZN(new_n695));
  INV_X1    g494(.A(new_n647), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n697), .A2(new_n537), .ZN(new_n698));
  NAND4_X1  g497(.A1(new_n693), .A2(new_n694), .A3(new_n277), .A4(new_n698), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(KEYINPUT45), .ZN(new_n700));
  INV_X1    g499(.A(new_n698), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n474), .A2(KEYINPUT106), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT106), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n664), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n616), .A2(KEYINPUT44), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n702), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(KEYINPUT44), .B1(new_n474), .B2(new_n616), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n701), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  AND2_X1   g507(.A1(new_n708), .A2(new_n277), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n700), .B1(new_n709), .B2(new_n694), .ZN(G1328gat));
  INV_X1    g509(.A(G36gat), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n697), .A2(new_n616), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n538), .A2(new_n711), .A3(new_n417), .A4(new_n712), .ZN(new_n713));
  XOR2_X1   g512(.A(new_n713), .B(KEYINPUT46), .Z(new_n714));
  AND2_X1   g513(.A1(new_n708), .A2(new_n417), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n714), .B1(new_n715), .B2(new_n711), .ZN(G1329gat));
  NOR3_X1   g515(.A1(new_n697), .A2(G43gat), .A3(new_n616), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n538), .A2(new_n343), .A3(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT107), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n718), .B(new_n719), .ZN(new_n720));
  AND2_X1   g519(.A1(new_n708), .A2(new_n682), .ZN(new_n721));
  OAI211_X1 g520(.A(KEYINPUT47), .B(new_n720), .C1(new_n721), .C2(new_n489), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT47), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n489), .B1(new_n708), .B2(new_n682), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n718), .B(KEYINPUT107), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n723), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n722), .A2(new_n726), .ZN(G1330gat));
  INV_X1    g526(.A(KEYINPUT109), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n428), .A2(G50gat), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n712), .B1(new_n728), .B2(new_n730), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n731), .B1(new_n728), .B2(new_n730), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n538), .A2(new_n732), .ZN(new_n733));
  AOI211_X1 g532(.A(new_n428), .B(new_n701), .C1(new_n706), .C2(new_n707), .ZN(new_n734));
  OAI211_X1 g533(.A(KEYINPUT48), .B(new_n733), .C1(new_n734), .C2(new_n490), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n708), .A2(new_n387), .ZN(new_n736));
  AOI22_X1  g535(.A1(new_n736), .A2(G50gat), .B1(new_n538), .B2(new_n732), .ZN(new_n737));
  XOR2_X1   g536(.A(KEYINPUT108), .B(KEYINPUT48), .Z(new_n738));
  OAI21_X1  g537(.A(new_n735), .B1(new_n737), .B2(new_n738), .ZN(G1331gat));
  AND2_X1   g538(.A1(new_n702), .A2(new_n704), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n617), .A2(new_n665), .A3(new_n696), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n276), .B(KEYINPUT110), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g543(.A(KEYINPUT111), .B(G57gat), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n744), .B(new_n745), .ZN(G1332gat));
  OR2_X1    g545(.A1(new_n417), .A2(KEYINPUT112), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n417), .A2(KEYINPUT112), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n742), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g550(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n752));
  AND2_X1   g551(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n751), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n754), .B1(new_n751), .B2(new_n752), .ZN(G1333gat));
  OAI21_X1  g554(.A(G71gat), .B1(new_n742), .B2(new_n442), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n344), .A2(G71gat), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n740), .A2(new_n741), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT50), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n756), .A2(KEYINPUT50), .A3(new_n758), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(G1334gat));
  NOR2_X1   g562(.A1(new_n742), .A2(new_n428), .ZN(new_n764));
  XOR2_X1   g563(.A(new_n764), .B(G78gat), .Z(G1335gat));
  NOR2_X1   g564(.A1(new_n570), .A2(new_n665), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n767), .A2(new_n696), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n769), .B1(new_n706), .B2(new_n707), .ZN(new_n770));
  AND2_X1   g569(.A1(new_n770), .A2(new_n277), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT51), .ZN(new_n772));
  NOR4_X1   g571(.A1(new_n474), .A2(new_n772), .A3(new_n616), .A4(new_n767), .ZN(new_n773));
  AOI21_X1  g572(.A(KEYINPUT51), .B1(new_n693), .B2(new_n766), .ZN(new_n774));
  OR2_X1    g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n277), .A2(new_n583), .A3(new_n647), .ZN(new_n777));
  OAI22_X1  g576(.A1(new_n771), .A2(new_n583), .B1(new_n776), .B2(new_n777), .ZN(G1336gat));
  NAND2_X1  g577(.A1(new_n770), .A2(new_n417), .ZN(new_n779));
  NOR3_X1   g578(.A1(new_n750), .A2(G92gat), .A3(new_n696), .ZN(new_n780));
  AOI22_X1  g579(.A1(new_n779), .A2(G92gat), .B1(new_n775), .B2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT52), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n584), .B1(new_n770), .B2(new_n749), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n775), .A2(new_n780), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(new_n782), .ZN(new_n785));
  OAI22_X1  g584(.A1(new_n781), .A2(new_n782), .B1(new_n783), .B2(new_n785), .ZN(G1337gat));
  INV_X1    g585(.A(KEYINPUT113), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n344), .A2(G99gat), .A3(new_n696), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n775), .A2(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(G99gat), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n791), .B1(new_n770), .B2(new_n682), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n787), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  AOI211_X1 g592(.A(new_n442), .B(new_n769), .C1(new_n706), .C2(new_n707), .ZN(new_n794));
  OAI211_X1 g593(.A(new_n789), .B(KEYINPUT113), .C1(new_n794), .C2(new_n791), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n793), .A2(new_n795), .ZN(G1338gat));
  NOR3_X1   g595(.A1(new_n428), .A2(G106gat), .A3(new_n696), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n797), .B1(new_n773), .B2(new_n774), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT114), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  OAI211_X1 g599(.A(KEYINPUT114), .B(new_n797), .C1(new_n773), .C2(new_n774), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(G106gat), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n803), .B1(new_n770), .B2(new_n387), .ZN(new_n804));
  OAI21_X1  g603(.A(KEYINPUT53), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  AOI21_X1  g604(.A(KEYINPUT53), .B1(new_n775), .B2(new_n797), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n770), .A2(new_n387), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n806), .B1(new_n807), .B2(new_n803), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n805), .A2(new_n808), .ZN(G1339gat));
  OAI211_X1 g608(.A(new_n636), .B(new_n618), .C1(new_n631), .C2(new_n633), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n638), .A2(KEYINPUT54), .A3(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT54), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n634), .A2(new_n812), .A3(new_n637), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n811), .A2(KEYINPUT55), .A3(new_n644), .A4(new_n813), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n814), .A2(new_n646), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT55), .ZN(new_n816));
  AND3_X1   g615(.A1(new_n638), .A2(KEYINPUT54), .A3(new_n810), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n813), .A2(new_n644), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n816), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n815), .A2(new_n536), .A3(new_n534), .A4(new_n819), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n522), .A2(new_n502), .A3(new_n520), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n503), .B1(new_n511), .B2(new_n513), .ZN(new_n822));
  INV_X1    g621(.A(new_n505), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n821), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(KEYINPUT115), .B1(new_n824), .B2(new_n529), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT115), .ZN(new_n826));
  INV_X1    g625(.A(new_n529), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n822), .A2(new_n823), .ZN(new_n828));
  OAI211_X1 g627(.A(new_n826), .B(new_n827), .C1(new_n828), .C2(new_n821), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n825), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n647), .A2(new_n533), .A3(new_n830), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n615), .B1(new_n820), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n819), .A2(new_n646), .A3(new_n814), .ZN(new_n833));
  INV_X1    g632(.A(new_n614), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n608), .A2(new_n610), .A3(new_n612), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n834), .A2(new_n830), .A3(new_n533), .A4(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(KEYINPUT116), .B1(new_n833), .B2(new_n836), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n533), .A2(new_n829), .A3(new_n825), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n838), .A2(new_n613), .A3(new_n614), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT116), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n815), .A2(new_n839), .A3(new_n840), .A4(new_n819), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n837), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n695), .B1(new_n832), .B2(new_n842), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n570), .A2(new_n537), .A3(new_n696), .A4(new_n616), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n743), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  AND3_X1   g644(.A1(new_n845), .A2(new_n388), .A3(new_n750), .ZN(new_n846));
  AOI21_X1  g645(.A(G113gat), .B1(new_n846), .B2(new_n665), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n749), .A2(new_n276), .A3(new_n344), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n387), .B1(new_n843), .B2(new_n844), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n665), .A2(G113gat), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n847), .B1(new_n850), .B2(new_n851), .ZN(G1340gat));
  INV_X1    g651(.A(new_n850), .ZN(new_n853));
  OAI21_X1  g652(.A(G120gat), .B1(new_n853), .B2(new_n696), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n696), .A2(G120gat), .ZN(new_n855));
  XOR2_X1   g654(.A(new_n855), .B(KEYINPUT117), .Z(new_n856));
  NAND2_X1  g655(.A1(new_n846), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n854), .A2(new_n857), .ZN(G1341gat));
  NAND3_X1  g657(.A1(new_n850), .A2(G127gat), .A3(new_n570), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n859), .B(KEYINPUT118), .ZN(new_n860));
  AOI21_X1  g659(.A(G127gat), .B1(new_n846), .B2(new_n570), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n860), .A2(new_n861), .ZN(G1342gat));
  OAI21_X1  g661(.A(G134gat), .B1(new_n853), .B2(new_n616), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n417), .A2(new_n616), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n845), .A2(new_n233), .A3(new_n388), .A4(new_n864), .ZN(new_n865));
  OR2_X1    g664(.A1(new_n865), .A2(KEYINPUT56), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(KEYINPUT56), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n863), .A2(new_n866), .A3(new_n867), .ZN(G1343gat));
  INV_X1    g667(.A(KEYINPUT121), .ZN(new_n869));
  AOI211_X1 g668(.A(new_n428), .B(new_n682), .C1(new_n845), .C2(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n870), .B1(new_n869), .B2(new_n845), .ZN(new_n871));
  NOR4_X1   g670(.A1(new_n871), .A2(G141gat), .A3(new_n537), .A4(new_n749), .ZN(new_n872));
  XNOR2_X1  g671(.A(KEYINPUT122), .B(KEYINPUT58), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NOR3_X1   g673(.A1(new_n749), .A2(new_n682), .A3(new_n276), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n843), .A2(new_n844), .ZN(new_n876));
  AOI21_X1  g675(.A(KEYINPUT57), .B1(new_n876), .B2(new_n387), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT57), .ZN(new_n878));
  AOI211_X1 g677(.A(new_n878), .B(new_n428), .C1(new_n843), .C2(new_n844), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n875), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(G141gat), .B1(new_n880), .B2(new_n537), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n874), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n880), .A2(KEYINPUT119), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT119), .ZN(new_n884));
  OAI211_X1 g683(.A(new_n884), .B(new_n875), .C1(new_n877), .C2(new_n879), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n883), .A2(new_n665), .A3(new_n885), .ZN(new_n886));
  AND3_X1   g685(.A1(new_n886), .A2(KEYINPUT120), .A3(G141gat), .ZN(new_n887));
  AOI21_X1  g686(.A(KEYINPUT120), .B1(new_n886), .B2(G141gat), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n887), .A2(new_n888), .A3(new_n872), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT58), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n882), .B1(new_n889), .B2(new_n890), .ZN(G1344gat));
  NOR3_X1   g690(.A1(new_n871), .A2(new_n696), .A3(new_n749), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT59), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n892), .A2(new_n893), .A3(G148gat), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n883), .A2(new_n885), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n893), .B1(new_n895), .B2(new_n696), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n833), .A2(new_n836), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n695), .B1(new_n832), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(new_n844), .ZN(new_n899));
  AOI21_X1  g698(.A(KEYINPUT57), .B1(new_n899), .B2(new_n387), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n900), .A2(new_n879), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n875), .A2(KEYINPUT59), .A3(new_n647), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n896), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n894), .B1(new_n903), .B2(G148gat), .ZN(G1345gat));
  NOR3_X1   g703(.A1(new_n895), .A2(new_n207), .A3(new_n695), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n871), .A2(new_n695), .A3(new_n749), .ZN(new_n906));
  OR2_X1    g705(.A1(new_n906), .A2(KEYINPUT123), .ZN(new_n907));
  AOI21_X1  g706(.A(G155gat), .B1(new_n906), .B2(KEYINPUT123), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n905), .B1(new_n907), .B2(new_n908), .ZN(G1346gat));
  OAI21_X1  g708(.A(G162gat), .B1(new_n895), .B2(new_n616), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n864), .A2(new_n208), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n910), .B1(new_n871), .B2(new_n911), .ZN(G1347gat));
  AOI21_X1  g711(.A(new_n277), .B1(new_n843), .B2(new_n844), .ZN(new_n913));
  AND3_X1   g712(.A1(new_n913), .A2(new_n388), .A3(new_n749), .ZN(new_n914));
  AOI21_X1  g713(.A(G169gat), .B1(new_n914), .B2(new_n665), .ZN(new_n915));
  AND4_X1   g714(.A1(new_n417), .A2(new_n849), .A3(new_n343), .A4(new_n743), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n665), .A2(G169gat), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n915), .B1(new_n916), .B2(new_n917), .ZN(G1348gat));
  NAND2_X1  g717(.A1(new_n916), .A2(new_n647), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n696), .A2(G176gat), .ZN(new_n920));
  AOI22_X1  g719(.A1(new_n919), .A2(G176gat), .B1(new_n914), .B2(new_n920), .ZN(new_n921));
  XOR2_X1   g720(.A(new_n921), .B(KEYINPUT124), .Z(G1349gat));
  INV_X1    g721(.A(KEYINPUT60), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n923), .A2(KEYINPUT125), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n307), .B1(new_n916), .B2(new_n570), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n695), .A2(new_n305), .ZN(new_n926));
  AOI211_X1 g725(.A(new_n924), .B(new_n925), .C1(new_n914), .C2(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n923), .A2(KEYINPUT125), .ZN(new_n928));
  XOR2_X1   g727(.A(new_n927), .B(new_n928), .Z(G1350gat));
  INV_X1    g728(.A(G190gat), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n930), .B1(new_n916), .B2(new_n615), .ZN(new_n931));
  XOR2_X1   g730(.A(new_n931), .B(KEYINPUT61), .Z(new_n932));
  NAND3_X1  g731(.A1(new_n914), .A2(new_n930), .A3(new_n615), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(G1351gat));
  NAND4_X1  g733(.A1(new_n913), .A2(new_n387), .A3(new_n442), .A4(new_n749), .ZN(new_n935));
  XNOR2_X1  g734(.A(new_n935), .B(KEYINPUT126), .ZN(new_n936));
  AOI21_X1  g735(.A(G197gat), .B1(new_n936), .B2(new_n665), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n743), .A2(new_n442), .A3(new_n417), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n901), .A2(new_n938), .ZN(new_n939));
  AND2_X1   g738(.A1(new_n665), .A2(G197gat), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n937), .B1(new_n939), .B2(new_n940), .ZN(G1352gat));
  NAND2_X1  g740(.A1(new_n939), .A2(new_n647), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(G204gat), .ZN(new_n943));
  NOR3_X1   g742(.A1(new_n935), .A2(G204gat), .A3(new_n696), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT62), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n944), .B1(KEYINPUT127), .B2(new_n945), .ZN(new_n946));
  XNOR2_X1  g745(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n947));
  OAI211_X1 g746(.A(new_n943), .B(new_n946), .C1(new_n944), .C2(new_n947), .ZN(G1353gat));
  NAND3_X1  g747(.A1(new_n936), .A2(new_n348), .A3(new_n570), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n939), .A2(new_n570), .ZN(new_n950));
  AND3_X1   g749(.A1(new_n950), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n951));
  AOI21_X1  g750(.A(KEYINPUT63), .B1(new_n950), .B2(G211gat), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n949), .B1(new_n951), .B2(new_n952), .ZN(G1354gat));
  AOI21_X1  g752(.A(G218gat), .B1(new_n936), .B2(new_n615), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n616), .A2(new_n347), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n954), .B1(new_n939), .B2(new_n955), .ZN(G1355gat));
endmodule


