//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 0 0 1 1 1 0 1 0 0 1 1 1 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 0 1 0 0 1 1 1 1 1 0 1 0 1 1 0 0 1 0 1 0 0 0 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:34 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n706,
    new_n707, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT66), .B(KEYINPUT1), .Z(new_n188));
  XNOR2_X1  g002(.A(G143), .B(G146), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n188), .A2(G128), .A3(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G125), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n192));
  INV_X1    g006(.A(G143), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n192), .A2(new_n193), .A3(G146), .ZN(new_n194));
  INV_X1    g008(.A(G146), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G143), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n193), .A2(G146), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G128), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n190), .A2(new_n191), .A3(new_n194), .A4(new_n200), .ZN(new_n201));
  AND4_X1   g015(.A1(KEYINPUT0), .A2(new_n196), .A3(new_n197), .A4(G128), .ZN(new_n202));
  NOR2_X1   g016(.A1(KEYINPUT0), .A2(G128), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT64), .ZN(new_n204));
  XNOR2_X1  g018(.A(new_n203), .B(new_n204), .ZN(new_n205));
  AOI22_X1  g019(.A1(new_n196), .A2(new_n197), .B1(KEYINPUT0), .B2(G128), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n202), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n201), .B1(new_n207), .B2(new_n191), .ZN(new_n208));
  INV_X1    g022(.A(G224), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n209), .A2(G953), .ZN(new_n210));
  XNOR2_X1  g024(.A(new_n208), .B(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G107), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G104), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(KEYINPUT3), .ZN(new_n214));
  INV_X1    g028(.A(G104), .ZN(new_n215));
  AOI21_X1  g029(.A(G101), .B1(new_n215), .B2(G107), .ZN(new_n216));
  XNOR2_X1  g030(.A(KEYINPUT83), .B(G107), .ZN(new_n217));
  OR2_X1    g031(.A1(new_n215), .A2(KEYINPUT3), .ZN(new_n218));
  OAI211_X1 g032(.A(new_n214), .B(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT85), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AND2_X1   g035(.A1(KEYINPUT83), .A2(G107), .ZN(new_n222));
  NOR2_X1   g036(.A1(KEYINPUT83), .A2(G107), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n215), .A2(KEYINPUT3), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n226), .A2(KEYINPUT85), .A3(new_n214), .A4(new_n216), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n213), .B1(new_n224), .B2(G104), .ZN(new_n228));
  AOI22_X1  g042(.A1(new_n221), .A2(new_n227), .B1(G101), .B2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G119), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G116), .ZN(new_n231));
  INV_X1    g045(.A(G116), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G119), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  XNOR2_X1  g048(.A(KEYINPUT2), .B(G113), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT5), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n234), .A2(KEYINPUT67), .ZN(new_n239));
  XNOR2_X1  g053(.A(G116), .B(G119), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT67), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n238), .B1(new_n239), .B2(new_n242), .ZN(new_n243));
  OAI21_X1  g057(.A(G113), .B1(new_n231), .B2(KEYINPUT5), .ZN(new_n244));
  OAI211_X1 g058(.A(new_n229), .B(new_n237), .C1(new_n243), .C2(new_n244), .ZN(new_n245));
  XNOR2_X1  g059(.A(G110), .B(G122), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n215), .A2(G107), .ZN(new_n247));
  OAI211_X1 g061(.A(new_n214), .B(new_n247), .C1(new_n217), .C2(new_n218), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(KEYINPUT84), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT84), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n226), .A2(new_n250), .A3(new_n214), .A4(new_n247), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n249), .A2(new_n251), .A3(G101), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n221), .A2(new_n227), .ZN(new_n253));
  AND3_X1   g067(.A1(new_n252), .A2(KEYINPUT4), .A3(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n249), .A2(new_n251), .A3(new_n255), .A4(G101), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n239), .A2(new_n242), .ZN(new_n257));
  INV_X1    g071(.A(new_n235), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n237), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n245), .B(new_n246), .C1(new_n254), .C2(new_n260), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n245), .B1(new_n254), .B2(new_n260), .ZN(new_n262));
  XOR2_X1   g076(.A(new_n246), .B(KEYINPUT89), .Z(new_n263));
  AOI22_X1  g077(.A1(new_n261), .A2(KEYINPUT6), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  AND3_X1   g078(.A1(new_n262), .A2(KEYINPUT6), .A3(new_n263), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n211), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT90), .ZN(new_n267));
  OAI21_X1  g081(.A(KEYINPUT7), .B1(new_n209), .B2(G953), .ZN(new_n268));
  AND3_X1   g082(.A1(new_n208), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n267), .B1(new_n208), .B2(new_n268), .ZN(new_n270));
  OAI22_X1  g084(.A1(new_n269), .A2(new_n270), .B1(new_n208), .B2(new_n268), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n246), .B(KEYINPUT8), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n237), .B1(new_n243), .B2(new_n244), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n272), .B1(new_n229), .B2(new_n273), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n234), .A2(new_n238), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n237), .B1(new_n275), .B2(new_n244), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n274), .B1(new_n229), .B2(new_n276), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n271), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(G902), .B1(new_n278), .B2(new_n261), .ZN(new_n279));
  OAI21_X1  g093(.A(G210), .B1(G237), .B2(G902), .ZN(new_n280));
  AND3_X1   g094(.A1(new_n266), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n280), .B1(new_n266), .B2(new_n279), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n187), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(KEYINPUT91), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n266), .A2(new_n279), .ZN(new_n285));
  INV_X1    g099(.A(new_n280), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n266), .A2(new_n279), .A3(new_n280), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT91), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n289), .A2(new_n290), .A3(new_n187), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n284), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g106(.A(G110), .B(G140), .ZN(new_n293));
  INV_X1    g107(.A(G953), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(G227), .ZN(new_n295));
  XNOR2_X1  g109(.A(new_n293), .B(new_n295), .ZN(new_n296));
  XNOR2_X1  g110(.A(KEYINPUT81), .B(KEYINPUT82), .ZN(new_n297));
  XNOR2_X1  g111(.A(new_n296), .B(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT87), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n252), .A2(KEYINPUT4), .A3(new_n253), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n301), .A2(new_n207), .A3(new_n256), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT11), .ZN(new_n303));
  INV_X1    g117(.A(G134), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n303), .B1(new_n304), .B2(G137), .ZN(new_n305));
  INV_X1    g119(.A(G137), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n306), .A2(KEYINPUT11), .A3(G134), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n304), .A2(G137), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n305), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(G131), .ZN(new_n310));
  INV_X1    g124(.A(G131), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n305), .A2(new_n307), .A3(new_n311), .A4(new_n308), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n228), .A2(G101), .ZN(new_n315));
  AOI21_X1  g129(.A(G128), .B1(new_n196), .B2(new_n197), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n193), .A2(KEYINPUT1), .A3(G146), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(KEYINPUT86), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT86), .ZN(new_n320));
  OAI211_X1 g134(.A(new_n320), .B(new_n317), .C1(new_n189), .C2(G128), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n319), .A2(new_n190), .A3(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n253), .A2(new_n315), .A3(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT10), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT69), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n194), .A2(new_n200), .ZN(new_n327));
  NOR3_X1   g141(.A1(new_n198), .A2(new_n192), .A3(new_n199), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n190), .A2(KEYINPUT69), .A3(new_n194), .A4(new_n200), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n229), .A2(KEYINPUT10), .A3(new_n329), .A4(new_n330), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n302), .A2(new_n314), .A3(new_n325), .A4(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n190), .A2(new_n194), .A3(new_n200), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n323), .B1(new_n333), .B2(new_n229), .ZN(new_n334));
  AND3_X1   g148(.A1(new_n334), .A2(KEYINPUT12), .A3(new_n313), .ZN(new_n335));
  AOI21_X1  g149(.A(KEYINPUT12), .B1(new_n334), .B2(new_n313), .ZN(new_n336));
  OAI211_X1 g150(.A(new_n300), .B(new_n332), .C1(new_n335), .C2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  AND3_X1   g152(.A1(new_n253), .A2(new_n315), .A3(new_n322), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n333), .B1(new_n253), .B2(new_n315), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n313), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT12), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n334), .A2(KEYINPUT12), .A3(new_n313), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n300), .B1(new_n345), .B2(new_n332), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n299), .B1(new_n338), .B2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n332), .ZN(new_n348));
  AND3_X1   g162(.A1(new_n329), .A2(KEYINPUT10), .A3(new_n330), .ZN(new_n349));
  AOI22_X1  g163(.A1(new_n349), .A2(new_n229), .B1(new_n323), .B2(new_n324), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n314), .B1(new_n350), .B2(new_n302), .ZN(new_n351));
  OR3_X1    g165(.A1(new_n348), .A2(new_n351), .A3(new_n299), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n347), .A2(G469), .A3(new_n352), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n298), .B(new_n332), .C1(new_n335), .C2(new_n336), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(KEYINPUT88), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT88), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n345), .A2(new_n356), .A3(new_n298), .A4(new_n332), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n299), .B1(new_n348), .B2(new_n351), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n355), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(G469), .ZN(new_n360));
  INV_X1    g174(.A(G902), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n359), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(G469), .A2(G902), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n353), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  XNOR2_X1  g178(.A(G125), .B(G140), .ZN(new_n365));
  XNOR2_X1  g179(.A(new_n365), .B(new_n195), .ZN(new_n366));
  NOR2_X1   g180(.A1(G237), .A2(G953), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n367), .A2(G143), .A3(G214), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  AOI21_X1  g183(.A(G143), .B1(new_n367), .B2(G214), .ZN(new_n370));
  OAI211_X1 g184(.A(KEYINPUT18), .B(G131), .C1(new_n369), .C2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(G237), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n372), .A2(new_n294), .A3(G214), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(new_n193), .ZN(new_n374));
  NAND2_X1  g188(.A1(KEYINPUT18), .A2(G131), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n374), .A2(new_n368), .A3(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n366), .A2(new_n371), .A3(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(G131), .B1(new_n369), .B2(new_n370), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n374), .A2(new_n311), .A3(new_n368), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n381), .A2(KEYINPUT17), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n365), .A2(KEYINPUT16), .ZN(new_n383));
  OR3_X1    g197(.A1(new_n191), .A2(KEYINPUT16), .A3(G140), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(new_n195), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n383), .A2(G146), .A3(new_n384), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n382), .A2(new_n388), .ZN(new_n389));
  OAI211_X1 g203(.A(KEYINPUT17), .B(G131), .C1(new_n369), .C2(new_n370), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n390), .B(KEYINPUT92), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n378), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  XNOR2_X1  g206(.A(G113), .B(G122), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n393), .B(new_n215), .ZN(new_n394));
  OAI21_X1  g208(.A(KEYINPUT93), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  XOR2_X1   g209(.A(new_n390), .B(KEYINPUT92), .Z(new_n396));
  OAI211_X1 g210(.A(new_n386), .B(new_n387), .C1(new_n381), .C2(KEYINPUT17), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n377), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT93), .ZN(new_n399));
  INV_X1    g213(.A(new_n394), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n398), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  AOI22_X1  g215(.A1(new_n395), .A2(new_n401), .B1(new_n394), .B2(new_n392), .ZN(new_n402));
  OAI21_X1  g216(.A(G475), .B1(new_n402), .B2(G902), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n394), .B(new_n377), .C1(new_n396), .C2(new_n397), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n387), .A2(KEYINPUT79), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n365), .B(KEYINPUT19), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(new_n195), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT79), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n383), .A2(new_n408), .A3(G146), .A4(new_n384), .ZN(new_n409));
  AND4_X1   g223(.A1(new_n405), .A2(new_n407), .A3(new_n409), .A4(new_n381), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n400), .B1(new_n410), .B2(new_n378), .ZN(new_n411));
  AND2_X1   g225(.A1(new_n404), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(G475), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(new_n361), .ZN(new_n414));
  OAI21_X1  g228(.A(KEYINPUT20), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n404), .A2(new_n411), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT20), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n416), .A2(new_n417), .A3(new_n413), .A4(new_n361), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n415), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n403), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(KEYINPUT13), .B1(new_n199), .B2(G143), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n421), .A2(new_n304), .ZN(new_n422));
  XNOR2_X1  g236(.A(G128), .B(G143), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n422), .B(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(G122), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(G116), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n232), .A2(G122), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n224), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT94), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n426), .A2(new_n427), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(new_n217), .ZN(new_n431));
  AND3_X1   g245(.A1(new_n428), .A2(new_n429), .A3(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n429), .B1(new_n428), .B2(new_n431), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n424), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT95), .ZN(new_n435));
  OR2_X1    g249(.A1(new_n428), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n427), .A2(KEYINPUT14), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(new_n426), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n427), .A2(KEYINPUT14), .ZN(new_n439));
  OAI21_X1  g253(.A(G107), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n428), .A2(new_n435), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n423), .B(new_n304), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n436), .A2(new_n440), .A3(new_n441), .A4(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n434), .A2(new_n443), .ZN(new_n444));
  XNOR2_X1  g258(.A(KEYINPUT9), .B(G234), .ZN(new_n445));
  INV_X1    g259(.A(G217), .ZN(new_n446));
  NOR3_X1   g260(.A1(new_n445), .A2(new_n446), .A3(G953), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n444), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n434), .A2(new_n443), .A3(new_n447), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(new_n361), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(KEYINPUT96), .ZN(new_n453));
  AOI21_X1  g267(.A(G902), .B1(new_n449), .B2(new_n450), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT96), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(G478), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n458), .A2(KEYINPUT15), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n459), .B1(new_n452), .B2(KEYINPUT96), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(G234), .ZN(new_n464));
  OAI211_X1 g278(.A(G902), .B(G953), .C1(new_n464), .C2(new_n372), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n465), .B(KEYINPUT97), .ZN(new_n466));
  XNOR2_X1  g280(.A(KEYINPUT21), .B(G898), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(G952), .ZN(new_n469));
  AOI211_X1 g283(.A(G953), .B(new_n469), .C1(G234), .C2(G237), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  XOR2_X1   g286(.A(new_n472), .B(KEYINPUT98), .Z(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  NOR3_X1   g288(.A1(new_n420), .A2(new_n463), .A3(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(G221), .ZN(new_n476));
  INV_X1    g290(.A(new_n445), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n476), .B1(new_n477), .B2(new_n361), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n364), .A2(new_n475), .A3(new_n479), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n292), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n306), .A2(G134), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(new_n308), .ZN(new_n483));
  AOI21_X1  g297(.A(KEYINPUT65), .B1(new_n483), .B2(G131), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT65), .ZN(new_n485));
  AOI211_X1 g299(.A(new_n485), .B(new_n311), .C1(new_n482), .C2(new_n308), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n312), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(KEYINPUT68), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT68), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n489), .B(new_n312), .C1(new_n484), .C2(new_n486), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n488), .A2(new_n329), .A3(new_n330), .A4(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n207), .A2(new_n313), .ZN(new_n492));
  INV_X1    g306(.A(new_n259), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n491), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n333), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n492), .B1(new_n496), .B2(new_n487), .ZN(new_n497));
  AND2_X1   g311(.A1(new_n497), .A2(new_n259), .ZN(new_n498));
  OAI21_X1  g312(.A(KEYINPUT28), .B1(new_n495), .B2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT28), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n494), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT74), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  XOR2_X1   g317(.A(KEYINPUT71), .B(KEYINPUT27), .Z(new_n504));
  NAND2_X1  g318(.A1(new_n367), .A2(G210), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n504), .B(new_n505), .ZN(new_n506));
  XNOR2_X1  g320(.A(KEYINPUT26), .B(G101), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n506), .B(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n494), .A2(KEYINPUT74), .A3(new_n500), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n499), .A2(new_n503), .A3(new_n508), .A4(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT29), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n491), .A2(KEYINPUT30), .A3(new_n492), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT30), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n493), .B1(new_n497), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT70), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n512), .A2(new_n514), .A3(KEYINPUT70), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n495), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  OAI211_X1 g333(.A(new_n510), .B(new_n511), .C1(new_n519), .C2(new_n508), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n491), .A2(new_n492), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n259), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n522), .A2(KEYINPUT75), .A3(new_n494), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT75), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n521), .A2(new_n524), .A3(new_n259), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n523), .A2(KEYINPUT28), .A3(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n509), .ZN(new_n527));
  AOI21_X1  g341(.A(KEYINPUT74), .B1(new_n494), .B2(new_n500), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n526), .A2(new_n529), .A3(KEYINPUT29), .A4(new_n508), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n520), .A2(new_n361), .A3(new_n530), .ZN(new_n531));
  AND3_X1   g345(.A1(new_n531), .A2(KEYINPUT76), .A3(G472), .ZN(new_n532));
  AOI21_X1  g346(.A(KEYINPUT76), .B1(new_n531), .B2(G472), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT32), .ZN(new_n534));
  AND2_X1   g348(.A1(new_n494), .A2(new_n508), .ZN(new_n535));
  XNOR2_X1  g349(.A(KEYINPUT72), .B(KEYINPUT31), .ZN(new_n536));
  AND3_X1   g350(.A1(new_n512), .A2(new_n514), .A3(KEYINPUT70), .ZN(new_n537));
  AOI21_X1  g351(.A(KEYINPUT70), .B1(new_n512), .B2(new_n514), .ZN(new_n538));
  OAI211_X1 g352(.A(new_n535), .B(new_n536), .C1(new_n537), .C2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(KEYINPUT73), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n517), .A2(new_n518), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT73), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n541), .A2(new_n542), .A3(new_n535), .A4(new_n536), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n540), .A2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n508), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n499), .A2(new_n503), .A3(new_n509), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n535), .B1(new_n537), .B2(new_n538), .ZN(new_n547));
  AOI22_X1  g361(.A1(new_n545), .A2(new_n546), .B1(new_n547), .B2(KEYINPUT31), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n544), .A2(new_n548), .ZN(new_n549));
  NOR2_X1   g363(.A1(G472), .A2(G902), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n534), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(new_n550), .ZN(new_n552));
  AOI211_X1 g366(.A(KEYINPUT32), .B(new_n552), .C1(new_n544), .C2(new_n548), .ZN(new_n553));
  OAI22_X1  g367(.A1(new_n532), .A2(new_n533), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(KEYINPUT22), .B(G137), .ZN(new_n555));
  NOR3_X1   g369(.A1(new_n476), .A2(new_n464), .A3(G953), .ZN(new_n556));
  XOR2_X1   g370(.A(new_n555), .B(new_n556), .Z(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n199), .A2(G119), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n230), .A2(G128), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  XNOR2_X1  g375(.A(KEYINPUT24), .B(G110), .ZN(new_n562));
  OR2_X1    g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AND3_X1   g377(.A1(new_n383), .A2(G146), .A3(new_n384), .ZN(new_n564));
  AOI21_X1  g378(.A(G146), .B1(new_n383), .B2(new_n384), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n563), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(KEYINPUT77), .A2(KEYINPUT23), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n559), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(new_n560), .ZN(new_n569));
  OR2_X1    g383(.A1(KEYINPUT77), .A2(KEYINPUT23), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n559), .B1(new_n570), .B2(new_n567), .ZN(new_n571));
  OAI21_X1  g385(.A(G110), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT78), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  OAI211_X1 g388(.A(KEYINPUT78), .B(G110), .C1(new_n569), .C2(new_n571), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n566), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n570), .A2(new_n567), .ZN(new_n577));
  INV_X1    g391(.A(new_n559), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(G110), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n579), .A2(new_n580), .A3(new_n560), .A4(new_n568), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n561), .A2(new_n562), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n365), .A2(new_n195), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n583), .A2(new_n405), .A3(new_n409), .A4(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n558), .B1(new_n576), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n574), .A2(new_n575), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n588), .A2(new_n563), .A3(new_n388), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n589), .A2(new_n585), .A3(new_n557), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n587), .A2(new_n361), .A3(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT25), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n587), .A2(KEYINPUT25), .A3(new_n361), .A4(new_n590), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n446), .B1(G234), .B2(new_n361), .ZN(new_n596));
  AOI21_X1  g410(.A(KEYINPUT80), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT80), .ZN(new_n598));
  INV_X1    g412(.A(new_n596), .ZN(new_n599));
  AOI211_X1 g413(.A(new_n598), .B(new_n599), .C1(new_n593), .C2(new_n594), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n587), .A2(new_n590), .ZN(new_n601));
  NOR3_X1   g415(.A1(new_n601), .A2(G902), .A3(new_n596), .ZN(new_n602));
  NOR3_X1   g416(.A1(new_n597), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n481), .A2(new_n554), .A3(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(G101), .ZN(G3));
  NAND2_X1  g419(.A1(new_n364), .A2(new_n479), .ZN(new_n606));
  OR3_X1    g420(.A1(new_n597), .A2(new_n600), .A3(new_n602), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(G472), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n609), .B1(new_n549), .B2(new_n361), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n552), .B1(new_n544), .B2(new_n548), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AND2_X1   g426(.A1(new_n608), .A2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n187), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n614), .B1(new_n287), .B2(new_n288), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT33), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n616), .B1(new_n448), .B2(KEYINPUT99), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n449), .A2(new_n450), .A3(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n617), .B1(new_n449), .B2(new_n450), .ZN(new_n620));
  OAI21_X1  g434(.A(G478), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n458), .A2(new_n361), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n622), .B1(new_n454), .B2(new_n458), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n624), .B1(new_n403), .B2(new_n419), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n615), .A2(new_n473), .A3(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n613), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g442(.A(KEYINPUT34), .B(G104), .Z(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G6));
  NOR2_X1   g444(.A1(new_n420), .A2(new_n474), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n613), .A2(new_n615), .A3(new_n631), .A4(new_n463), .ZN(new_n632));
  XOR2_X1   g446(.A(KEYINPUT35), .B(G107), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G9));
  NAND2_X1  g448(.A1(new_n589), .A2(new_n585), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(KEYINPUT100), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n635), .A2(KEYINPUT100), .ZN(new_n638));
  OAI22_X1  g452(.A1(new_n637), .A2(new_n638), .B1(KEYINPUT36), .B2(new_n558), .ZN(new_n639));
  INV_X1    g453(.A(new_n638), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n558), .A2(KEYINPUT36), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n640), .A2(new_n641), .A3(new_n636), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n596), .A2(G902), .ZN(new_n643));
  AND3_X1   g457(.A1(new_n639), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  OR3_X1    g458(.A1(new_n597), .A2(new_n600), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n549), .A2(new_n550), .ZN(new_n646));
  AOI21_X1  g460(.A(G902), .B1(new_n544), .B2(new_n548), .ZN(new_n647));
  OAI211_X1 g461(.A(new_n645), .B(new_n646), .C1(new_n609), .C2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT101), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n610), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n651), .A2(KEYINPUT101), .A3(new_n646), .A4(new_n645), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n481), .A2(new_n650), .A3(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT37), .B(G110), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G12));
  AOI21_X1  g469(.A(new_n461), .B1(new_n457), .B2(new_n459), .ZN(new_n656));
  INV_X1    g470(.A(G900), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n470), .B1(new_n466), .B2(new_n657), .ZN(new_n658));
  NOR3_X1   g472(.A1(new_n420), .A2(new_n656), .A3(new_n658), .ZN(new_n659));
  AND4_X1   g473(.A1(new_n615), .A2(new_n364), .A3(new_n479), .A4(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n554), .A2(new_n660), .A3(new_n645), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G128), .ZN(G30));
  AND3_X1   g476(.A1(new_n420), .A2(new_n463), .A3(new_n187), .ZN(new_n663));
  NOR3_X1   g477(.A1(new_n597), .A2(new_n600), .A3(new_n644), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(KEYINPUT102), .ZN(new_n666));
  AND2_X1   g480(.A1(new_n523), .A2(new_n525), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n361), .B1(new_n667), .B2(new_n508), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n519), .A2(new_n545), .ZN(new_n669));
  OAI21_X1  g483(.A(G472), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n670), .B1(new_n551), .B2(new_n553), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n289), .B(KEYINPUT38), .ZN(new_n672));
  AND3_X1   g486(.A1(new_n666), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT103), .ZN(new_n674));
  OR2_X1    g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n606), .ZN(new_n676));
  XOR2_X1   g490(.A(new_n658), .B(KEYINPUT39), .Z(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g492(.A(new_n678), .B(KEYINPUT40), .Z(new_n679));
  NAND2_X1  g493(.A1(new_n673), .A2(new_n674), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n675), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G143), .ZN(G45));
  INV_X1    g496(.A(KEYINPUT104), .ZN(new_n683));
  INV_X1    g497(.A(new_n624), .ZN(new_n684));
  INV_X1    g498(.A(new_n658), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n420), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n683), .B1(new_n283), .B2(new_n686), .ZN(new_n687));
  AOI211_X1 g501(.A(new_n658), .B(new_n624), .C1(new_n403), .C2(new_n419), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n688), .A2(new_n289), .A3(KEYINPUT104), .A4(new_n187), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n554), .A2(new_n676), .A3(new_n645), .A4(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G146), .ZN(G48));
  NOR2_X1   g506(.A1(new_n626), .A2(new_n607), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n359), .A2(new_n361), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(G469), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT105), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n695), .A2(new_n696), .A3(new_n479), .A4(new_n362), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n695), .A2(new_n479), .A3(new_n362), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(KEYINPUT105), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n554), .A2(new_n693), .A3(new_n697), .A4(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(KEYINPUT41), .B(G113), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(G15));
  AND4_X1   g516(.A1(new_n603), .A2(new_n615), .A3(new_n631), .A4(new_n463), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n554), .A2(new_n697), .A3(new_n699), .A4(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G116), .ZN(G18));
  AND3_X1   g519(.A1(new_n699), .A2(new_n615), .A3(new_n697), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n706), .A2(new_n554), .A3(new_n475), .A4(new_n645), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G119), .ZN(G21));
  NAND2_X1  g522(.A1(new_n663), .A2(new_n289), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n709), .A2(new_n474), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n526), .A2(new_n529), .ZN(new_n711));
  AOI22_X1  g525(.A1(new_n711), .A2(new_n545), .B1(KEYINPUT31), .B2(new_n547), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n552), .B1(new_n712), .B2(new_n544), .ZN(new_n713));
  NOR3_X1   g527(.A1(new_n610), .A2(new_n607), .A3(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n710), .A2(new_n714), .A3(new_n697), .A4(new_n699), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G122), .ZN(G24));
  NOR4_X1   g530(.A1(new_n610), .A2(new_n713), .A3(new_n664), .A4(new_n686), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n717), .A2(new_n615), .A3(new_n697), .A4(new_n699), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G125), .ZN(G27));
  XNOR2_X1  g533(.A(new_n611), .B(new_n534), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n531), .A2(G472), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT76), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n531), .A2(KEYINPUT76), .A3(G472), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n607), .B1(new_n720), .B2(new_n725), .ZN(new_n726));
  NOR3_X1   g540(.A1(new_n281), .A2(new_n282), .A3(new_n614), .ZN(new_n727));
  AND3_X1   g541(.A1(new_n364), .A2(new_n727), .A3(new_n479), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n726), .A2(KEYINPUT42), .A3(new_n688), .A4(new_n728), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n554), .A2(new_n603), .A3(new_n688), .A4(new_n728), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT42), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n729), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G131), .ZN(G33));
  INV_X1    g548(.A(KEYINPUT106), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n726), .A2(new_n735), .A3(new_n659), .A4(new_n728), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n554), .A2(new_n603), .A3(new_n659), .A4(new_n728), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(KEYINPUT106), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G134), .ZN(G36));
  INV_X1    g554(.A(new_n420), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(new_n684), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(KEYINPUT43), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(KEYINPUT110), .ZN(new_n744));
  OAI211_X1 g558(.A(new_n744), .B(new_n645), .C1(new_n611), .C2(new_n610), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT44), .ZN(new_n746));
  OR2_X1    g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n745), .A2(new_n746), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n747), .A2(new_n727), .A3(new_n748), .ZN(new_n749));
  AND2_X1   g563(.A1(new_n347), .A2(new_n352), .ZN(new_n750));
  OAI21_X1  g564(.A(G469), .B1(new_n750), .B2(KEYINPUT45), .ZN(new_n751));
  AOI22_X1  g565(.A1(new_n751), .A2(KEYINPUT107), .B1(KEYINPUT45), .B2(new_n750), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT107), .ZN(new_n753));
  OAI211_X1 g567(.A(new_n753), .B(G469), .C1(new_n750), .C2(KEYINPUT45), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n755), .A2(KEYINPUT46), .A3(new_n363), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(KEYINPUT108), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n755), .A2(new_n363), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT46), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT108), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n755), .A2(new_n761), .A3(KEYINPUT46), .A4(new_n363), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n757), .A2(new_n760), .A3(new_n362), .A4(new_n762), .ZN(new_n763));
  AND3_X1   g577(.A1(new_n763), .A2(new_n479), .A3(new_n677), .ZN(new_n764));
  OR2_X1    g578(.A1(new_n764), .A2(KEYINPUT109), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(KEYINPUT109), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n749), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(new_n306), .ZN(G39));
  AND2_X1   g582(.A1(KEYINPUT111), .A2(KEYINPUT47), .ZN(new_n769));
  NOR2_X1   g583(.A1(KEYINPUT111), .A2(KEYINPUT47), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n771), .B1(new_n763), .B2(new_n479), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(new_n769), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n763), .A2(new_n479), .A3(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(new_n727), .ZN(new_n776));
  NOR4_X1   g590(.A1(new_n554), .A2(new_n603), .A3(new_n686), .A4(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(KEYINPUT112), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n773), .A2(new_n775), .A3(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G140), .ZN(G42));
  NOR2_X1   g594(.A1(new_n743), .A2(new_n471), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(new_n714), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n699), .A2(new_n615), .A3(new_n697), .ZN(new_n783));
  OAI211_X1 g597(.A(G952), .B(new_n294), .C1(new_n782), .C2(new_n783), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n699), .A2(new_n697), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n727), .ZN(new_n786));
  NOR3_X1   g600(.A1(new_n786), .A2(new_n471), .A3(new_n743), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(new_n726), .ZN(new_n788));
  XOR2_X1   g602(.A(new_n788), .B(KEYINPUT48), .Z(new_n789));
  NOR4_X1   g603(.A1(new_n786), .A2(new_n607), .A3(new_n471), .A4(new_n671), .ZN(new_n790));
  AOI211_X1 g604(.A(new_n784), .B(new_n789), .C1(new_n625), .C2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT51), .ZN(new_n792));
  AND3_X1   g606(.A1(new_n763), .A2(new_n479), .A3(new_n774), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n695), .A2(new_n362), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(KEYINPUT113), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  OAI22_X1  g610(.A1(new_n793), .A2(new_n772), .B1(new_n479), .B2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(new_n782), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n798), .A2(new_n727), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(KEYINPUT116), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n797), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n420), .A2(new_n684), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n610), .A2(new_n713), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(new_n645), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  AOI22_X1  g619(.A1(new_n790), .A2(new_n802), .B1(new_n787), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n672), .A2(new_n187), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n785), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(KEYINPUT117), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT117), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n785), .A2(new_n807), .A3(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n798), .A2(new_n809), .A3(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT50), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n812), .A2(new_n813), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n806), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n792), .B1(new_n801), .B2(new_n817), .ZN(new_n818));
  AOI211_X1 g632(.A(KEYINPUT51), .B(new_n816), .C1(new_n797), .C2(new_n800), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n791), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT114), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n700), .A2(new_n704), .A3(new_n715), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n554), .A2(new_n645), .ZN(new_n823));
  INV_X1    g637(.A(new_n475), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n823), .A2(new_n783), .A3(new_n824), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n821), .B1(new_n822), .B2(new_n825), .ZN(new_n826));
  OAI211_X1 g640(.A(new_n785), .B(new_n554), .C1(new_n693), .C2(new_n703), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n707), .A2(new_n827), .A3(KEYINPUT114), .A4(new_n715), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(new_n292), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n741), .A2(new_n463), .ZN(new_n831));
  INV_X1    g645(.A(new_n625), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n474), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n830), .A2(new_n608), .A3(new_n612), .A4(new_n833), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n653), .A2(new_n604), .A3(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(new_n728), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n420), .A2(new_n463), .A3(new_n658), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n554), .A2(new_n645), .A3(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(new_n717), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n836), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(new_n840), .ZN(new_n841));
  AND4_X1   g655(.A1(new_n733), .A2(new_n739), .A3(new_n835), .A4(new_n841), .ZN(new_n842));
  AND4_X1   g656(.A1(new_n289), .A2(new_n663), .A3(new_n664), .A4(new_n685), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n843), .A2(new_n671), .A3(new_n676), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n718), .A2(new_n691), .A3(new_n661), .A4(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT52), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n845), .B(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n829), .A2(new_n842), .A3(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT53), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n848), .B(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(KEYINPUT54), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n845), .B(KEYINPUT52), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n653), .A2(new_n604), .A3(new_n834), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n853), .A2(new_n840), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n849), .B1(new_n736), .B2(new_n738), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n852), .A2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT115), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n729), .A2(new_n732), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n707), .A2(new_n827), .A3(new_n715), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n858), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n822), .A2(new_n825), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n862), .A2(KEYINPUT115), .A3(new_n733), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT54), .B1(new_n857), .B2(new_n864), .ZN(new_n865));
  AOI22_X1  g679(.A1(new_n732), .A2(new_n729), .B1(new_n736), .B2(new_n738), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n718), .A2(new_n661), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n691), .A2(new_n844), .ZN(new_n868));
  AOI21_X1  g682(.A(KEYINPUT52), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n845), .A2(new_n846), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n866), .B(new_n854), .C1(new_n869), .C2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n826), .A2(new_n828), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n849), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n865), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n851), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g689(.A(KEYINPUT118), .B1(new_n820), .B2(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(G952), .A2(G953), .ZN(new_n877));
  XNOR2_X1  g691(.A(new_n877), .B(KEYINPUT119), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n820), .A2(new_n875), .A3(KEYINPUT118), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n796), .A2(KEYINPUT49), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n796), .A2(KEYINPUT49), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n603), .A2(new_n187), .A3(new_n479), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n672), .A2(new_n742), .A3(new_n883), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n882), .A2(new_n720), .A3(new_n670), .A4(new_n884), .ZN(new_n885));
  OAI22_X1  g699(.A1(new_n879), .A2(new_n880), .B1(new_n881), .B2(new_n885), .ZN(G75));
  NOR2_X1   g700(.A1(new_n294), .A2(G952), .ZN(new_n887));
  INV_X1    g701(.A(new_n887), .ZN(new_n888));
  AOI22_X1  g702(.A1(new_n848), .A2(new_n849), .B1(new_n857), .B2(new_n864), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n889), .A2(new_n361), .ZN(new_n890));
  AOI21_X1  g704(.A(KEYINPUT56), .B1(new_n890), .B2(G210), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n264), .A2(new_n265), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(new_n211), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(KEYINPUT55), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n888), .B1(new_n891), .B2(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n895), .B1(new_n891), .B2(new_n894), .ZN(G51));
  INV_X1    g710(.A(KEYINPUT121), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n889), .A2(new_n361), .A3(new_n755), .ZN(new_n898));
  XOR2_X1   g712(.A(new_n363), .B(KEYINPUT57), .Z(new_n899));
  INV_X1    g713(.A(KEYINPUT120), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n854), .A2(new_n855), .ZN(new_n901));
  AND3_X1   g715(.A1(new_n700), .A2(new_n704), .A3(new_n715), .ZN(new_n902));
  AND4_X1   g716(.A1(KEYINPUT115), .A2(new_n733), .A3(new_n707), .A4(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(KEYINPUT115), .B1(new_n862), .B2(new_n733), .ZN(new_n904));
  OAI211_X1 g718(.A(new_n847), .B(new_n901), .C1(new_n903), .C2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT54), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n873), .A2(new_n900), .A3(new_n905), .A4(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n907), .B1(new_n906), .B2(new_n889), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n900), .B1(new_n865), .B2(new_n873), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n899), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n898), .B1(new_n910), .B2(new_n359), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n897), .B1(new_n911), .B2(new_n887), .ZN(new_n912));
  INV_X1    g726(.A(new_n359), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n874), .A2(KEYINPUT120), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n873), .A2(new_n905), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(KEYINPUT54), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n914), .A2(new_n907), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n913), .B1(new_n917), .B2(new_n899), .ZN(new_n918));
  OAI211_X1 g732(.A(KEYINPUT121), .B(new_n888), .C1(new_n918), .C2(new_n898), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n912), .A2(new_n919), .ZN(G54));
  AND3_X1   g734(.A1(new_n890), .A2(KEYINPUT58), .A3(G475), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n888), .B1(new_n921), .B2(new_n416), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n922), .B1(new_n416), .B2(new_n921), .ZN(G60));
  OR2_X1    g737(.A1(new_n619), .A2(new_n620), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n622), .B(KEYINPUT59), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n887), .B1(new_n917), .B2(new_n926), .ZN(new_n927));
  AND2_X1   g741(.A1(new_n927), .A2(KEYINPUT122), .ZN(new_n928));
  AOI22_X1  g742(.A1(new_n850), .A2(KEYINPUT54), .B1(new_n873), .B2(new_n865), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n924), .B1(new_n929), .B2(new_n925), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n930), .B1(new_n927), .B2(KEYINPUT122), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n928), .A2(new_n931), .ZN(G63));
  OR3_X1    g746(.A1(new_n446), .A2(new_n361), .A3(KEYINPUT60), .ZN(new_n933));
  OAI21_X1  g747(.A(KEYINPUT60), .B1(new_n446), .B2(new_n361), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n915), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n887), .B1(new_n935), .B2(new_n601), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n639), .A2(new_n642), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n936), .B1(new_n937), .B2(new_n935), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n938), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g753(.A(G953), .B1(new_n467), .B2(new_n209), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n872), .A2(new_n853), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n940), .B1(new_n941), .B2(G953), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n892), .B1(G898), .B2(new_n294), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT124), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(KEYINPUT123), .Z(new_n945));
  XNOR2_X1  g759(.A(new_n942), .B(new_n945), .ZN(G69));
  AND2_X1   g760(.A1(new_n867), .A2(new_n691), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n681), .A2(new_n947), .ZN(new_n948));
  OR2_X1    g762(.A1(new_n948), .A2(KEYINPUT62), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(KEYINPUT62), .ZN(new_n950));
  INV_X1    g764(.A(new_n726), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n831), .A2(new_n832), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(new_n727), .ZN(new_n953));
  NOR3_X1   g767(.A1(new_n951), .A2(new_n678), .A3(new_n953), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT126), .Z(new_n955));
  NAND4_X1  g769(.A1(new_n949), .A2(new_n779), .A3(new_n950), .A4(new_n955), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n294), .B1(new_n956), .B2(new_n767), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n497), .A2(new_n513), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n512), .A2(new_n958), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT125), .Z(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(new_n406), .ZN(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n957), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n765), .A2(new_n766), .ZN(new_n964));
  INV_X1    g778(.A(new_n749), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n951), .A2(new_n709), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n964), .A2(new_n967), .ZN(new_n968));
  AND3_X1   g782(.A1(new_n779), .A2(new_n866), .A3(new_n947), .ZN(new_n969));
  AND4_X1   g783(.A1(new_n294), .A2(new_n966), .A3(new_n968), .A4(new_n969), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n961), .B1(new_n657), .B2(new_n294), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n963), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n294), .B1(G227), .B2(G900), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(new_n973), .ZN(new_n975));
  OAI211_X1 g789(.A(new_n963), .B(new_n975), .C1(new_n970), .C2(new_n971), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n974), .A2(new_n976), .ZN(G72));
  NAND2_X1  g791(.A1(G472), .A2(G902), .ZN(new_n978));
  XOR2_X1   g792(.A(new_n978), .B(KEYINPUT63), .Z(new_n979));
  OAI21_X1  g793(.A(new_n547), .B1(new_n519), .B2(new_n508), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n850), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(new_n888), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n519), .A2(new_n545), .ZN(new_n983));
  NAND4_X1  g797(.A1(new_n966), .A2(new_n968), .A3(new_n941), .A4(new_n969), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n979), .B(KEYINPUT127), .Z(new_n985));
  AOI21_X1  g799(.A(new_n983), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n956), .A2(new_n767), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n987), .A2(new_n941), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n988), .A2(new_n985), .ZN(new_n989));
  AOI211_X1 g803(.A(new_n982), .B(new_n986), .C1(new_n669), .C2(new_n989), .ZN(G57));
endmodule


