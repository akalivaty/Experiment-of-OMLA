

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587;

  XOR2_X1 U325 ( .A(n440), .B(n439), .Z(n293) );
  XOR2_X1 U326 ( .A(n366), .B(KEYINPUT91), .Z(n294) );
  INV_X1 U327 ( .A(KEYINPUT93), .ZN(n350) );
  XNOR2_X1 U328 ( .A(n441), .B(n293), .ZN(n442) );
  XNOR2_X1 U329 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U330 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U331 ( .A(n353), .B(n352), .ZN(n355) );
  XOR2_X1 U332 ( .A(n359), .B(n358), .Z(n514) );
  XNOR2_X1 U333 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U334 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n450) );
  XNOR2_X1 U335 ( .A(G99GAT), .B(KEYINPUT102), .ZN(n448) );
  XNOR2_X1 U336 ( .A(n474), .B(n473), .ZN(G1351GAT) );
  XNOR2_X1 U337 ( .A(n449), .B(n448), .ZN(G1338GAT) );
  XNOR2_X1 U338 ( .A(G176GAT), .B(KEYINPUT18), .ZN(n295) );
  XNOR2_X1 U339 ( .A(n295), .B(KEYINPUT17), .ZN(n296) );
  XOR2_X1 U340 ( .A(n296), .B(KEYINPUT19), .Z(n298) );
  XNOR2_X1 U341 ( .A(G169GAT), .B(G190GAT), .ZN(n297) );
  XNOR2_X1 U342 ( .A(n298), .B(n297), .ZN(n357) );
  XOR2_X1 U343 ( .A(KEYINPUT79), .B(KEYINPUT20), .Z(n300) );
  XNOR2_X1 U344 ( .A(KEYINPUT80), .B(KEYINPUT78), .ZN(n299) );
  XNOR2_X1 U345 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U346 ( .A(n357), .B(n301), .ZN(n310) );
  XOR2_X1 U347 ( .A(G99GAT), .B(G71GAT), .Z(n433) );
  XNOR2_X1 U348 ( .A(G43GAT), .B(G15GAT), .ZN(n302) );
  XNOR2_X1 U349 ( .A(n302), .B(G113GAT), .ZN(n428) );
  XOR2_X1 U350 ( .A(n433), .B(n428), .Z(n304) );
  NAND2_X1 U351 ( .A1(G227GAT), .A2(G233GAT), .ZN(n303) );
  XNOR2_X1 U352 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U353 ( .A(n305), .B(G120GAT), .Z(n308) );
  XNOR2_X1 U354 ( .A(G134GAT), .B(G127GAT), .ZN(n306) );
  XNOR2_X1 U355 ( .A(n306), .B(KEYINPUT0), .ZN(n328) );
  XNOR2_X1 U356 ( .A(n328), .B(G183GAT), .ZN(n307) );
  XNOR2_X1 U357 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U358 ( .A(n310), .B(n309), .ZN(n520) );
  INV_X1 U359 ( .A(n520), .ZN(n505) );
  XOR2_X1 U360 ( .A(KEYINPUT13), .B(G78GAT), .Z(n312) );
  XNOR2_X1 U361 ( .A(G8GAT), .B(G155GAT), .ZN(n311) );
  XNOR2_X1 U362 ( .A(n312), .B(n311), .ZN(n316) );
  XOR2_X1 U363 ( .A(KEYINPUT76), .B(KEYINPUT77), .Z(n314) );
  XNOR2_X1 U364 ( .A(KEYINPUT15), .B(KEYINPUT14), .ZN(n313) );
  XNOR2_X1 U365 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U366 ( .A(n316), .B(n315), .ZN(n327) );
  XOR2_X1 U367 ( .A(G1GAT), .B(G57GAT), .Z(n329) );
  XOR2_X1 U368 ( .A(G71GAT), .B(G127GAT), .Z(n318) );
  XNOR2_X1 U369 ( .A(G15GAT), .B(G22GAT), .ZN(n317) );
  XNOR2_X1 U370 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U371 ( .A(n329), .B(n319), .Z(n321) );
  NAND2_X1 U372 ( .A1(G231GAT), .A2(G233GAT), .ZN(n320) );
  XNOR2_X1 U373 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U374 ( .A(n322), .B(KEYINPUT12), .Z(n325) );
  XNOR2_X1 U375 ( .A(G183GAT), .B(G211GAT), .ZN(n323) );
  XNOR2_X1 U376 ( .A(n323), .B(KEYINPUT75), .ZN(n354) );
  XNOR2_X1 U377 ( .A(G64GAT), .B(n354), .ZN(n324) );
  XNOR2_X1 U378 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U379 ( .A(n327), .B(n326), .ZN(n545) );
  XOR2_X1 U380 ( .A(n329), .B(n328), .Z(n331) );
  NAND2_X1 U381 ( .A1(G225GAT), .A2(G233GAT), .ZN(n330) );
  XNOR2_X1 U382 ( .A(n331), .B(n330), .ZN(n342) );
  XOR2_X1 U383 ( .A(KEYINPUT5), .B(KEYINPUT88), .Z(n333) );
  XNOR2_X1 U384 ( .A(KEYINPUT1), .B(KEYINPUT89), .ZN(n332) );
  XNOR2_X1 U385 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U386 ( .A(G120GAT), .B(G148GAT), .Z(n437) );
  XOR2_X1 U387 ( .A(n334), .B(n437), .Z(n336) );
  XNOR2_X1 U388 ( .A(G113GAT), .B(G141GAT), .ZN(n335) );
  XNOR2_X1 U389 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U390 ( .A(n337), .B(KEYINPUT4), .Z(n340) );
  XNOR2_X1 U391 ( .A(G29GAT), .B(KEYINPUT74), .ZN(n338) );
  XNOR2_X1 U392 ( .A(n338), .B(G85GAT), .ZN(n399) );
  XNOR2_X1 U393 ( .A(n399), .B(KEYINPUT6), .ZN(n339) );
  XNOR2_X1 U394 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U395 ( .A(n342), .B(n341), .ZN(n346) );
  XOR2_X1 U396 ( .A(KEYINPUT85), .B(G162GAT), .Z(n344) );
  XNOR2_X1 U397 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n343) );
  XNOR2_X1 U398 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U399 ( .A(KEYINPUT2), .B(n345), .ZN(n376) );
  XNOR2_X1 U400 ( .A(n346), .B(n376), .ZN(n387) );
  XNOR2_X1 U401 ( .A(KEYINPUT90), .B(n387), .ZN(n465) );
  INV_X1 U402 ( .A(n465), .ZN(n566) );
  XOR2_X1 U403 ( .A(KEYINPUT84), .B(KEYINPUT21), .Z(n348) );
  XNOR2_X1 U404 ( .A(G197GAT), .B(G218GAT), .ZN(n347) );
  XNOR2_X1 U405 ( .A(n348), .B(n347), .ZN(n366) );
  NAND2_X1 U406 ( .A1(G226GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U407 ( .A(n294), .B(n349), .ZN(n353) );
  XOR2_X1 U408 ( .A(G36GAT), .B(G8GAT), .Z(n416) );
  XNOR2_X1 U409 ( .A(n416), .B(KEYINPUT92), .ZN(n351) );
  XOR2_X1 U410 ( .A(n355), .B(n354), .Z(n359) );
  XNOR2_X1 U411 ( .A(G204GAT), .B(G92GAT), .ZN(n356) );
  XNOR2_X1 U412 ( .A(n356), .B(G64GAT), .ZN(n434) );
  XNOR2_X1 U413 ( .A(n357), .B(n434), .ZN(n358) );
  XNOR2_X1 U414 ( .A(n514), .B(KEYINPUT94), .ZN(n360) );
  XNOR2_X1 U415 ( .A(KEYINPUT27), .B(n360), .ZN(n383) );
  NAND2_X1 U416 ( .A1(n566), .A2(n383), .ZN(n516) );
  XNOR2_X1 U417 ( .A(KEYINPUT81), .B(n520), .ZN(n361) );
  NOR2_X1 U418 ( .A1(n516), .A2(n361), .ZN(n379) );
  XOR2_X1 U419 ( .A(G106GAT), .B(G78GAT), .Z(n438) );
  XNOR2_X1 U420 ( .A(G50GAT), .B(G22GAT), .ZN(n362) );
  XNOR2_X1 U421 ( .A(n362), .B(G141GAT), .ZN(n427) );
  XOR2_X1 U422 ( .A(n438), .B(n427), .Z(n364) );
  NAND2_X1 U423 ( .A1(G228GAT), .A2(G233GAT), .ZN(n363) );
  XNOR2_X1 U424 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U425 ( .A(n365), .B(KEYINPUT83), .Z(n368) );
  XNOR2_X1 U426 ( .A(n366), .B(KEYINPUT23), .ZN(n367) );
  XNOR2_X1 U427 ( .A(n368), .B(n367), .ZN(n372) );
  XOR2_X1 U428 ( .A(KEYINPUT22), .B(KEYINPUT82), .Z(n370) );
  XNOR2_X1 U429 ( .A(G211GAT), .B(KEYINPUT87), .ZN(n369) );
  XNOR2_X1 U430 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U431 ( .A(n372), .B(n371), .Z(n378) );
  XOR2_X1 U432 ( .A(G148GAT), .B(G204GAT), .Z(n374) );
  XNOR2_X1 U433 ( .A(KEYINPUT24), .B(KEYINPUT86), .ZN(n373) );
  XNOR2_X1 U434 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U435 ( .A(n376), .B(n375), .Z(n377) );
  XNOR2_X1 U436 ( .A(n378), .B(n377), .ZN(n467) );
  XOR2_X1 U437 ( .A(n467), .B(KEYINPUT28), .Z(n518) );
  NAND2_X1 U438 ( .A1(n379), .A2(n518), .ZN(n389) );
  AND2_X1 U439 ( .A1(n505), .A2(n514), .ZN(n380) );
  NOR2_X1 U440 ( .A1(n467), .A2(n380), .ZN(n381) );
  XNOR2_X1 U441 ( .A(n381), .B(KEYINPUT25), .ZN(n385) );
  NAND2_X1 U442 ( .A1(n467), .A2(n520), .ZN(n382) );
  XOR2_X1 U443 ( .A(n382), .B(KEYINPUT26), .Z(n564) );
  NAND2_X1 U444 ( .A1(n383), .A2(n564), .ZN(n384) );
  NAND2_X1 U445 ( .A1(n385), .A2(n384), .ZN(n386) );
  NAND2_X1 U446 ( .A1(n387), .A2(n386), .ZN(n388) );
  NAND2_X1 U447 ( .A1(n389), .A2(n388), .ZN(n390) );
  XNOR2_X1 U448 ( .A(n390), .B(KEYINPUT95), .ZN(n476) );
  XOR2_X1 U449 ( .A(KEYINPUT64), .B(KEYINPUT9), .Z(n392) );
  XNOR2_X1 U450 ( .A(KEYINPUT73), .B(KEYINPUT11), .ZN(n391) );
  XNOR2_X1 U451 ( .A(n392), .B(n391), .ZN(n410) );
  XOR2_X1 U452 ( .A(G106GAT), .B(G162GAT), .Z(n394) );
  XNOR2_X1 U453 ( .A(G134GAT), .B(G99GAT), .ZN(n393) );
  XNOR2_X1 U454 ( .A(n394), .B(n393), .ZN(n398) );
  XOR2_X1 U455 ( .A(G92GAT), .B(G36GAT), .Z(n396) );
  XNOR2_X1 U456 ( .A(G43GAT), .B(G50GAT), .ZN(n395) );
  XNOR2_X1 U457 ( .A(n396), .B(n395), .ZN(n397) );
  XOR2_X1 U458 ( .A(n398), .B(n397), .Z(n404) );
  XOR2_X1 U459 ( .A(KEYINPUT10), .B(n399), .Z(n401) );
  NAND2_X1 U460 ( .A1(G232GAT), .A2(G233GAT), .ZN(n400) );
  XNOR2_X1 U461 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U462 ( .A(G218GAT), .B(n402), .ZN(n403) );
  XNOR2_X1 U463 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U464 ( .A(n405), .B(KEYINPUT72), .Z(n408) );
  XNOR2_X1 U465 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n406) );
  XNOR2_X1 U466 ( .A(n406), .B(KEYINPUT68), .ZN(n420) );
  XNOR2_X1 U467 ( .A(n420), .B(G190GAT), .ZN(n407) );
  XNOR2_X1 U468 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U469 ( .A(n410), .B(n409), .ZN(n470) );
  XNOR2_X1 U470 ( .A(KEYINPUT36), .B(n470), .ZN(n582) );
  NOR2_X1 U471 ( .A1(n476), .A2(n582), .ZN(n411) );
  NAND2_X1 U472 ( .A1(n545), .A2(n411), .ZN(n412) );
  XOR2_X1 U473 ( .A(KEYINPUT37), .B(n412), .Z(n488) );
  XOR2_X1 U474 ( .A(G1GAT), .B(G197GAT), .Z(n414) );
  XNOR2_X1 U475 ( .A(G169GAT), .B(G29GAT), .ZN(n413) );
  XNOR2_X1 U476 ( .A(n414), .B(n413), .ZN(n415) );
  XOR2_X1 U477 ( .A(n416), .B(n415), .Z(n418) );
  NAND2_X1 U478 ( .A1(G229GAT), .A2(G233GAT), .ZN(n417) );
  XNOR2_X1 U479 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U480 ( .A(n419), .B(KEYINPUT65), .Z(n422) );
  XNOR2_X1 U481 ( .A(n420), .B(KEYINPUT69), .ZN(n421) );
  XNOR2_X1 U482 ( .A(n422), .B(n421), .ZN(n426) );
  XOR2_X1 U483 ( .A(KEYINPUT29), .B(KEYINPUT67), .Z(n424) );
  XNOR2_X1 U484 ( .A(KEYINPUT66), .B(KEYINPUT30), .ZN(n423) );
  XNOR2_X1 U485 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U486 ( .A(n426), .B(n425), .Z(n430) );
  XNOR2_X1 U487 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U488 ( .A(n430), .B(n429), .ZN(n569) );
  INV_X1 U489 ( .A(n569), .ZN(n446) );
  XOR2_X1 U490 ( .A(KEYINPUT13), .B(G57GAT), .Z(n432) );
  XNOR2_X1 U491 ( .A(G176GAT), .B(G85GAT), .ZN(n431) );
  XNOR2_X1 U492 ( .A(n432), .B(n431), .ZN(n445) );
  XNOR2_X1 U493 ( .A(n434), .B(n433), .ZN(n436) );
  AND2_X1 U494 ( .A1(G230GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U495 ( .A(n436), .B(n435), .ZN(n443) );
  XNOR2_X1 U496 ( .A(n438), .B(n437), .ZN(n441) );
  XOR2_X1 U497 ( .A(KEYINPUT32), .B(KEYINPUT31), .Z(n440) );
  XNOR2_X1 U498 ( .A(KEYINPUT71), .B(KEYINPUT33), .ZN(n439) );
  XOR2_X1 U499 ( .A(n445), .B(n444), .Z(n574) );
  XNOR2_X1 U500 ( .A(n574), .B(KEYINPUT41), .ZN(n554) );
  NAND2_X1 U501 ( .A1(n446), .A2(n554), .ZN(n500) );
  NOR2_X1 U502 ( .A1(n488), .A2(n500), .ZN(n447) );
  XOR2_X1 U503 ( .A(KEYINPUT101), .B(n447), .Z(n513) );
  NAND2_X1 U504 ( .A1(n505), .A2(n513), .ZN(n449) );
  INV_X1 U505 ( .A(n518), .ZN(n508) );
  NAND2_X1 U506 ( .A1(n508), .A2(n513), .ZN(n451) );
  XNOR2_X1 U507 ( .A(n451), .B(n450), .ZN(G1339GAT) );
  XNOR2_X1 U508 ( .A(n545), .B(KEYINPUT103), .ZN(n560) );
  NAND2_X1 U509 ( .A1(n569), .A2(n554), .ZN(n452) );
  XOR2_X1 U510 ( .A(KEYINPUT46), .B(n452), .Z(n453) );
  NOR2_X1 U511 ( .A1(n560), .A2(n453), .ZN(n454) );
  XNOR2_X1 U512 ( .A(n454), .B(KEYINPUT104), .ZN(n455) );
  NAND2_X1 U513 ( .A1(n455), .A2(n470), .ZN(n456) );
  XNOR2_X1 U514 ( .A(n456), .B(KEYINPUT47), .ZN(n461) );
  XNOR2_X1 U515 ( .A(n569), .B(KEYINPUT70), .ZN(n552) );
  NOR2_X1 U516 ( .A1(n582), .A2(n545), .ZN(n457) );
  XNOR2_X1 U517 ( .A(KEYINPUT45), .B(n457), .ZN(n458) );
  NAND2_X1 U518 ( .A1(n458), .A2(n574), .ZN(n459) );
  NOR2_X1 U519 ( .A1(n552), .A2(n459), .ZN(n460) );
  NOR2_X1 U520 ( .A1(n461), .A2(n460), .ZN(n462) );
  XNOR2_X1 U521 ( .A(KEYINPUT48), .B(n462), .ZN(n517) );
  XOR2_X1 U522 ( .A(n514), .B(KEYINPUT118), .Z(n463) );
  NOR2_X1 U523 ( .A1(n517), .A2(n463), .ZN(n464) );
  XNOR2_X1 U524 ( .A(n464), .B(KEYINPUT54), .ZN(n568) );
  NAND2_X1 U525 ( .A1(n568), .A2(n465), .ZN(n466) );
  NOR2_X1 U526 ( .A1(n467), .A2(n466), .ZN(n468) );
  XNOR2_X1 U527 ( .A(n468), .B(KEYINPUT55), .ZN(n469) );
  NOR2_X2 U528 ( .A1(n520), .A2(n469), .ZN(n559) );
  INV_X1 U529 ( .A(n470), .ZN(n548) );
  NAND2_X1 U530 ( .A1(n559), .A2(n548), .ZN(n474) );
  XOR2_X1 U531 ( .A(KEYINPUT58), .B(KEYINPUT120), .Z(n472) );
  INV_X1 U532 ( .A(G190GAT), .ZN(n471) );
  NAND2_X1 U533 ( .A1(n574), .A2(n552), .ZN(n487) );
  NOR2_X1 U534 ( .A1(n548), .A2(n545), .ZN(n475) );
  XNOR2_X1 U535 ( .A(n475), .B(KEYINPUT16), .ZN(n478) );
  INV_X1 U536 ( .A(n476), .ZN(n477) );
  NAND2_X1 U537 ( .A1(n478), .A2(n477), .ZN(n499) );
  NOR2_X1 U538 ( .A1(n487), .A2(n499), .ZN(n485) );
  NAND2_X1 U539 ( .A1(n566), .A2(n485), .ZN(n481) );
  XNOR2_X1 U540 ( .A(G1GAT), .B(KEYINPUT96), .ZN(n479) );
  XNOR2_X1 U541 ( .A(n479), .B(KEYINPUT34), .ZN(n480) );
  XNOR2_X1 U542 ( .A(n481), .B(n480), .ZN(G1324GAT) );
  NAND2_X1 U543 ( .A1(n514), .A2(n485), .ZN(n482) );
  XNOR2_X1 U544 ( .A(n482), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U545 ( .A(G15GAT), .B(KEYINPUT35), .Z(n484) );
  NAND2_X1 U546 ( .A1(n485), .A2(n505), .ZN(n483) );
  XNOR2_X1 U547 ( .A(n484), .B(n483), .ZN(G1326GAT) );
  NAND2_X1 U548 ( .A1(n508), .A2(n485), .ZN(n486) );
  XNOR2_X1 U549 ( .A(n486), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U550 ( .A(KEYINPUT39), .B(KEYINPUT97), .Z(n491) );
  NOR2_X1 U551 ( .A1(n488), .A2(n487), .ZN(n489) );
  XNOR2_X1 U552 ( .A(n489), .B(KEYINPUT38), .ZN(n496) );
  NAND2_X1 U553 ( .A1(n496), .A2(n566), .ZN(n490) );
  XNOR2_X1 U554 ( .A(n491), .B(n490), .ZN(n492) );
  XOR2_X1 U555 ( .A(G29GAT), .B(n492), .Z(G1328GAT) );
  NAND2_X1 U556 ( .A1(n496), .A2(n514), .ZN(n493) );
  XNOR2_X1 U557 ( .A(n493), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U558 ( .A1(n505), .A2(n496), .ZN(n494) );
  XNOR2_X1 U559 ( .A(KEYINPUT40), .B(n494), .ZN(n495) );
  XNOR2_X1 U560 ( .A(G43GAT), .B(n495), .ZN(G1330GAT) );
  XNOR2_X1 U561 ( .A(G50GAT), .B(KEYINPUT98), .ZN(n498) );
  NAND2_X1 U562 ( .A1(n508), .A2(n496), .ZN(n497) );
  XNOR2_X1 U563 ( .A(n498), .B(n497), .ZN(G1331GAT) );
  XOR2_X1 U564 ( .A(KEYINPUT99), .B(KEYINPUT42), .Z(n502) );
  NOR2_X1 U565 ( .A1(n500), .A2(n499), .ZN(n509) );
  NAND2_X1 U566 ( .A1(n509), .A2(n566), .ZN(n501) );
  XNOR2_X1 U567 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U568 ( .A(G57GAT), .B(n503), .ZN(G1332GAT) );
  NAND2_X1 U569 ( .A1(n514), .A2(n509), .ZN(n504) );
  XNOR2_X1 U570 ( .A(n504), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U571 ( .A1(n505), .A2(n509), .ZN(n506) );
  XNOR2_X1 U572 ( .A(n506), .B(KEYINPUT100), .ZN(n507) );
  XNOR2_X1 U573 ( .A(G71GAT), .B(n507), .ZN(G1334GAT) );
  XOR2_X1 U574 ( .A(G78GAT), .B(KEYINPUT43), .Z(n511) );
  NAND2_X1 U575 ( .A1(n509), .A2(n508), .ZN(n510) );
  XNOR2_X1 U576 ( .A(n511), .B(n510), .ZN(G1335GAT) );
  NAND2_X1 U577 ( .A1(n513), .A2(n566), .ZN(n512) );
  XNOR2_X1 U578 ( .A(G85GAT), .B(n512), .ZN(G1336GAT) );
  NAND2_X1 U579 ( .A1(n514), .A2(n513), .ZN(n515) );
  XNOR2_X1 U580 ( .A(n515), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U581 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n522) );
  NOR2_X1 U582 ( .A1(n517), .A2(n516), .ZN(n537) );
  NAND2_X1 U583 ( .A1(n537), .A2(n518), .ZN(n519) );
  NOR2_X1 U584 ( .A1(n520), .A2(n519), .ZN(n532) );
  NAND2_X1 U585 ( .A1(n532), .A2(n552), .ZN(n521) );
  XNOR2_X1 U586 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U587 ( .A(G113GAT), .B(n523), .ZN(G1340GAT) );
  XOR2_X1 U588 ( .A(KEYINPUT107), .B(KEYINPUT49), .Z(n525) );
  NAND2_X1 U589 ( .A1(n532), .A2(n554), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n525), .B(n524), .ZN(n526) );
  XOR2_X1 U591 ( .A(G120GAT), .B(n526), .Z(G1341GAT) );
  XOR2_X1 U592 ( .A(KEYINPUT50), .B(KEYINPUT110), .Z(n528) );
  XNOR2_X1 U593 ( .A(G127GAT), .B(KEYINPUT109), .ZN(n527) );
  XNOR2_X1 U594 ( .A(n528), .B(n527), .ZN(n531) );
  NAND2_X1 U595 ( .A1(n560), .A2(n532), .ZN(n529) );
  XNOR2_X1 U596 ( .A(n529), .B(KEYINPUT108), .ZN(n530) );
  XNOR2_X1 U597 ( .A(n531), .B(n530), .ZN(G1342GAT) );
  XOR2_X1 U598 ( .A(KEYINPUT111), .B(KEYINPUT51), .Z(n534) );
  NAND2_X1 U599 ( .A1(n532), .A2(n548), .ZN(n533) );
  XNOR2_X1 U600 ( .A(n534), .B(n533), .ZN(n536) );
  XOR2_X1 U601 ( .A(G134GAT), .B(KEYINPUT112), .Z(n535) );
  XNOR2_X1 U602 ( .A(n536), .B(n535), .ZN(G1343GAT) );
  AND2_X1 U603 ( .A1(n564), .A2(n537), .ZN(n549) );
  NAND2_X1 U604 ( .A1(n569), .A2(n549), .ZN(n538) );
  XNOR2_X1 U605 ( .A(G141GAT), .B(n538), .ZN(G1344GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT115), .B(KEYINPUT114), .Z(n540) );
  XNOR2_X1 U607 ( .A(KEYINPUT113), .B(KEYINPUT53), .ZN(n539) );
  XNOR2_X1 U608 ( .A(n540), .B(n539), .ZN(n544) );
  XNOR2_X1 U609 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n542) );
  NAND2_X1 U610 ( .A1(n549), .A2(n554), .ZN(n541) );
  XNOR2_X1 U611 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U612 ( .A(n544), .B(n543), .ZN(G1345GAT) );
  INV_X1 U613 ( .A(n545), .ZN(n578) );
  NAND2_X1 U614 ( .A1(n578), .A2(n549), .ZN(n546) );
  XNOR2_X1 U615 ( .A(n546), .B(KEYINPUT116), .ZN(n547) );
  XNOR2_X1 U616 ( .A(G155GAT), .B(n547), .ZN(G1346GAT) );
  XOR2_X1 U617 ( .A(G162GAT), .B(KEYINPUT117), .Z(n551) );
  NAND2_X1 U618 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U619 ( .A(n551), .B(n550), .ZN(G1347GAT) );
  NAND2_X1 U620 ( .A1(n559), .A2(n552), .ZN(n553) );
  XNOR2_X1 U621 ( .A(G169GAT), .B(n553), .ZN(G1348GAT) );
  XOR2_X1 U622 ( .A(KEYINPUT57), .B(KEYINPUT119), .Z(n556) );
  NAND2_X1 U623 ( .A1(n559), .A2(n554), .ZN(n555) );
  XNOR2_X1 U624 ( .A(n556), .B(n555), .ZN(n558) );
  XOR2_X1 U625 ( .A(G176GAT), .B(KEYINPUT56), .Z(n557) );
  XNOR2_X1 U626 ( .A(n558), .B(n557), .ZN(G1349GAT) );
  NAND2_X1 U627 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n561), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U629 ( .A(KEYINPUT123), .B(KEYINPUT60), .Z(n563) );
  XNOR2_X1 U630 ( .A(KEYINPUT121), .B(KEYINPUT122), .ZN(n562) );
  XNOR2_X1 U631 ( .A(n563), .B(n562), .ZN(n573) );
  XOR2_X1 U632 ( .A(G197GAT), .B(KEYINPUT59), .Z(n571) );
  INV_X1 U633 ( .A(n564), .ZN(n565) );
  NOR2_X1 U634 ( .A1(n566), .A2(n565), .ZN(n567) );
  AND2_X1 U635 ( .A1(n568), .A2(n567), .ZN(n579) );
  NAND2_X1 U636 ( .A1(n579), .A2(n569), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(n572) );
  XOR2_X1 U638 ( .A(n573), .B(n572), .Z(G1352GAT) );
  XOR2_X1 U639 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n576) );
  INV_X1 U640 ( .A(n579), .ZN(n581) );
  OR2_X1 U641 ( .A1(n581), .A2(n574), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U643 ( .A(G204GAT), .B(n577), .ZN(G1353GAT) );
  NAND2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(G211GAT), .B(n580), .ZN(G1354GAT) );
  NOR2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n584) );
  XNOR2_X1 U647 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n584), .B(n583), .ZN(n585) );
  XOR2_X1 U649 ( .A(n585), .B(KEYINPUT126), .Z(n587) );
  XNOR2_X1 U650 ( .A(G218GAT), .B(KEYINPUT125), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n587), .B(n586), .ZN(G1355GAT) );
endmodule

