//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 1 0 0 1 0 1 0 1 1 1 0 1 1 0 0 0 0 1 0 1 0 1 1 0 0 1 1 1 0 1 0 0 1 1 1 1 1 0 0 1 0 1 1 1 1 0 0 0 1 0 0 0 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:02 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1283, new_n1284;
  XOR2_X1   g0000(.A(KEYINPUT64), .B(G50), .Z(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT65), .Z(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  INV_X1    g0014(.A(new_n202), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G50), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n218), .A2(new_n209), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g0020(.A(KEYINPUT66), .B(G238), .ZN(new_n221));
  INV_X1    g0021(.A(G68), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G107), .A2(G264), .ZN(new_n227));
  NAND4_X1  g0027(.A1(new_n224), .A2(new_n225), .A3(new_n226), .A4(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n211), .B1(new_n223), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n214), .B(new_n220), .C1(KEYINPUT1), .C2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G68), .B(G77), .Z(new_n240));
  XOR2_X1   g0040(.A(G50), .B(G58), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G87), .B(G97), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  NAND3_X1  g0046(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(new_n218), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n203), .A2(G20), .ZN(new_n250));
  XNOR2_X1  g0050(.A(KEYINPUT8), .B(G58), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n209), .A2(G33), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  NOR2_X1   g0054(.A1(G20), .A2(G33), .ZN(new_n255));
  AOI22_X1  g0055(.A1(new_n252), .A2(new_n254), .B1(G150), .B2(new_n255), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n249), .B1(new_n250), .B2(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n259), .A2(new_n248), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n208), .A2(G20), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n260), .A2(G50), .A3(new_n261), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n262), .B1(G50), .B2(new_n258), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n257), .A2(new_n263), .ZN(new_n264));
  OR2_X1    g0064(.A1(KEYINPUT3), .A2(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(KEYINPUT3), .A2(G33), .ZN(new_n266));
  AOI21_X1  g0066(.A(G1698), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G222), .ZN(new_n268));
  INV_X1    g0068(.A(G77), .ZN(new_n269));
  XNOR2_X1  g0069(.A(KEYINPUT3), .B(G33), .ZN(new_n270));
  INV_X1    g0070(.A(G223), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(G1698), .ZN(new_n272));
  OAI221_X1 g0072(.A(new_n268), .B1(new_n269), .B2(new_n270), .C1(new_n271), .C2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(G33), .A2(G41), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n274), .A2(G1), .A3(G13), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n275), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G41), .ZN(new_n281));
  INV_X1    g0081(.A(G45), .ZN(new_n282));
  AOI21_X1  g0082(.A(G1), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  AND2_X1   g0083(.A1(new_n275), .A2(G274), .ZN(new_n284));
  AOI22_X1  g0084(.A1(new_n280), .A2(G226), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n277), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G169), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n264), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n288), .B1(G179), .B2(new_n286), .ZN(new_n289));
  INV_X1    g0089(.A(G190), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n286), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT68), .ZN(new_n292));
  XNOR2_X1  g0092(.A(new_n291), .B(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT9), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n264), .B(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n286), .A2(G200), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT10), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT69), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n299), .B1(new_n296), .B2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  AND3_X1   g0102(.A1(new_n293), .A2(new_n298), .A3(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n302), .B1(new_n293), .B2(new_n298), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n289), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G226), .ZN(new_n306));
  INV_X1    g0106(.A(G1698), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n270), .B(new_n308), .C1(G232), .C2(new_n307), .ZN(new_n309));
  NAND2_X1  g0109(.A1(G33), .A2(G97), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n275), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n283), .A2(new_n275), .A3(G274), .ZN(new_n312));
  INV_X1    g0112(.A(G238), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n312), .B1(new_n313), .B2(new_n279), .ZN(new_n314));
  OAI21_X1  g0114(.A(KEYINPUT13), .B1(new_n311), .B2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT70), .ZN(new_n316));
  XNOR2_X1  g0116(.A(new_n315), .B(new_n316), .ZN(new_n317));
  OR3_X1    g0117(.A1(new_n311), .A2(KEYINPUT13), .A3(new_n314), .ZN(new_n318));
  OR2_X1    g0118(.A1(new_n318), .A2(KEYINPUT71), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(KEYINPUT71), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n317), .A2(new_n319), .A3(G179), .A4(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n318), .A2(new_n315), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(G169), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(KEYINPUT14), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT14), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n322), .A2(new_n325), .A3(G169), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n321), .A2(new_n324), .A3(new_n326), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n260), .A2(G68), .A3(new_n261), .ZN(new_n328));
  XNOR2_X1  g0128(.A(new_n328), .B(KEYINPUT72), .ZN(new_n329));
  AOI22_X1  g0129(.A1(new_n255), .A2(G50), .B1(G20), .B2(new_n222), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n330), .B1(new_n269), .B2(new_n253), .ZN(new_n331));
  AND2_X1   g0131(.A1(new_n331), .A2(new_n248), .ZN(new_n332));
  OR2_X1    g0132(.A1(new_n332), .A2(KEYINPUT11), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n259), .A2(new_n222), .ZN(new_n334));
  XNOR2_X1  g0134(.A(new_n334), .B(KEYINPUT12), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n332), .A2(KEYINPUT11), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n329), .A2(new_n333), .A3(new_n335), .A4(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n327), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(G244), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n312), .B1(new_n339), .B2(new_n279), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n270), .A2(G232), .A3(new_n307), .ZN(new_n341));
  INV_X1    g0141(.A(G107), .ZN(new_n342));
  OAI221_X1 g0142(.A(new_n341), .B1(new_n342), .B2(new_n270), .C1(new_n272), .C2(new_n221), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n340), .B1(new_n343), .B2(new_n276), .ZN(new_n344));
  OAI21_X1  g0144(.A(KEYINPUT67), .B1(new_n344), .B2(G169), .ZN(new_n345));
  INV_X1    g0145(.A(new_n344), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n345), .B1(G179), .B2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(G179), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n344), .A2(KEYINPUT67), .A3(new_n348), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n252), .A2(new_n255), .B1(G20), .B2(G77), .ZN(new_n350));
  XNOR2_X1  g0150(.A(KEYINPUT15), .B(G87), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n350), .B1(new_n253), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n248), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n269), .B1(new_n208), .B2(G20), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n260), .A2(new_n354), .B1(new_n269), .B2(new_n259), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  AND2_X1   g0156(.A1(new_n349), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n347), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n356), .B1(new_n346), .B2(G200), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n359), .B1(new_n290), .B2(new_n346), .ZN(new_n360));
  AND2_X1   g0160(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n317), .A2(new_n319), .A3(G190), .A4(new_n320), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n337), .B1(G200), .B2(new_n322), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n338), .A2(new_n361), .A3(new_n364), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n305), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT18), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n251), .B1(new_n208), .B2(G20), .ZN(new_n368));
  AOI22_X1  g0168(.A1(new_n368), .A2(new_n260), .B1(new_n259), .B2(new_n251), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n265), .A2(new_n209), .A3(new_n266), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT7), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT73), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n265), .A2(KEYINPUT7), .A3(new_n209), .A4(new_n266), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n373), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n375), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(KEYINPUT73), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n376), .A2(G68), .A3(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(G58), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n380), .A2(new_n222), .ZN(new_n381));
  OAI21_X1  g0181(.A(G20), .B1(new_n381), .B2(new_n202), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n255), .A2(G159), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n379), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT16), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n222), .B1(new_n373), .B2(new_n375), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n389), .A2(new_n384), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n249), .B1(new_n390), .B2(KEYINPUT16), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n370), .B1(new_n388), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n271), .A2(new_n307), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n306), .A2(G1698), .ZN(new_n394));
  AND2_X1   g0194(.A1(KEYINPUT3), .A2(G33), .ZN(new_n395));
  NOR2_X1   g0195(.A1(KEYINPUT3), .A2(G33), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n393), .B(new_n394), .C1(new_n395), .C2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(G33), .A2(G87), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n275), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n275), .A2(G232), .A3(new_n278), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n312), .A2(new_n400), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(G179), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n403), .B1(new_n287), .B2(new_n402), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n367), .B1(new_n392), .B2(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(KEYINPUT16), .B1(new_n379), .B2(new_n385), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n395), .A2(new_n396), .ZN(new_n408));
  AOI21_X1  g0208(.A(KEYINPUT7), .B1(new_n408), .B2(new_n209), .ZN(new_n409));
  OAI21_X1  g0209(.A(G68), .B1(new_n409), .B2(new_n377), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n410), .A2(KEYINPUT16), .A3(new_n385), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n248), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n369), .B1(new_n407), .B2(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n413), .A2(new_n404), .A3(KEYINPUT18), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n406), .A2(KEYINPUT74), .A3(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(G200), .ZN(new_n416));
  INV_X1    g0216(.A(new_n399), .ZN(new_n417));
  INV_X1    g0217(.A(new_n401), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n416), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NOR3_X1   g0219(.A1(new_n399), .A2(new_n401), .A3(new_n290), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n421), .B(new_n369), .C1(new_n407), .C2(new_n412), .ZN(new_n422));
  XNOR2_X1  g0222(.A(new_n422), .B(KEYINPUT17), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT74), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n424), .B(new_n367), .C1(new_n392), .C2(new_n405), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n415), .A2(new_n423), .A3(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n366), .A2(new_n427), .ZN(new_n428));
  XNOR2_X1  g0228(.A(new_n428), .B(KEYINPUT75), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n209), .B(G68), .C1(new_n395), .C2(new_n396), .ZN(new_n430));
  OR2_X1    g0230(.A1(KEYINPUT76), .A2(G97), .ZN(new_n431));
  NAND2_X1  g0231(.A1(KEYINPUT76), .A2(G97), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n253), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n430), .B1(new_n433), .B2(KEYINPUT19), .ZN(new_n434));
  NOR2_X1   g0234(.A1(G87), .A2(G107), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n431), .A2(new_n432), .A3(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT19), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n209), .B1(new_n310), .B2(new_n437), .ZN(new_n438));
  AND2_X1   g0238(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n248), .B1(new_n434), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n351), .A2(new_n259), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n208), .A2(G33), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n258), .A2(new_n442), .A3(new_n218), .A4(new_n247), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(G87), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n440), .A2(new_n441), .A3(new_n445), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n282), .A2(G1), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n275), .A2(G274), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n208), .A2(G45), .ZN(new_n449));
  AND2_X1   g0249(.A1(G33), .A2(G41), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n449), .B(G250), .C1(new_n450), .C2(new_n218), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n448), .A2(new_n451), .ZN(new_n452));
  OAI211_X1 g0252(.A(G244), .B(G1698), .C1(new_n395), .C2(new_n396), .ZN(new_n453));
  OAI211_X1 g0253(.A(G238), .B(new_n307), .C1(new_n395), .C2(new_n396), .ZN(new_n454));
  NAND2_X1  g0254(.A1(G33), .A2(G116), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  AOI211_X1 g0256(.A(new_n290), .B(new_n452), .C1(new_n276), .C2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n276), .ZN(new_n458));
  INV_X1    g0258(.A(new_n452), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n416), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NOR3_X1   g0260(.A1(new_n446), .A2(new_n457), .A3(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n351), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n444), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n440), .A2(new_n441), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(KEYINPUT80), .ZN(new_n465));
  AND2_X1   g0265(.A1(KEYINPUT76), .A2(G97), .ZN(new_n466));
  NOR2_X1   g0266(.A1(KEYINPUT76), .A2(G97), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n437), .B1(new_n468), .B2(new_n253), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n436), .A2(new_n438), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n469), .A2(new_n470), .A3(new_n430), .ZN(new_n471));
  AOI22_X1  g0271(.A1(new_n471), .A2(new_n248), .B1(new_n259), .B2(new_n351), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT80), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n472), .A2(new_n473), .A3(new_n463), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n465), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n452), .B1(new_n456), .B2(new_n276), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n476), .A2(G169), .ZN(new_n477));
  AOI211_X1 g0277(.A(G179), .B(new_n452), .C1(new_n276), .C2(new_n456), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n461), .B1(new_n475), .B2(new_n479), .ZN(new_n480));
  AND3_X1   g0280(.A1(KEYINPUT79), .A2(G33), .A3(G283), .ZN(new_n481));
  AOI21_X1  g0281(.A(KEYINPUT79), .B1(G33), .B2(G283), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n307), .B1(new_n265), .B2(new_n266), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n483), .B1(new_n484), .B2(G250), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT78), .ZN(new_n486));
  OAI211_X1 g0286(.A(G244), .B(new_n307), .C1(new_n395), .C2(new_n396), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT4), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n267), .A2(KEYINPUT78), .A3(KEYINPUT4), .A4(G244), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n485), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT77), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n487), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n270), .A2(KEYINPUT77), .A3(G244), .A4(new_n307), .ZN(new_n494));
  AND3_X1   g0294(.A1(new_n493), .A2(new_n494), .A3(new_n488), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n276), .B1(new_n491), .B2(new_n495), .ZN(new_n496));
  XNOR2_X1  g0296(.A(KEYINPUT5), .B(G41), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n276), .B1(new_n447), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(G257), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n284), .A2(new_n447), .A3(new_n497), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n496), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n287), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n376), .A2(G107), .A3(new_n378), .ZN(new_n505));
  XOR2_X1   g0305(.A(G97), .B(G107), .Z(new_n506));
  NAND2_X1  g0306(.A1(new_n342), .A2(KEYINPUT6), .ZN(new_n507));
  OAI22_X1  g0307(.A1(new_n506), .A2(KEYINPUT6), .B1(new_n468), .B2(new_n507), .ZN(new_n508));
  AOI22_X1  g0308(.A1(new_n508), .A2(G20), .B1(G77), .B2(new_n255), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n505), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(new_n248), .ZN(new_n511));
  INV_X1    g0311(.A(G97), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n259), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n513), .B1(new_n443), .B2(new_n512), .ZN(new_n514));
  INV_X1    g0314(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n511), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n493), .A2(new_n494), .A3(new_n488), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n517), .A2(new_n490), .A3(new_n489), .A4(new_n485), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n501), .B1(new_n518), .B2(new_n276), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(new_n348), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n504), .A2(new_n516), .A3(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n496), .A2(G190), .A3(new_n502), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n514), .B1(new_n510), .B2(new_n248), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n522), .B(new_n523), .C1(new_n416), .C2(new_n519), .ZN(new_n524));
  AND3_X1   g0324(.A1(new_n480), .A2(new_n521), .A3(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT82), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT21), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n258), .A2(G116), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n528), .B1(new_n444), .B2(G116), .ZN(new_n529));
  INV_X1    g0329(.A(G33), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n530), .B1(new_n466), .B2(new_n467), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n531), .B(new_n209), .C1(new_n482), .C2(new_n481), .ZN(new_n532));
  INV_X1    g0332(.A(G116), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n247), .A2(new_n218), .B1(G20), .B2(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(KEYINPUT20), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n209), .B1(new_n481), .B2(new_n482), .ZN(new_n536));
  AOI21_X1  g0336(.A(G33), .B1(new_n431), .B2(new_n432), .ZN(new_n537));
  OAI211_X1 g0337(.A(KEYINPUT20), .B(new_n534), .C1(new_n536), .C2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n529), .B1(new_n535), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(G169), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n497), .A2(new_n447), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n542), .A2(G270), .A3(new_n275), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n500), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n270), .A2(G264), .A3(G1698), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n408), .A2(G303), .ZN(new_n546));
  OAI211_X1 g0346(.A(G257), .B(new_n307), .C1(new_n395), .C2(new_n396), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT81), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n275), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n545), .A2(new_n546), .A3(KEYINPUT81), .A4(new_n547), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n544), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n526), .B(new_n527), .C1(new_n541), .C2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n550), .A2(new_n551), .ZN(new_n554));
  INV_X1    g0354(.A(new_n544), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n526), .A2(new_n527), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n556), .A2(G169), .A3(new_n557), .A4(new_n540), .ZN(new_n558));
  AOI211_X1 g0358(.A(new_n348), .B(new_n544), .C1(new_n550), .C2(new_n551), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n540), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n553), .A2(new_n558), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(KEYINPUT25), .B1(new_n259), .B2(new_n342), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n259), .A2(KEYINPUT25), .A3(new_n342), .ZN(new_n564));
  AOI22_X1  g0364(.A1(new_n563), .A2(new_n564), .B1(G107), .B2(new_n444), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n270), .A2(new_n209), .A3(G87), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(KEYINPUT22), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT22), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n270), .A2(new_n568), .A3(new_n209), .A4(G87), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT83), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n571), .B1(new_n209), .B2(G107), .ZN(new_n572));
  OR2_X1    g0372(.A1(new_n572), .A2(KEYINPUT23), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(KEYINPUT23), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n573), .A2(new_n574), .B1(G116), .B2(new_n254), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n570), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(KEYINPUT24), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT24), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n570), .A2(new_n578), .A3(new_n575), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g0380(.A(KEYINPUT84), .B1(new_n580), .B2(new_n248), .ZN(new_n581));
  AND3_X1   g0381(.A1(new_n570), .A2(new_n578), .A3(new_n575), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n578), .B1(new_n570), .B2(new_n575), .ZN(new_n583));
  OAI211_X1 g0383(.A(KEYINPUT84), .B(new_n248), .C1(new_n582), .C2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n584), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n565), .B1(new_n581), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n270), .A2(G257), .A3(G1698), .ZN(new_n587));
  NAND2_X1  g0387(.A1(G33), .A2(G294), .ZN(new_n588));
  OAI211_X1 g0388(.A(G250), .B(new_n307), .C1(new_n395), .C2(new_n396), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n276), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n498), .A2(G264), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n591), .A2(new_n500), .A3(new_n592), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n593), .A2(G179), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n594), .B1(new_n287), .B2(new_n593), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n561), .B1(new_n586), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n556), .A2(new_n290), .ZN(new_n597));
  INV_X1    g0397(.A(new_n540), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n598), .B1(new_n552), .B2(new_n416), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(new_n565), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n248), .B1(new_n582), .B2(new_n583), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT84), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n601), .B1(new_n604), .B2(new_n584), .ZN(new_n605));
  OR3_X1    g0405(.A1(new_n593), .A2(KEYINPUT85), .A3(G190), .ZN(new_n606));
  OAI21_X1  g0406(.A(KEYINPUT85), .B1(new_n593), .B2(G190), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n593), .A2(new_n416), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n600), .B1(new_n605), .B2(new_n609), .ZN(new_n610));
  AND4_X1   g0410(.A1(new_n429), .A2(new_n525), .A3(new_n596), .A4(new_n610), .ZN(G372));
  XNOR2_X1  g0411(.A(KEYINPUT88), .B(KEYINPUT18), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n413), .A2(new_n404), .A3(KEYINPUT87), .ZN(new_n614));
  INV_X1    g0414(.A(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(KEYINPUT87), .B1(new_n413), .B2(new_n404), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n613), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n616), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n618), .A2(new_n614), .A3(new_n612), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  AND2_X1   g0421(.A1(new_n362), .A2(new_n363), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n338), .B1(new_n358), .B2(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n621), .B1(new_n423), .B2(new_n623), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n303), .A2(new_n304), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n289), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n605), .A2(new_n609), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n586), .A2(new_n595), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n525), .B(new_n627), .C1(new_n629), .C2(new_n561), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT26), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n464), .A2(KEYINPUT80), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n473), .B1(new_n472), .B2(new_n463), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n479), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n461), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n631), .B1(new_n636), .B2(new_n521), .ZN(new_n637));
  AND3_X1   g0437(.A1(new_n496), .A2(new_n348), .A3(new_n502), .ZN(new_n638));
  AOI21_X1  g0438(.A(G169), .B1(new_n496), .B2(new_n502), .ZN(new_n639));
  NOR3_X1   g0439(.A1(new_n638), .A2(new_n639), .A3(new_n523), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n640), .A2(new_n480), .A3(KEYINPUT26), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n637), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(KEYINPUT86), .B1(new_n642), .B2(new_n634), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT86), .ZN(new_n644));
  INV_X1    g0444(.A(new_n634), .ZN(new_n645));
  AOI211_X1 g0445(.A(new_n644), .B(new_n645), .C1(new_n637), .C2(new_n641), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n630), .B1(new_n643), .B2(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n626), .B1(new_n429), .B2(new_n647), .ZN(new_n648));
  XNOR2_X1  g0448(.A(new_n648), .B(KEYINPUT89), .ZN(G369));
  NAND3_X1  g0449(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n650));
  OR2_X1    g0450(.A1(new_n650), .A2(KEYINPUT27), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(KEYINPUT27), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n651), .A2(G213), .A3(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(G343), .ZN(new_n655));
  XNOR2_X1  g0455(.A(new_n655), .B(KEYINPUT90), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n656), .A2(new_n598), .ZN(new_n657));
  XNOR2_X1  g0457(.A(new_n561), .B(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n658), .B1(new_n597), .B2(new_n599), .ZN(new_n659));
  XOR2_X1   g0459(.A(new_n659), .B(KEYINPUT91), .Z(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(G330), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n627), .B1(new_n605), .B2(new_n656), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(new_n628), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n629), .A2(new_n656), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n561), .A2(new_n656), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n669), .B1(new_n629), .B2(new_n656), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n667), .A2(new_n670), .ZN(G399));
  INV_X1    g0471(.A(new_n212), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n672), .A2(G41), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(G1), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n468), .A2(new_n533), .A3(new_n435), .ZN(new_n676));
  OAI22_X1  g0476(.A1(new_n675), .A2(new_n676), .B1(new_n216), .B2(new_n674), .ZN(new_n677));
  XNOR2_X1  g0477(.A(new_n677), .B(KEYINPUT28), .ZN(new_n678));
  INV_X1    g0478(.A(new_n656), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n645), .B1(new_n637), .B2(new_n641), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n679), .B1(new_n630), .B2(new_n680), .ZN(new_n681));
  AND2_X1   g0481(.A1(new_n681), .A2(KEYINPUT29), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT29), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n647), .A2(new_n656), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n682), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n596), .A2(new_n525), .A3(new_n610), .A4(new_n656), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT30), .ZN(new_n687));
  AND3_X1   g0487(.A1(new_n476), .A2(new_n591), .A3(new_n592), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n519), .A2(new_n688), .A3(G179), .A4(new_n552), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n476), .A2(G179), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(new_n593), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n691), .A2(new_n552), .ZN(new_n692));
  AOI22_X1  g0492(.A1(new_n687), .A2(new_n689), .B1(new_n692), .B2(new_n503), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n559), .A2(KEYINPUT30), .A3(new_n519), .A4(new_n688), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n656), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(KEYINPUT31), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n689), .A2(new_n687), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n692), .A2(new_n503), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(new_n694), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(new_n679), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT31), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n686), .A2(new_n696), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(G330), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n685), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n678), .B1(new_n706), .B2(G1), .ZN(G364));
  NOR2_X1   g0507(.A1(new_n660), .A2(G330), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n209), .A2(G13), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n208), .B1(new_n709), .B2(G45), .ZN(new_n710));
  AOI211_X1 g0510(.A(new_n708), .B(new_n662), .C1(new_n674), .C2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n710), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n673), .A2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n212), .A2(G116), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n672), .A2(new_n270), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n716), .B1(G45), .B2(new_n216), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n717), .B1(G45), .B2(new_n242), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n672), .A2(new_n408), .ZN(new_n719));
  AOI211_X1 g0519(.A(new_n715), .B(new_n718), .C1(G355), .C2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(G13), .A2(G33), .ZN(new_n722));
  XNOR2_X1  g0522(.A(new_n722), .B(KEYINPUT92), .ZN(new_n723));
  OR2_X1    g0523(.A1(new_n723), .A2(G20), .ZN(new_n724));
  XOR2_X1   g0524(.A(new_n724), .B(KEYINPUT93), .Z(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n218), .B1(G20), .B2(new_n287), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n714), .B1(new_n721), .B2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n209), .A2(new_n348), .ZN(new_n730));
  NOR2_X1   g0530(.A1(G190), .A2(G200), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n290), .A2(G200), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  OAI221_X1 g0534(.A(new_n270), .B1(new_n732), .B2(new_n269), .C1(new_n380), .C2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT32), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n209), .A2(G179), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(new_n731), .ZN(new_n738));
  INV_X1    g0538(.A(G159), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n736), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n738), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n741), .A2(KEYINPUT32), .A3(G159), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n735), .B1(new_n740), .B2(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n209), .B1(new_n733), .B2(new_n348), .ZN(new_n744));
  XOR2_X1   g0544(.A(new_n744), .B(KEYINPUT94), .Z(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(G97), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n737), .A2(G190), .A3(G200), .ZN(new_n747));
  INV_X1    g0547(.A(G87), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n730), .A2(G200), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(G190), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n749), .B1(G68), .B2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n750), .A2(new_n290), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n737), .A2(new_n290), .A3(G200), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  AOI22_X1  g0555(.A1(new_n753), .A2(G50), .B1(new_n755), .B2(G107), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n743), .A2(new_n746), .A3(new_n752), .A4(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT95), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(G303), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n408), .B1(new_n747), .B2(new_n760), .ZN(new_n761));
  XNOR2_X1  g0561(.A(new_n761), .B(KEYINPUT96), .ZN(new_n762));
  INV_X1    g0562(.A(G311), .ZN(new_n763));
  INV_X1    g0563(.A(G329), .ZN(new_n764));
  OAI22_X1  g0564(.A1(new_n732), .A2(new_n763), .B1(new_n738), .B2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n734), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n765), .B1(G322), .B2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n744), .ZN(new_n768));
  AOI22_X1  g0568(.A1(G326), .A2(new_n753), .B1(new_n768), .B2(G294), .ZN(new_n769));
  XNOR2_X1  g0569(.A(KEYINPUT33), .B(G317), .ZN(new_n770));
  AOI22_X1  g0570(.A1(new_n751), .A2(new_n770), .B1(new_n755), .B2(G283), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n767), .A2(new_n769), .A3(new_n771), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n759), .B1(new_n762), .B2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n757), .A2(new_n758), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n727), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n729), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n776), .B1(new_n659), .B2(new_n726), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n711), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(G396));
  NAND3_X1  g0579(.A1(new_n647), .A2(new_n361), .A3(new_n656), .ZN(new_n780));
  INV_X1    g0580(.A(new_n684), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n679), .A2(new_n356), .ZN(new_n782));
  AND3_X1   g0582(.A1(new_n358), .A2(new_n360), .A3(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n782), .B1(new_n358), .B2(new_n360), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT99), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n780), .B1(new_n781), .B2(new_n786), .ZN(new_n787));
  OR2_X1    g0587(.A1(new_n787), .A2(new_n704), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n713), .B1(new_n787), .B2(new_n704), .ZN(new_n789));
  AND2_X1   g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  OR2_X1    g0590(.A1(new_n727), .A2(new_n722), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n713), .B1(G77), .B2(new_n791), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n732), .A2(new_n533), .B1(new_n738), .B2(new_n763), .ZN(new_n793));
  AOI211_X1 g0593(.A(new_n270), .B(new_n793), .C1(G294), .C2(new_n766), .ZN(new_n794));
  INV_X1    g0594(.A(new_n747), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n753), .A2(G303), .B1(new_n795), .B2(G107), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n754), .A2(new_n748), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n797), .B1(G283), .B2(new_n751), .ZN(new_n798));
  NAND4_X1  g0598(.A1(new_n794), .A2(new_n746), .A3(new_n796), .A4(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n754), .A2(new_n222), .ZN(new_n800));
  AOI211_X1 g0600(.A(new_n408), .B(new_n800), .C1(G132), .C2(new_n741), .ZN(new_n801));
  AOI22_X1  g0601(.A1(G58), .A2(new_n768), .B1(new_n795), .B2(G50), .ZN(new_n802));
  INV_X1    g0602(.A(new_n732), .ZN(new_n803));
  AOI22_X1  g0603(.A1(G143), .A2(new_n766), .B1(new_n803), .B2(G159), .ZN(new_n804));
  INV_X1    g0604(.A(new_n751), .ZN(new_n805));
  INV_X1    g0605(.A(G150), .ZN(new_n806));
  INV_X1    g0606(.A(G137), .ZN(new_n807));
  INV_X1    g0607(.A(new_n753), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n804), .B1(new_n805), .B2(new_n806), .C1(new_n807), .C2(new_n808), .ZN(new_n809));
  XNOR2_X1  g0609(.A(KEYINPUT97), .B(KEYINPUT34), .ZN(new_n810));
  OAI211_X1 g0610(.A(new_n801), .B(new_n802), .C1(new_n809), .C2(new_n810), .ZN(new_n811));
  AND2_X1   g0611(.A1(new_n809), .A2(new_n810), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n799), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n792), .B1(new_n813), .B2(new_n727), .ZN(new_n814));
  INV_X1    g0614(.A(new_n785), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n814), .B1(new_n815), .B2(new_n723), .ZN(new_n816));
  XOR2_X1   g0616(.A(new_n816), .B(KEYINPUT98), .Z(new_n817));
  NOR2_X1   g0617(.A1(new_n790), .A2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(G384));
  OR2_X1    g0619(.A1(new_n508), .A2(KEYINPUT35), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n508), .A2(KEYINPUT35), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n820), .A2(G116), .A3(new_n219), .A4(new_n821), .ZN(new_n822));
  XOR2_X1   g0622(.A(new_n822), .B(KEYINPUT36), .Z(new_n823));
  OR3_X1    g0623(.A1(new_n216), .A2(new_n269), .A3(new_n381), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n201), .A2(G68), .ZN(new_n825));
  AOI211_X1 g0625(.A(new_n208), .B(G13), .C1(new_n824), .C2(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n823), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n338), .A2(new_n679), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT39), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n387), .B1(new_n389), .B2(new_n384), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n830), .A2(new_n411), .A3(new_n248), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(new_n369), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(new_n404), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(new_n422), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n834), .A2(KEYINPUT101), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT101), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n833), .A2(new_n836), .A3(new_n422), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n832), .A2(new_n654), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n835), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(KEYINPUT37), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n413), .A2(new_n654), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(new_n422), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n392), .A2(new_n405), .ZN(new_n843));
  NOR3_X1   g0643(.A1(new_n842), .A2(new_n843), .A3(KEYINPUT37), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n840), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n838), .ZN(new_n847));
  AND3_X1   g0647(.A1(new_n413), .A2(new_n404), .A3(KEYINPUT18), .ZN(new_n848));
  AOI21_X1  g0648(.A(KEYINPUT18), .B1(new_n413), .B2(new_n404), .ZN(new_n849));
  NOR3_X1   g0649(.A1(new_n848), .A2(new_n849), .A3(new_n424), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT17), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n422), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n392), .A2(KEYINPUT17), .A3(new_n421), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n425), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  OAI211_X1 g0654(.A(KEYINPUT100), .B(new_n847), .C1(new_n850), .C2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(KEYINPUT100), .B1(new_n426), .B2(new_n847), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n846), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT38), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  OAI211_X1 g0660(.A(KEYINPUT38), .B(new_n846), .C1(new_n856), .C2(new_n857), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n829), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n841), .B1(new_n620), .B2(new_n423), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n422), .B(new_n841), .C1(new_n615), .C2(new_n616), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n844), .B1(new_n864), .B2(KEYINPUT37), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n859), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n861), .A2(new_n866), .A3(new_n829), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  NOR3_X1   g0668(.A1(new_n862), .A2(new_n868), .A3(KEYINPUT102), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT102), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n847), .B1(new_n850), .B2(new_n854), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT100), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(new_n855), .ZN(new_n874));
  AOI21_X1  g0674(.A(KEYINPUT38), .B1(new_n874), .B2(new_n846), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n844), .B1(new_n839), .B2(KEYINPUT37), .ZN(new_n876));
  AOI211_X1 g0676(.A(new_n859), .B(new_n876), .C1(new_n873), .C2(new_n855), .ZN(new_n877));
  OAI21_X1  g0677(.A(KEYINPUT39), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n870), .B1(new_n878), .B2(new_n867), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n828), .B1(new_n869), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n679), .A2(new_n337), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n338), .A2(new_n364), .A3(new_n881), .ZN(new_n882));
  OAI211_X1 g0682(.A(new_n337), .B(new_n679), .C1(new_n622), .C2(new_n327), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n358), .A2(new_n679), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n885), .B1(new_n780), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n860), .A2(new_n861), .ZN(new_n889));
  AOI22_X1  g0689(.A1(new_n888), .A2(new_n889), .B1(new_n621), .B2(new_n653), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n880), .A2(KEYINPUT103), .A3(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT103), .ZN(new_n892));
  INV_X1    g0692(.A(new_n828), .ZN(new_n893));
  OAI21_X1  g0693(.A(KEYINPUT102), .B1(new_n862), .B2(new_n868), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n878), .A2(new_n870), .A3(new_n867), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n893), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n890), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n892), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n891), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n626), .B1(new_n429), .B2(new_n685), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n899), .B(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n861), .A2(new_n866), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT104), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n903), .B1(new_n695), .B2(KEYINPUT31), .ZN(new_n904));
  AND4_X1   g0704(.A1(new_n903), .A2(new_n699), .A3(KEYINPUT31), .A4(new_n679), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n686), .B(new_n702), .C1(new_n904), .C2(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n785), .B1(new_n882), .B2(new_n883), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n902), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(KEYINPUT40), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n908), .A2(KEYINPUT105), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT105), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n906), .B(new_n907), .C1(new_n913), .C2(KEYINPUT40), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n912), .B(new_n914), .C1(new_n877), .C2(new_n875), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n911), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n916), .A2(new_n429), .A3(new_n906), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n429), .A2(new_n906), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n918), .A2(new_n911), .A3(new_n915), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n917), .A2(new_n919), .A3(G330), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n901), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(new_n208), .B2(new_n709), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n901), .A2(new_n920), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n827), .B1(new_n922), .B2(new_n923), .ZN(G367));
  NAND2_X1  g0724(.A1(new_n679), .A2(new_n516), .ZN(new_n925));
  NOR3_X1   g0725(.A1(new_n925), .A2(new_n638), .A3(new_n639), .ZN(new_n926));
  AND2_X1   g0726(.A1(new_n926), .A2(KEYINPUT107), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n925), .A2(new_n521), .A3(new_n524), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n926), .A2(KEYINPUT107), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n927), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n669), .A2(new_n930), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n931), .B(KEYINPUT42), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n640), .B1(new_n930), .B2(new_n629), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n656), .B1(new_n933), .B2(KEYINPUT108), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n934), .B1(KEYINPUT108), .B2(new_n933), .ZN(new_n935));
  OR2_X1    g0735(.A1(new_n932), .A2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT109), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n938), .B(KEYINPUT43), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n679), .A2(new_n446), .ZN(new_n940));
  XOR2_X1   g0740(.A(new_n940), .B(KEYINPUT106), .Z(new_n941));
  NOR2_X1   g0741(.A1(new_n941), .A2(new_n645), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n942), .B1(new_n636), .B2(new_n941), .ZN(new_n943));
  AND3_X1   g0743(.A1(new_n939), .A2(new_n943), .A3(new_n936), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n939), .A2(new_n943), .ZN(new_n945));
  INV_X1    g0745(.A(new_n930), .ZN(new_n946));
  OAI22_X1  g0746(.A1(new_n944), .A2(new_n945), .B1(new_n667), .B2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n706), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n670), .A2(new_n930), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(KEYINPUT44), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n670), .A2(new_n930), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT45), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n951), .B(new_n952), .ZN(new_n953));
  AND3_X1   g0753(.A1(new_n950), .A2(new_n667), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n667), .B1(new_n950), .B2(new_n953), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(KEYINPUT110), .B1(new_n666), .B2(new_n668), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n661), .B(new_n957), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(new_n669), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n948), .B1(new_n956), .B2(new_n959), .ZN(new_n960));
  XOR2_X1   g0760(.A(new_n673), .B(KEYINPUT41), .Z(new_n961));
  OAI21_X1  g0761(.A(new_n710), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n939), .A2(new_n943), .A3(new_n936), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n667), .A2(new_n946), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n963), .B(new_n964), .C1(new_n943), .C2(new_n939), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n947), .A2(new_n962), .A3(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(new_n728), .ZN(new_n967));
  INV_X1    g0767(.A(new_n716), .ZN(new_n968));
  OAI22_X1  g0768(.A1(new_n968), .A2(new_n238), .B1(new_n212), .B2(new_n351), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n713), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  OAI22_X1  g0770(.A1(new_n734), .A2(new_n806), .B1(new_n738), .B2(new_n807), .ZN(new_n971));
  INV_X1    g0771(.A(new_n201), .ZN(new_n972));
  AOI211_X1 g0772(.A(new_n408), .B(new_n971), .C1(new_n972), .C2(new_n803), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n745), .A2(G68), .ZN(new_n974));
  AOI22_X1  g0774(.A1(new_n751), .A2(G159), .B1(new_n753), .B2(G143), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n754), .A2(new_n269), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n976), .B1(G58), .B2(new_n795), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n973), .A2(new_n974), .A3(new_n975), .A4(new_n977), .ZN(new_n978));
  AOI22_X1  g0778(.A1(G294), .A2(new_n751), .B1(new_n768), .B2(G107), .ZN(new_n979));
  INV_X1    g0779(.A(new_n468), .ZN(new_n980));
  AOI22_X1  g0780(.A1(new_n753), .A2(G311), .B1(new_n755), .B2(new_n980), .ZN(new_n981));
  AOI22_X1  g0781(.A1(G283), .A2(new_n803), .B1(new_n766), .B2(G303), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n270), .B1(new_n741), .B2(G317), .ZN(new_n983));
  NAND4_X1  g0783(.A1(new_n979), .A2(new_n981), .A3(new_n982), .A4(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n747), .A2(new_n533), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(KEYINPUT46), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n978), .B1(new_n984), .B2(new_n986), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT47), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n970), .B1(new_n988), .B2(new_n727), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(new_n943), .B2(new_n725), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n966), .A2(new_n990), .ZN(G387));
  NAND2_X1  g0791(.A1(new_n959), .A2(new_n712), .ZN(new_n992));
  INV_X1    g0792(.A(G50), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n270), .B1(new_n738), .B2(new_n806), .C1(new_n734), .C2(new_n993), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n808), .A2(new_n739), .B1(new_n747), .B2(new_n269), .ZN(new_n995));
  AOI211_X1 g0795(.A(new_n994), .B(new_n995), .C1(G97), .C2(new_n755), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n751), .A2(new_n252), .B1(new_n803), .B2(G68), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT112), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n745), .A2(new_n462), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n996), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n270), .B1(new_n741), .B2(G326), .ZN(new_n1001));
  INV_X1    g0801(.A(G283), .ZN(new_n1002));
  INV_X1    g0802(.A(G294), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n744), .A2(new_n1002), .B1(new_n747), .B2(new_n1003), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(G303), .A2(new_n803), .B1(new_n766), .B2(G317), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n753), .A2(G322), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n1005), .B(new_n1006), .C1(new_n763), .C2(new_n805), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT48), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1004), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(new_n1008), .B2(new_n1007), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT49), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n1001), .B1(new_n533), .B2(new_n754), .C1(new_n1010), .C2(new_n1011), .ZN(new_n1012));
  AND2_X1   g0812(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1000), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(new_n727), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n719), .A2(new_n676), .B1(new_n342), .B2(new_n672), .ZN(new_n1016));
  AOI211_X1 g0816(.A(G45), .B(new_n676), .C1(G68), .C2(G77), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n251), .A2(G50), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT50), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n968), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT111), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n1020), .A2(new_n1021), .B1(new_n282), .B2(new_n235), .ZN(new_n1022));
  AND2_X1   g0822(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1016), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n714), .B1(new_n1024), .B2(new_n728), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n1015), .B(new_n1025), .C1(new_n666), .C2(new_n725), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n959), .A2(new_n706), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1027), .A2(new_n673), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n959), .A2(new_n706), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n992), .B(new_n1026), .C1(new_n1028), .C2(new_n1029), .ZN(G393));
  NAND3_X1  g0830(.A1(new_n956), .A2(new_n706), .A3(new_n959), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1027), .B1(new_n954), .B2(new_n955), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1031), .A2(new_n673), .A3(new_n1032), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n753), .A2(G150), .B1(new_n766), .B2(G159), .ZN(new_n1034));
  XOR2_X1   g0834(.A(new_n1034), .B(KEYINPUT51), .Z(new_n1035));
  NAND2_X1  g0835(.A1(new_n745), .A2(G77), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n408), .B1(new_n741), .B2(G143), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n251), .B2(new_n732), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n1038), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n747), .A2(new_n222), .ZN(new_n1040));
  AOI211_X1 g0840(.A(new_n797), .B(new_n1040), .C1(new_n972), .C2(new_n751), .ZN(new_n1041));
  NAND4_X1  g0841(.A1(new_n1035), .A2(new_n1036), .A3(new_n1039), .A4(new_n1041), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n753), .A2(G317), .B1(new_n766), .B2(G311), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n1043), .B(KEYINPUT52), .Z(new_n1044));
  NOR2_X1   g0844(.A1(new_n732), .A2(new_n1003), .ZN(new_n1045));
  AOI211_X1 g0845(.A(new_n270), .B(new_n1045), .C1(G322), .C2(new_n741), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n751), .A2(G303), .B1(new_n755), .B2(G107), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(G116), .A2(new_n768), .B1(new_n795), .B2(G283), .ZN(new_n1048));
  NAND4_X1  g0848(.A1(new_n1044), .A2(new_n1046), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1049), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1042), .B1(new_n1050), .B2(KEYINPUT113), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT113), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n1049), .A2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n727), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n716), .A2(new_n245), .B1(new_n672), .B2(new_n980), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n714), .B1(new_n728), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n1057), .B(KEYINPUT114), .Z(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(new_n726), .B2(new_n946), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(new_n956), .B2(new_n712), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1033), .A2(new_n1060), .ZN(G390));
  NAND2_X1  g0861(.A1(new_n780), .A2(new_n887), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1062), .A2(new_n884), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT115), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1063), .A2(new_n1064), .A3(new_n893), .ZN(new_n1065));
  OAI21_X1  g0865(.A(KEYINPUT115), .B1(new_n888), .B2(new_n828), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n1065), .A2(new_n894), .A3(new_n1066), .A4(new_n895), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n886), .B1(new_n681), .B2(new_n361), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n902), .B(new_n893), .C1(new_n1068), .C2(new_n885), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n906), .A2(G330), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(new_n907), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1070), .A2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n705), .A2(new_n815), .A3(new_n884), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1067), .A2(new_n1069), .A3(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n429), .A2(new_n1072), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1076), .A2(new_n1068), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1072), .A2(KEYINPUT116), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT116), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1071), .A2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1081), .A2(new_n786), .A3(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1080), .B1(new_n1084), .B2(new_n885), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n885), .B1(new_n704), .B2(new_n785), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1073), .A2(new_n1086), .ZN(new_n1087));
  AND2_X1   g0887(.A1(new_n1087), .A2(new_n1062), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n900), .B(new_n1079), .C1(new_n1085), .C2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1078), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1089), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1075), .A2(new_n1091), .A3(new_n1077), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1090), .A2(new_n673), .A3(new_n1092), .ZN(new_n1093));
  AND3_X1   g0893(.A1(new_n1067), .A2(new_n1069), .A3(new_n1076), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1073), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n712), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n713), .B1(new_n252), .B2(new_n791), .ZN(new_n1098));
  INV_X1    g0898(.A(G128), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n1099), .A2(new_n808), .B1(new_n805), .B2(new_n807), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1100), .B1(new_n972), .B2(new_n755), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(KEYINPUT54), .B(G143), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n732), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(G132), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n270), .B1(new_n734), .B2(new_n1104), .ZN(new_n1105));
  AOI211_X1 g0905(.A(new_n1103), .B(new_n1105), .C1(G125), .C2(new_n741), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n745), .A2(G159), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n747), .A2(new_n806), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(new_n1108), .B(new_n1109), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n1101), .A2(new_n1106), .A3(new_n1107), .A4(new_n1110), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1036), .B1(new_n533), .B2(new_n734), .ZN(new_n1112));
  XOR2_X1   g0912(.A(new_n1112), .B(KEYINPUT119), .Z(new_n1113));
  NOR2_X1   g0913(.A1(new_n749), .A2(new_n270), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n1114), .B(KEYINPUT118), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n732), .A2(new_n468), .B1(new_n738), .B2(new_n1003), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n342), .A2(new_n805), .B1(new_n808), .B2(new_n1002), .ZN(new_n1117));
  OR4_X1    g0917(.A1(new_n800), .A2(new_n1115), .A3(new_n1116), .A4(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1111), .B1(new_n1113), .B2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1098), .B1(new_n1119), .B2(new_n727), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n869), .A2(new_n879), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1120), .B1(new_n1122), .B2(new_n723), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1093), .A2(new_n1097), .A3(new_n1123), .ZN(G378));
  OAI21_X1  g0924(.A(new_n713), .B1(new_n972), .B2(new_n791), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n993), .B1(G33), .B2(G41), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1126), .B1(new_n408), .B2(new_n281), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n512), .A2(new_n805), .B1(new_n808), .B2(new_n533), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n380), .A2(new_n754), .B1(new_n747), .B2(new_n269), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  AOI211_X1 g0930(.A(G41), .B(new_n270), .C1(new_n741), .C2(G283), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(G107), .A2(new_n766), .B1(new_n803), .B2(new_n462), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1130), .A2(new_n974), .A3(new_n1131), .A4(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT58), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1127), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n734), .A2(new_n1099), .B1(new_n732), .B2(new_n807), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(G132), .B2(new_n751), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1102), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n753), .A2(G125), .B1(new_n795), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n745), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n1137), .B(new_n1139), .C1(new_n1140), .C2(new_n806), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(KEYINPUT59), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n755), .A2(G159), .ZN(new_n1143));
  AOI211_X1 g0943(.A(G33), .B(G41), .C1(new_n741), .C2(G124), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1142), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1141), .A2(KEYINPUT59), .ZN(new_n1146));
  OAI221_X1 g0946(.A(new_n1135), .B1(new_n1134), .B2(new_n1133), .C1(new_n1145), .C2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1125), .B1(new_n1147), .B2(new_n727), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n264), .A2(new_n653), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n305), .A2(new_n1149), .ZN(new_n1150));
  OAI221_X1 g0950(.A(new_n289), .B1(new_n264), .B2(new_n653), .C1(new_n303), .C2(new_n304), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1152));
  AND3_X1   g0952(.A1(new_n1150), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1152), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1148), .B1(new_n1156), .B2(new_n723), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(new_n1157), .B(KEYINPUT120), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1156), .B1(new_n916), .B2(G330), .ZN(new_n1160));
  INV_X1    g0960(.A(G330), .ZN(new_n1161));
  AOI211_X1 g0961(.A(new_n1161), .B(new_n1155), .C1(new_n911), .C2(new_n915), .ZN(new_n1162));
  OR2_X1    g0962(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(KEYINPUT103), .B1(new_n880), .B2(new_n890), .ZN(new_n1164));
  NOR3_X1   g0964(.A1(new_n896), .A2(new_n892), .A3(new_n897), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1163), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n891), .A2(new_n1167), .A3(new_n898), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1159), .B1(new_n1169), .B2(new_n710), .ZN(new_n1170));
  NOR3_X1   g0970(.A1(new_n1094), .A2(new_n1095), .A3(new_n1089), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n900), .A2(new_n1079), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1168), .B(new_n1166), .C1(new_n1171), .C2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT57), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n674), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  AND3_X1   g0975(.A1(new_n891), .A2(new_n1167), .A3(new_n898), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1167), .B1(new_n898), .B2(new_n891), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1172), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1092), .A2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1178), .A2(KEYINPUT57), .A3(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1170), .B1(new_n1175), .B2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(G375));
  OR2_X1    g0983(.A1(new_n1085), .A2(new_n1088), .ZN(new_n1184));
  XOR2_X1   g0984(.A(new_n710), .B(KEYINPUT121), .Z(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n885), .A2(new_n722), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n713), .B1(G68), .B2(new_n791), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(new_n1188), .B(KEYINPUT122), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n734), .A2(new_n1002), .B1(new_n732), .B2(new_n342), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n270), .B(new_n1190), .C1(G303), .C2(new_n741), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n976), .B1(G116), .B2(new_n751), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n753), .A2(G294), .B1(new_n795), .B2(G97), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1191), .A2(new_n999), .A3(new_n1192), .A4(new_n1193), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n751), .A2(new_n1138), .B1(new_n755), .B2(G58), .ZN(new_n1195));
  OAI221_X1 g0995(.A(new_n1195), .B1(new_n739), .B2(new_n747), .C1(new_n1140), .C2(new_n993), .ZN(new_n1196));
  OR3_X1    g0996(.A1(new_n808), .A2(KEYINPUT123), .A3(new_n1104), .ZN(new_n1197));
  OAI21_X1  g0997(.A(KEYINPUT123), .B1(new_n808), .B2(new_n1104), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n408), .B1(new_n803), .B2(G150), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(G137), .A2(new_n766), .B1(new_n741), .B2(G128), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1197), .A2(new_n1198), .A3(new_n1199), .A4(new_n1200), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1194), .B1(new_n1196), .B2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1189), .B1(new_n1202), .B2(new_n727), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n1184), .A2(new_n1186), .B1(new_n1187), .B2(new_n1203), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1184), .A2(new_n1179), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n961), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1089), .A2(new_n1206), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1204), .B1(new_n1205), .B2(new_n1207), .ZN(G381));
  INV_X1    g1008(.A(G390), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1209), .A2(new_n818), .ZN(new_n1210));
  OR4_X1    g1010(.A1(G396), .A2(new_n1210), .A3(G393), .A4(G381), .ZN(new_n1211));
  INV_X1    g1011(.A(G378), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1182), .A2(new_n1212), .ZN(new_n1213));
  OR3_X1    g1013(.A1(new_n1211), .A2(G387), .A3(new_n1213), .ZN(G407));
  OAI211_X1 g1014(.A(G407), .B(G213), .C1(G343), .C2(new_n1213), .ZN(G409));
  XNOR2_X1  g1015(.A(G393), .B(new_n778), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  AND3_X1   g1017(.A1(new_n966), .A2(new_n990), .A3(G390), .ZN(new_n1218));
  AOI21_X1  g1018(.A(G390), .B1(new_n966), .B2(new_n990), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1217), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(G387), .A2(new_n1209), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n966), .A2(new_n990), .A3(G390), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1221), .A2(new_n1216), .A3(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1220), .A2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1178), .A2(new_n1186), .ZN(new_n1225));
  AND2_X1   g1025(.A1(new_n1225), .A2(new_n1157), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1178), .A2(new_n1206), .A3(new_n1180), .ZN(new_n1227));
  AOI21_X1  g1027(.A(G378), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(KEYINPUT124), .B1(new_n1182), .B2(G378), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1172), .B1(new_n1096), .B2(new_n1184), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1174), .B1(new_n1231), .B2(new_n1169), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1232), .A2(new_n673), .A3(new_n1181), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1170), .ZN(new_n1234));
  AND4_X1   g1034(.A1(KEYINPUT124), .A2(new_n1233), .A3(G378), .A4(new_n1234), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1229), .B1(new_n1230), .B2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT62), .ZN(new_n1237));
  INV_X1    g1037(.A(G343), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1238), .A2(G213), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1089), .B1(new_n1205), .B2(KEYINPUT60), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT125), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  OAI211_X1 g1042(.A(KEYINPUT125), .B(new_n1089), .C1(new_n1205), .C2(KEYINPUT60), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n674), .B1(new_n1205), .B2(KEYINPUT60), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1242), .A2(new_n1243), .A3(new_n1244), .ZN(new_n1245));
  AND3_X1   g1045(.A1(new_n1245), .A2(G384), .A3(new_n1204), .ZN(new_n1246));
  AOI21_X1  g1046(.A(G384), .B1(new_n1245), .B2(new_n1204), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1236), .A2(new_n1237), .A3(new_n1239), .A4(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1239), .ZN(new_n1250));
  OAI211_X1 g1050(.A(G2897), .B(new_n1250), .C1(new_n1246), .C2(new_n1247), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1247), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1245), .A2(G384), .A3(new_n1204), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1250), .A2(G2897), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1252), .A2(new_n1253), .A3(new_n1254), .ZN(new_n1255));
  AND2_X1   g1055(.A1(new_n1251), .A2(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1233), .A2(G378), .A3(new_n1234), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT124), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1233), .A2(G378), .A3(KEYINPUT124), .A4(new_n1234), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1228), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1256), .B1(new_n1261), .B2(new_n1250), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT61), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1249), .A2(new_n1262), .A3(new_n1263), .ZN(new_n1264));
  XNOR2_X1  g1064(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1250), .B1(new_n1266), .B2(new_n1229), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1265), .B1(new_n1267), .B2(new_n1248), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1224), .B1(new_n1264), .B2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1236), .A2(new_n1239), .ZN(new_n1270));
  AOI21_X1  g1070(.A(KEYINPUT61), .B1(new_n1270), .B2(new_n1256), .ZN(new_n1271));
  AND2_X1   g1071(.A1(new_n1220), .A2(new_n1223), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1236), .A2(new_n1239), .A3(new_n1248), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT63), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1267), .A2(KEYINPUT63), .A3(new_n1248), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1271), .A2(new_n1272), .A3(new_n1275), .A4(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1269), .A2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT127), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1269), .A2(new_n1277), .A3(KEYINPUT127), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(G405));
  OAI21_X1  g1082(.A(new_n1266), .B1(G378), .B2(new_n1182), .ZN(new_n1283));
  XNOR2_X1  g1083(.A(new_n1283), .B(new_n1248), .ZN(new_n1284));
  XNOR2_X1  g1084(.A(new_n1284), .B(new_n1224), .ZN(G402));
endmodule


