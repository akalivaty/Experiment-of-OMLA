//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 1 1 1 1 1 1 0 0 0 0 0 0 1 1 0 0 0 0 0 0 0 0 0 1 1 1 0 0 0 0 0 1 0 0 0 1 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:14 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n207, new_n208,
    new_n209, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XOR2_X1   g0003(.A(new_n203), .B(KEYINPUT64), .Z(new_n204));
  INV_X1    g0004(.A(G77), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(G353));
  INV_X1    g0006(.A(G97), .ZN(new_n207));
  INV_X1    g0007(.A(G107), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n209), .A2(G87), .ZN(G355));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n211), .A2(KEYINPUT65), .ZN(new_n212));
  INV_X1    g0012(.A(KEYINPUT65), .ZN(new_n213));
  NAND3_X1  g0013(.A1(new_n213), .A2(G1), .A3(G13), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G20), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT66), .ZN(new_n217));
  INV_X1    g0017(.A(KEYINPUT67), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n201), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(KEYINPUT67), .B1(G58), .B2(G68), .ZN(new_n220));
  NAND3_X1  g0020(.A1(new_n219), .A2(G50), .A3(new_n220), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n217), .A2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(G1), .ZN(new_n223));
  INV_X1    g0023(.A(G20), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n226), .A2(G13), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n227), .B(G250), .C1(G257), .C2(G264), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT0), .ZN(new_n229));
  XOR2_X1   g0029(.A(KEYINPUT68), .B(G244), .Z(new_n230));
  NOR2_X1   g0030(.A1(new_n230), .A2(new_n205), .ZN(new_n231));
  AOI22_X1  g0031(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n232));
  AOI22_X1  g0032(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n233));
  AOI22_X1  g0033(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n234));
  NAND2_X1  g0034(.A1(G107), .A2(G264), .ZN(new_n235));
  NAND4_X1  g0035(.A1(new_n232), .A2(new_n233), .A3(new_n234), .A4(new_n235), .ZN(new_n236));
  OAI21_X1  g0036(.A(new_n226), .B1(new_n231), .B2(new_n236), .ZN(new_n237));
  OAI21_X1  g0037(.A(new_n229), .B1(KEYINPUT1), .B2(new_n237), .ZN(new_n238));
  AOI211_X1 g0038(.A(new_n222), .B(new_n238), .C1(KEYINPUT1), .C2(new_n237), .ZN(G361));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  INV_X1    g0040(.A(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(KEYINPUT2), .B(G226), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G264), .B(G270), .Z(new_n245));
  XNOR2_X1  g0045(.A(G250), .B(G257), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G358));
  XNOR2_X1  g0048(.A(G50), .B(G68), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G58), .B(G77), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n249), .B(new_n250), .Z(new_n251));
  XOR2_X1   g0051(.A(G87), .B(G97), .Z(new_n252));
  XNOR2_X1  g0052(.A(G107), .B(G116), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n251), .B(new_n254), .ZN(G351));
  INV_X1    g0055(.A(G169), .ZN(new_n256));
  OR2_X1    g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G1698), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n259), .A2(G257), .A3(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G303), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n259), .A2(G1698), .ZN(new_n263));
  INV_X1    g0063(.A(G264), .ZN(new_n264));
  OAI221_X1 g0064(.A(new_n261), .B1(new_n262), .B2(new_n259), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(G33), .A2(G41), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n215), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g0069(.A(KEYINPUT5), .B(G41), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n266), .A2(G1), .A3(G13), .ZN(new_n271));
  INV_X1    g0071(.A(G45), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n272), .A2(G1), .ZN(new_n273));
  AND4_X1   g0073(.A1(G274), .A2(new_n270), .A3(new_n271), .A4(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n211), .B1(G33), .B2(G41), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n275), .B1(new_n273), .B2(new_n270), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n274), .B1(G270), .B2(new_n276), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n256), .B1(new_n269), .B2(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n223), .A2(G13), .A3(G20), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(KEYINPUT72), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT72), .ZN(new_n281));
  NAND4_X1  g0081(.A1(new_n281), .A2(new_n223), .A3(G13), .A4(G20), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n283), .A2(G116), .ZN(new_n284));
  AOI21_X1  g0084(.A(G20), .B1(G33), .B2(G283), .ZN(new_n285));
  INV_X1    g0085(.A(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G97), .ZN(new_n287));
  INV_X1    g0087(.A(G116), .ZN(new_n288));
  AOI22_X1  g0088(.A1(new_n285), .A2(new_n287), .B1(G20), .B2(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n212), .A2(new_n214), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT20), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n289), .A2(new_n291), .A3(KEYINPUT20), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n284), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT70), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n291), .A2(new_n297), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n212), .A2(new_n214), .A3(KEYINPUT70), .A4(new_n290), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n223), .A2(G33), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n300), .A2(G116), .A3(new_n283), .A4(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT85), .ZN(new_n303));
  AND3_X1   g0103(.A1(new_n296), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n303), .B1(new_n296), .B2(new_n302), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n278), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT21), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT86), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n309), .B1(new_n306), .B2(new_n307), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n296), .A2(new_n302), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(KEYINPUT85), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n296), .A2(new_n302), .A3(new_n303), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n269), .A2(new_n277), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n314), .A2(G179), .A3(new_n316), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n314), .A2(KEYINPUT86), .A3(KEYINPUT21), .A4(new_n278), .ZN(new_n318));
  AND4_X1   g0118(.A1(new_n308), .A2(new_n310), .A3(new_n317), .A4(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT71), .ZN(new_n320));
  INV_X1    g0120(.A(G58), .ZN(new_n321));
  NOR3_X1   g0121(.A1(new_n320), .A2(new_n321), .A3(KEYINPUT8), .ZN(new_n322));
  XNOR2_X1  g0122(.A(KEYINPUT8), .B(G58), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n322), .B1(new_n320), .B2(new_n323), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n286), .A2(G20), .ZN(new_n325));
  NOR2_X1   g0125(.A1(G20), .A2(G33), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n324), .A2(new_n325), .B1(G150), .B2(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n327), .B1(new_n224), .B2(new_n204), .ZN(new_n328));
  AND2_X1   g0128(.A1(new_n298), .A2(new_n299), .ZN(new_n329));
  AND2_X1   g0129(.A1(new_n280), .A2(new_n282), .ZN(new_n330));
  AOI22_X1  g0130(.A1(new_n328), .A2(new_n329), .B1(new_n202), .B2(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n330), .B1(new_n298), .B2(new_n299), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n223), .A2(G20), .ZN(new_n333));
  XNOR2_X1  g0133(.A(new_n333), .B(KEYINPUT73), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n332), .A2(G50), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n331), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(G1698), .B1(new_n257), .B2(new_n258), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(G222), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n259), .A2(G223), .A3(G1698), .ZN(new_n339));
  AND2_X1   g0139(.A1(KEYINPUT3), .A2(G33), .ZN(new_n340));
  NOR2_X1   g0140(.A1(KEYINPUT3), .A2(G33), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(G77), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n338), .A2(new_n339), .A3(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT69), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n338), .A2(new_n339), .A3(KEYINPUT69), .A4(new_n343), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n346), .A2(new_n268), .A3(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(G41), .ZN(new_n349));
  AOI21_X1  g0149(.A(G1), .B1(new_n349), .B2(new_n272), .ZN(new_n350));
  AND3_X1   g0150(.A1(new_n350), .A2(new_n271), .A3(G274), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n275), .A2(new_n350), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n351), .B1(G226), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n348), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(new_n256), .ZN(new_n355));
  OAI211_X1 g0155(.A(new_n336), .B(new_n355), .C1(G179), .C2(new_n354), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n337), .A2(G232), .B1(new_n342), .B2(G107), .ZN(new_n357));
  INV_X1    g0157(.A(G238), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n357), .B1(new_n358), .B2(new_n263), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n268), .ZN(new_n360));
  INV_X1    g0160(.A(new_n230), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n351), .B1(new_n361), .B2(new_n352), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(G190), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(new_n323), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n366), .A2(new_n326), .B1(G20), .B2(G77), .ZN(new_n367));
  XNOR2_X1  g0167(.A(KEYINPUT15), .B(G87), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n369), .A2(KEYINPUT74), .A3(new_n325), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n367), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(KEYINPUT74), .B1(new_n369), .B2(new_n325), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n329), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n332), .A2(G77), .A3(new_n334), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n373), .B(new_n374), .C1(G77), .C2(new_n283), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n365), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n363), .A2(G200), .ZN(new_n377));
  AND2_X1   g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n363), .A2(new_n256), .ZN(new_n379));
  INV_X1    g0179(.A(G179), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n360), .A2(new_n380), .A3(new_n362), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n379), .A2(new_n375), .A3(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n378), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT9), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n336), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n354), .A2(G200), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n331), .A2(KEYINPUT9), .A3(new_n335), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n348), .A2(G190), .A3(new_n353), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n386), .A2(new_n387), .A3(new_n388), .A4(new_n389), .ZN(new_n390));
  AND2_X1   g0190(.A1(new_n390), .A2(KEYINPUT10), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n390), .A2(KEYINPUT10), .ZN(new_n392));
  OAI211_X1 g0192(.A(new_n356), .B(new_n384), .C1(new_n391), .C2(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n351), .B1(G232), .B2(new_n352), .ZN(new_n394));
  INV_X1    g0194(.A(G226), .ZN(new_n395));
  INV_X1    g0195(.A(G87), .ZN(new_n396));
  OAI22_X1  g0196(.A1(new_n263), .A2(new_n395), .B1(new_n286), .B2(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(KEYINPUT81), .B1(new_n337), .B2(G223), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n337), .A2(KEYINPUT81), .A3(G223), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n397), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n364), .B(new_n394), .C1(new_n401), .C2(new_n267), .ZN(new_n402));
  INV_X1    g0202(.A(new_n394), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n342), .A2(new_n260), .ZN(new_n404));
  AOI22_X1  g0204(.A1(new_n404), .A2(G226), .B1(G33), .B2(G87), .ZN(new_n405));
  INV_X1    g0205(.A(new_n400), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n405), .B1(new_n406), .B2(new_n398), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n403), .B1(new_n407), .B2(new_n268), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n402), .B1(G200), .B2(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n257), .A2(new_n224), .A3(new_n258), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT7), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n257), .A2(KEYINPUT7), .A3(new_n224), .A4(new_n258), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(G68), .ZN(new_n415));
  INV_X1    g0215(.A(G68), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n321), .A2(new_n416), .ZN(new_n417));
  OR2_X1    g0217(.A1(new_n417), .A2(new_n201), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n418), .A2(G20), .B1(G159), .B2(new_n326), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n415), .A2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT16), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n415), .A2(KEYINPUT16), .A3(new_n419), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n422), .A2(new_n329), .A3(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n322), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n425), .B1(new_n366), .B2(KEYINPUT71), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n426), .B1(new_n300), .B2(new_n283), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n330), .B1(new_n334), .B2(new_n324), .ZN(new_n428));
  OAI21_X1  g0228(.A(KEYINPUT79), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT80), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n324), .A2(new_n334), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n283), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT79), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n432), .B(new_n433), .C1(new_n332), .C2(new_n426), .ZN(new_n434));
  AND3_X1   g0234(.A1(new_n429), .A2(new_n430), .A3(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n430), .B1(new_n429), .B2(new_n434), .ZN(new_n436));
  OAI211_X1 g0236(.A(new_n409), .B(new_n424), .C1(new_n435), .C2(new_n436), .ZN(new_n437));
  XNOR2_X1  g0237(.A(new_n437), .B(KEYINPUT17), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n408), .A2(new_n256), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n439), .B1(G179), .B2(new_n408), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n424), .B1(new_n435), .B2(new_n436), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(KEYINPUT18), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT18), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n442), .A2(new_n445), .A3(new_n441), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n438), .A2(new_n444), .A3(new_n446), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n393), .A2(new_n447), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n325), .A2(G77), .B1(G20), .B2(new_n416), .ZN(new_n449));
  INV_X1    g0249(.A(new_n326), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n449), .B1(new_n202), .B2(new_n450), .ZN(new_n451));
  AND2_X1   g0251(.A1(new_n329), .A2(new_n451), .ZN(new_n452));
  OR2_X1    g0252(.A1(new_n452), .A2(KEYINPUT11), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n330), .A2(new_n416), .ZN(new_n454));
  XNOR2_X1  g0254(.A(new_n454), .B(KEYINPUT12), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n452), .A2(KEYINPUT11), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n332), .A2(G68), .A3(new_n334), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n453), .A2(new_n455), .A3(new_n456), .A4(new_n457), .ZN(new_n458));
  AOI22_X1  g0258(.A1(new_n351), .A2(KEYINPUT75), .B1(new_n352), .B2(G238), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  NOR2_X1   g0260(.A1(G226), .A2(G1698), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n461), .B1(new_n241), .B2(G1698), .ZN(new_n462));
  AOI22_X1  g0262(.A1(new_n462), .A2(new_n259), .B1(G33), .B2(G97), .ZN(new_n463));
  OAI22_X1  g0263(.A1(new_n463), .A2(new_n267), .B1(new_n351), .B2(KEYINPUT75), .ZN(new_n464));
  OAI21_X1  g0264(.A(KEYINPUT13), .B1(new_n460), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n462), .A2(new_n259), .ZN(new_n466));
  NAND2_X1  g0266(.A1(G33), .A2(G97), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  AND2_X1   g0268(.A1(new_n271), .A2(G274), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(new_n350), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT75), .ZN(new_n471));
  AOI22_X1  g0271(.A1(new_n468), .A2(new_n268), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT13), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n472), .A2(new_n473), .A3(new_n459), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n256), .B1(new_n465), .B2(new_n474), .ZN(new_n475));
  XNOR2_X1  g0275(.A(new_n475), .B(KEYINPUT14), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT76), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n472), .A2(KEYINPUT76), .A3(new_n473), .A4(new_n459), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n478), .A2(G179), .A3(new_n465), .A4(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(KEYINPUT77), .B1(new_n476), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n465), .A2(new_n474), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(G169), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(KEYINPUT14), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT14), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n475), .A2(new_n485), .ZN(new_n486));
  AND4_X1   g0286(.A1(KEYINPUT77), .A2(new_n484), .A3(new_n480), .A4(new_n486), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n458), .B1(new_n481), .B2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n458), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n478), .A2(G190), .A3(new_n465), .A4(new_n479), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n482), .A2(G200), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n489), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n488), .A2(KEYINPUT78), .A3(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT78), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n476), .A2(KEYINPUT77), .A3(new_n480), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n484), .A2(new_n480), .A3(new_n486), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT77), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n489), .B1(new_n495), .B2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(new_n492), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n494), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  AND3_X1   g0301(.A1(new_n448), .A2(new_n493), .A3(new_n501), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n304), .A2(new_n305), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n315), .A2(G200), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n503), .B(new_n504), .C1(new_n364), .C2(new_n315), .ZN(new_n505));
  XNOR2_X1  g0305(.A(new_n505), .B(KEYINPUT87), .ZN(new_n506));
  AND3_X1   g0306(.A1(new_n208), .A2(KEYINPUT6), .A3(G97), .ZN(new_n507));
  XNOR2_X1  g0307(.A(G97), .B(G107), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT6), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  OAI22_X1  g0310(.A1(new_n510), .A2(new_n224), .B1(new_n205), .B2(new_n450), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n208), .B1(new_n412), .B2(new_n413), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n329), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n300), .A2(G97), .A3(new_n283), .A4(new_n301), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n283), .A2(G97), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  AND3_X1   g0316(.A1(new_n513), .A2(new_n514), .A3(new_n516), .ZN(new_n517));
  OAI211_X1 g0317(.A(G244), .B(new_n260), .C1(new_n340), .C2(new_n341), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT4), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n518), .A2(new_n519), .B1(G33), .B2(G283), .ZN(new_n520));
  OAI211_X1 g0320(.A(G250), .B(G1698), .C1(new_n340), .C2(new_n341), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT83), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n259), .A2(KEYINPUT83), .A3(G250), .A4(G1698), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n520), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT82), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n526), .B1(new_n518), .B2(new_n519), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n337), .A2(KEYINPUT82), .A3(KEYINPUT4), .A4(G244), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n268), .B1(new_n525), .B2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(new_n274), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n276), .A2(G257), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n530), .A2(G190), .A3(new_n534), .ZN(new_n535));
  AND2_X1   g0335(.A1(new_n523), .A2(new_n524), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n536), .A2(new_n520), .A3(new_n527), .A4(new_n528), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n533), .B1(new_n537), .B2(new_n268), .ZN(new_n538));
  INV_X1    g0338(.A(G200), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n517), .B(new_n535), .C1(new_n538), .C2(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n530), .A2(new_n380), .A3(new_n534), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n513), .A2(new_n514), .A3(new_n516), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n541), .B(new_n542), .C1(new_n538), .C2(G169), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n224), .B(G87), .C1(new_n340), .C2(new_n341), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(KEYINPUT22), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT22), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n259), .A2(new_n546), .A3(new_n224), .A4(G87), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT24), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n224), .A2(G33), .A3(G116), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT23), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n551), .A2(new_n208), .A3(G20), .ZN(new_n552));
  OAI21_X1  g0352(.A(KEYINPUT23), .B1(new_n224), .B2(G107), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT88), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n550), .B(new_n552), .C1(new_n553), .C2(new_n554), .ZN(new_n555));
  AND2_X1   g0355(.A1(new_n553), .A2(new_n554), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AND3_X1   g0357(.A1(new_n548), .A2(new_n549), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n549), .B1(new_n548), .B2(new_n557), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n329), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  OAI211_X1 g0360(.A(G257), .B(G1698), .C1(new_n340), .C2(new_n341), .ZN(new_n561));
  OAI211_X1 g0361(.A(G250), .B(new_n260), .C1(new_n340), .C2(new_n341), .ZN(new_n562));
  INV_X1    g0362(.A(G294), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n561), .B(new_n562), .C1(new_n286), .C2(new_n563), .ZN(new_n564));
  AOI22_X1  g0364(.A1(new_n564), .A2(new_n268), .B1(new_n276), .B2(G264), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n531), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(G200), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n300), .A2(G107), .A3(new_n283), .A4(new_n301), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n280), .A2(new_n208), .A3(new_n282), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT25), .ZN(new_n570));
  XNOR2_X1  g0370(.A(new_n569), .B(new_n570), .ZN(new_n571));
  AND2_X1   g0371(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n565), .A2(G190), .A3(new_n531), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n560), .A2(new_n567), .A3(new_n572), .A4(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n540), .A2(new_n543), .A3(new_n574), .ZN(new_n575));
  OAI211_X1 g0375(.A(G238), .B(new_n260), .C1(new_n340), .C2(new_n341), .ZN(new_n576));
  OAI211_X1 g0376(.A(G244), .B(G1698), .C1(new_n340), .C2(new_n341), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n576), .B(new_n577), .C1(new_n286), .C2(new_n288), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n268), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT84), .ZN(new_n580));
  INV_X1    g0380(.A(G250), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n273), .A2(new_n581), .ZN(new_n582));
  AOI22_X1  g0382(.A1(new_n469), .A2(new_n273), .B1(new_n271), .B2(new_n582), .ZN(new_n583));
  AND3_X1   g0383(.A1(new_n579), .A2(new_n580), .A3(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n580), .B1(new_n579), .B2(new_n583), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n256), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n579), .A2(new_n583), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(KEYINPUT84), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n579), .A2(new_n580), .A3(new_n583), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n588), .A2(new_n380), .A3(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n332), .A2(new_n301), .A3(new_n369), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT19), .ZN(new_n592));
  INV_X1    g0392(.A(new_n325), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n592), .B1(new_n593), .B2(new_n207), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n259), .A2(new_n224), .A3(G68), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n224), .B1(new_n467), .B2(new_n592), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n596), .B1(G87), .B2(new_n209), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n594), .A2(new_n595), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n329), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n330), .A2(new_n368), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n591), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n586), .A2(new_n590), .A3(new_n601), .ZN(new_n602));
  OAI21_X1  g0402(.A(G200), .B1(new_n584), .B2(new_n585), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n588), .A2(G190), .A3(new_n589), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n300), .A2(G87), .A3(new_n283), .A4(new_n301), .ZN(new_n605));
  AND3_X1   g0405(.A1(new_n599), .A2(new_n605), .A3(new_n600), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n603), .A2(new_n604), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n602), .A2(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(G169), .B1(new_n565), .B2(new_n531), .ZN(new_n609));
  INV_X1    g0409(.A(new_n566), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n609), .B1(new_n610), .B2(new_n380), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n560), .A2(new_n572), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  NOR3_X1   g0414(.A1(new_n575), .A2(new_n608), .A3(new_n614), .ZN(new_n615));
  AND4_X1   g0415(.A1(new_n319), .A2(new_n502), .A3(new_n506), .A4(new_n615), .ZN(G372));
  XNOR2_X1  g0416(.A(new_n390), .B(KEYINPUT10), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n488), .B1(new_n382), .B2(new_n500), .ZN(new_n618));
  AND2_X1   g0418(.A1(new_n618), .A2(new_n438), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n444), .A2(new_n446), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n617), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  AND2_X1   g0421(.A1(new_n621), .A2(new_n356), .ZN(new_n622));
  INV_X1    g0422(.A(new_n502), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n587), .A2(new_n256), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n590), .A2(new_n601), .A3(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n530), .A2(new_n534), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n450), .A2(new_n205), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n508), .A2(new_n509), .ZN(new_n629));
  INV_X1    g0429(.A(new_n507), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n628), .B1(new_n631), .B2(G20), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n414), .A2(G107), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n515), .B1(new_n634), .B2(new_n329), .ZN(new_n635));
  AOI22_X1  g0435(.A1(new_n256), .A2(new_n627), .B1(new_n635), .B2(new_n514), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n636), .A2(new_n602), .A3(new_n607), .A4(new_n541), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n626), .B1(new_n637), .B2(KEYINPUT26), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n587), .A2(G200), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n604), .A2(new_n606), .A3(new_n639), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n625), .A2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT89), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n636), .A2(new_n642), .A3(new_n541), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n543), .A2(KEYINPUT89), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n641), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n638), .B1(KEYINPUT26), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(KEYINPUT90), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT90), .ZN(new_n648));
  OAI211_X1 g0448(.A(new_n638), .B(new_n648), .C1(KEYINPUT26), .C2(new_n645), .ZN(new_n649));
  AOI22_X1  g0449(.A1(new_n306), .A2(new_n307), .B1(new_n611), .B2(new_n612), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n650), .A2(new_n310), .A3(new_n317), .A4(new_n318), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n625), .A2(new_n640), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n575), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n647), .A2(new_n649), .A3(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n622), .B1(new_n623), .B2(new_n656), .ZN(G369));
  NAND3_X1  g0457(.A1(new_n223), .A2(new_n224), .A3(G13), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n658), .A2(KEYINPUT27), .ZN(new_n659));
  XNOR2_X1  g0459(.A(new_n659), .B(KEYINPUT91), .ZN(new_n660));
  INV_X1    g0460(.A(G213), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n661), .B1(new_n658), .B2(KEYINPUT27), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(G343), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n314), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n506), .A2(new_n319), .A3(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n667), .B1(new_n319), .B2(new_n666), .ZN(new_n668));
  INV_X1    g0468(.A(new_n665), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n614), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n574), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n669), .B1(new_n560), .B2(new_n572), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n613), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n668), .A2(G330), .A3(new_n674), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n319), .A2(new_n665), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n674), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n675), .A2(new_n670), .A3(new_n677), .ZN(G399));
  NAND2_X1  g0478(.A1(new_n227), .A2(new_n349), .ZN(new_n679));
  NOR3_X1   g0479(.A1(new_n209), .A2(G87), .A3(G116), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n679), .A2(G1), .A3(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n681), .B1(new_n221), .B2(new_n679), .ZN(new_n682));
  XNOR2_X1  g0482(.A(new_n682), .B(KEYINPUT28), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT29), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n684), .B1(new_n656), .B2(new_n665), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n608), .A2(new_n543), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT26), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n626), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n645), .A2(KEYINPUT26), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT93), .ZN(new_n691));
  AND3_X1   g0491(.A1(new_n651), .A2(new_n653), .A3(new_n691), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n691), .B1(new_n651), .B2(new_n653), .ZN(new_n693));
  NOR3_X1   g0493(.A1(new_n690), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(KEYINPUT94), .B1(new_n694), .B2(new_n665), .ZN(new_n695));
  INV_X1    g0495(.A(new_n693), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n651), .A2(new_n653), .A3(new_n691), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n696), .A2(new_n697), .A3(new_n689), .A4(new_n688), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT94), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n698), .A2(new_n699), .A3(new_n669), .ZN(new_n700));
  AND2_X1   g0500(.A1(new_n695), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n685), .B1(new_n701), .B2(new_n684), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n506), .A2(new_n319), .A3(new_n615), .A4(new_n669), .ZN(new_n703));
  AND4_X1   g0503(.A1(G179), .A2(new_n269), .A3(new_n277), .A4(new_n565), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n584), .A2(new_n585), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n704), .A2(new_n538), .A3(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT30), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n316), .A2(G179), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n709), .A2(new_n627), .A3(new_n566), .A4(new_n587), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n704), .A2(KEYINPUT30), .A3(new_n705), .A4(new_n538), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n708), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n712), .A2(KEYINPUT31), .A3(new_n665), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(KEYINPUT92), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n712), .A2(new_n665), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT31), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT92), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n712), .A2(new_n718), .A3(KEYINPUT31), .A4(new_n665), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n703), .A2(new_n714), .A3(new_n717), .A4(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(G330), .ZN(new_n721));
  AND2_X1   g0521(.A1(new_n702), .A2(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n683), .B1(new_n722), .B2(G1), .ZN(G364));
  INV_X1    g0523(.A(new_n679), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n224), .A2(G13), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n223), .B1(new_n726), .B2(G45), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n724), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n227), .A2(new_n259), .ZN(new_n730));
  INV_X1    g0530(.A(G355), .ZN(new_n731));
  OAI22_X1  g0531(.A1(new_n730), .A2(new_n731), .B1(G116), .B2(new_n227), .ZN(new_n732));
  OR2_X1    g0532(.A1(new_n251), .A2(new_n272), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n227), .A2(new_n342), .ZN(new_n734));
  INV_X1    g0534(.A(new_n221), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n734), .B1(new_n735), .B2(new_n272), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n732), .B1(new_n733), .B2(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n215), .B1(new_n224), .B2(G169), .ZN(new_n738));
  NOR2_X1   g0538(.A1(G13), .A2(G33), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(G20), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n738), .A2(new_n742), .ZN(new_n743));
  XOR2_X1   g0543(.A(new_n743), .B(KEYINPUT95), .Z(new_n744));
  OAI21_X1  g0544(.A(new_n729), .B1(new_n737), .B2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n224), .A2(new_n380), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n746), .A2(G190), .A3(new_n539), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n224), .A2(G179), .ZN(new_n748));
  NOR2_X1   g0548(.A1(G190), .A2(G200), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(G159), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT32), .ZN(new_n753));
  OAI221_X1 g0553(.A(new_n259), .B1(new_n321), .B2(new_n747), .C1(new_n752), .C2(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n754), .B1(new_n753), .B2(new_n752), .ZN(new_n755));
  NOR3_X1   g0555(.A1(new_n364), .A2(G179), .A3(G200), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(new_n224), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n539), .A2(G190), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n746), .A2(new_n758), .ZN(new_n759));
  OAI22_X1  g0559(.A1(new_n757), .A2(new_n207), .B1(new_n759), .B2(new_n416), .ZN(new_n760));
  XNOR2_X1  g0560(.A(new_n760), .B(KEYINPUT96), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n364), .A2(new_n539), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(new_n748), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n748), .A2(new_n758), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AOI22_X1  g0566(.A1(G87), .A2(new_n764), .B1(new_n766), .B2(G107), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n746), .A2(new_n762), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n746), .A2(new_n749), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  AOI22_X1  g0571(.A1(G50), .A2(new_n769), .B1(new_n771), .B2(G77), .ZN(new_n772));
  NAND4_X1  g0572(.A1(new_n755), .A2(new_n761), .A3(new_n767), .A4(new_n772), .ZN(new_n773));
  XNOR2_X1  g0573(.A(new_n768), .B(KEYINPUT97), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  XNOR2_X1  g0575(.A(KEYINPUT98), .B(G326), .ZN(new_n776));
  INV_X1    g0576(.A(new_n757), .ZN(new_n777));
  AOI22_X1  g0577(.A1(new_n775), .A2(new_n776), .B1(G294), .B2(new_n777), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n778), .B(KEYINPUT99), .ZN(new_n779));
  INV_X1    g0579(.A(new_n759), .ZN(new_n780));
  INV_X1    g0580(.A(G317), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(KEYINPUT33), .ZN(new_n782));
  OR2_X1    g0582(.A1(new_n781), .A2(KEYINPUT33), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n780), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n784), .B1(new_n262), .B2(new_n763), .ZN(new_n785));
  INV_X1    g0585(.A(new_n750), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n785), .B1(G329), .B2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n747), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n259), .B1(new_n788), .B2(G322), .ZN(new_n789));
  AOI22_X1  g0589(.A1(G311), .A2(new_n771), .B1(new_n766), .B2(G283), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n787), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n773), .B1(new_n779), .B2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n738), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n745), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n794), .B1(new_n668), .B2(new_n742), .ZN(new_n795));
  XOR2_X1   g0595(.A(new_n795), .B(KEYINPUT100), .Z(new_n796));
  AOI21_X1  g0596(.A(new_n729), .B1(new_n668), .B2(G330), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n797), .B1(G330), .B2(new_n668), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  XOR2_X1   g0599(.A(new_n799), .B(KEYINPUT101), .Z(G396));
  NAND2_X1  g0600(.A1(new_n655), .A2(new_n669), .ZN(new_n801));
  AND2_X1   g0601(.A1(new_n375), .A2(new_n665), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n382), .B1(new_n378), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n383), .A2(new_n669), .ZN(new_n804));
  AND2_X1   g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  XOR2_X1   g0605(.A(new_n801), .B(new_n805), .Z(new_n806));
  AOI21_X1  g0606(.A(new_n729), .B1(new_n806), .B2(new_n721), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n807), .B1(new_n721), .B2(new_n806), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n738), .A2(new_n740), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n729), .B1(new_n809), .B2(G77), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n788), .A2(G143), .B1(new_n771), .B2(G159), .ZN(new_n811));
  INV_X1    g0611(.A(G137), .ZN(new_n812));
  INV_X1    g0612(.A(G150), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n811), .B1(new_n812), .B2(new_n768), .C1(new_n813), .C2(new_n759), .ZN(new_n814));
  INV_X1    g0614(.A(KEYINPUT34), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(G132), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n259), .B1(new_n750), .B2(new_n817), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n763), .A2(new_n202), .B1(new_n765), .B2(new_n416), .ZN(new_n819));
  AOI211_X1 g0619(.A(new_n818), .B(new_n819), .C1(G58), .C2(new_n777), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n816), .A2(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n814), .A2(new_n815), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  AOI22_X1  g0623(.A1(G283), .A2(new_n780), .B1(new_n766), .B2(G87), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n259), .B1(new_n771), .B2(G116), .ZN(new_n825));
  OAI211_X1 g0625(.A(new_n824), .B(new_n825), .C1(new_n207), .C2(new_n757), .ZN(new_n826));
  INV_X1    g0626(.A(G311), .ZN(new_n827));
  OAI22_X1  g0627(.A1(new_n763), .A2(new_n208), .B1(new_n750), .B2(new_n827), .ZN(new_n828));
  OAI22_X1  g0628(.A1(new_n747), .A2(new_n563), .B1(new_n768), .B2(new_n262), .ZN(new_n829));
  NOR3_X1   g0629(.A1(new_n826), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n823), .B1(KEYINPUT102), .B2(new_n831), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n832), .B1(KEYINPUT102), .B2(new_n831), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n810), .B1(new_n833), .B2(new_n793), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n834), .B1(new_n805), .B2(new_n740), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n808), .A2(new_n835), .ZN(G384));
  INV_X1    g0636(.A(KEYINPUT39), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT37), .ZN(new_n838));
  INV_X1    g0638(.A(new_n424), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n429), .A2(new_n434), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(KEYINPUT80), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n429), .A2(new_n434), .A3(new_n430), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n839), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n437), .B(new_n838), .C1(new_n843), .C2(new_n440), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT104), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n846), .B1(new_n843), .B2(new_n663), .ZN(new_n847));
  INV_X1    g0647(.A(new_n663), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n442), .A2(KEYINPUT104), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  AND3_X1   g0650(.A1(new_n845), .A2(new_n850), .A3(KEYINPUT105), .ZN(new_n851));
  AOI21_X1  g0651(.A(KEYINPUT105), .B1(new_n845), .B2(new_n850), .ZN(new_n852));
  OAI21_X1  g0652(.A(KEYINPUT106), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT105), .ZN(new_n854));
  AND3_X1   g0654(.A1(new_n442), .A2(KEYINPUT104), .A3(new_n848), .ZN(new_n855));
  AOI21_X1  g0655(.A(KEYINPUT104), .B1(new_n442), .B2(new_n848), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n854), .B1(new_n857), .B2(new_n844), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n845), .A2(new_n850), .A3(KEYINPUT105), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT106), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n443), .A2(new_n437), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n838), .B1(new_n863), .B2(new_n850), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n853), .A2(new_n861), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n447), .A2(new_n857), .ZN(new_n867));
  AOI21_X1  g0667(.A(KEYINPUT38), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n423), .A2(new_n329), .ZN(new_n869));
  OR2_X1    g0669(.A1(new_n420), .A2(KEYINPUT103), .ZN(new_n870));
  AOI21_X1  g0670(.A(KEYINPUT16), .B1(new_n420), .B2(KEYINPUT103), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n869), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  OR2_X1    g0672(.A1(new_n872), .A2(new_n840), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n873), .B1(new_n441), .B2(new_n848), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n838), .B1(new_n874), .B2(new_n437), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n875), .B1(new_n858), .B2(new_n859), .ZN(new_n876));
  AND2_X1   g0676(.A1(new_n873), .A2(new_n848), .ZN(new_n877));
  AND2_X1   g0677(.A1(new_n447), .A2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT38), .ZN(new_n879));
  NOR3_X1   g0679(.A1(new_n876), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n837), .B1(new_n868), .B2(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n488), .A2(new_n665), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n879), .B1(new_n876), .B2(new_n878), .ZN(new_n883));
  INV_X1    g0683(.A(new_n875), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n884), .B1(new_n851), .B2(new_n852), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n447), .A2(new_n877), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n885), .A2(KEYINPUT38), .A3(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n883), .A2(new_n887), .A3(KEYINPUT39), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n881), .A2(new_n882), .A3(new_n888), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n489), .A2(new_n669), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n890), .B1(new_n499), .B2(new_n500), .ZN(new_n891));
  INV_X1    g0691(.A(new_n890), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n488), .A2(new_n492), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n655), .A2(new_n669), .A3(new_n805), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n895), .B1(new_n896), .B2(new_n804), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n883), .A2(new_n887), .ZN(new_n898));
  AOI22_X1  g0698(.A1(new_n897), .A2(new_n898), .B1(new_n620), .B2(new_n663), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n889), .A2(new_n899), .ZN(new_n900));
  OAI211_X1 g0700(.A(new_n502), .B(new_n685), .C1(new_n701), .C2(new_n684), .ZN(new_n901));
  AND2_X1   g0701(.A1(new_n901), .A2(new_n622), .ZN(new_n902));
  XOR2_X1   g0702(.A(new_n900), .B(new_n902), .Z(new_n903));
  INV_X1    g0703(.A(G330), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT107), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n703), .A2(new_n713), .A3(new_n717), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n894), .A2(new_n805), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n907), .B1(new_n883), .B2(new_n887), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n905), .B1(new_n908), .B2(KEYINPUT40), .ZN(new_n909));
  AND3_X1   g0709(.A1(new_n894), .A2(new_n805), .A3(new_n906), .ZN(new_n910));
  AOI21_X1  g0710(.A(KEYINPUT38), .B1(new_n885), .B2(new_n886), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n910), .B1(new_n880), .B2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT40), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n912), .A2(KEYINPUT107), .A3(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n867), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n858), .A2(new_n859), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n864), .B1(new_n916), .B2(KEYINPUT106), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n915), .B1(new_n917), .B2(new_n861), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n887), .B1(new_n918), .B2(KEYINPUT38), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n907), .A2(new_n913), .ZN(new_n920));
  AOI22_X1  g0720(.A1(new_n909), .A2(new_n914), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n448), .A2(new_n906), .A3(new_n493), .A4(new_n501), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n904), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n924), .B1(new_n921), .B2(new_n923), .ZN(new_n925));
  AOI22_X1  g0725(.A1(new_n903), .A2(new_n925), .B1(G1), .B2(new_n725), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n903), .B2(new_n925), .ZN(new_n927));
  OAI21_X1  g0727(.A(G116), .B1(new_n631), .B2(KEYINPUT35), .ZN(new_n928));
  AOI211_X1 g0728(.A(new_n928), .B(new_n217), .C1(KEYINPUT35), .C2(new_n631), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n929), .B(KEYINPUT36), .ZN(new_n930));
  OR3_X1    g0730(.A1(new_n221), .A2(new_n205), .A3(new_n417), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n202), .A2(G68), .ZN(new_n932));
  AOI211_X1 g0732(.A(new_n223), .B(G13), .C1(new_n931), .C2(new_n932), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n930), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n927), .A2(new_n934), .ZN(G367));
  OAI22_X1  g0735(.A1(new_n247), .A2(new_n734), .B1(new_n227), .B2(new_n368), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n729), .B1(new_n744), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n775), .A2(G143), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n765), .A2(new_n205), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n259), .B1(new_n763), .B2(new_n321), .ZN(new_n940));
  AOI211_X1 g0740(.A(new_n939), .B(new_n940), .C1(G137), .C2(new_n786), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n777), .A2(G68), .ZN(new_n942));
  OAI22_X1  g0742(.A1(new_n747), .A2(new_n813), .B1(new_n759), .B2(new_n751), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n943), .B1(G50), .B2(new_n771), .ZN(new_n944));
  NAND4_X1  g0744(.A1(new_n938), .A2(new_n941), .A3(new_n942), .A4(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT111), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n763), .B2(new_n288), .ZN(new_n947));
  AOI22_X1  g0747(.A1(new_n775), .A2(G311), .B1(KEYINPUT46), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n342), .B1(new_n759), .B2(new_n563), .ZN(new_n949));
  OAI22_X1  g0749(.A1(new_n765), .A2(new_n207), .B1(new_n750), .B2(new_n781), .ZN(new_n950));
  AOI211_X1 g0750(.A(new_n949), .B(new_n950), .C1(G303), .C2(new_n788), .ZN(new_n951));
  OAI211_X1 g0751(.A(new_n948), .B(new_n951), .C1(KEYINPUT46), .C2(new_n947), .ZN(new_n952));
  INV_X1    g0752(.A(G283), .ZN(new_n953));
  OAI22_X1  g0753(.A1(new_n757), .A2(new_n208), .B1(new_n770), .B2(new_n953), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n954), .B(KEYINPUT110), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n945), .B1(new_n952), .B2(new_n955), .ZN(new_n956));
  XOR2_X1   g0756(.A(new_n956), .B(KEYINPUT47), .Z(new_n957));
  NOR2_X1   g0757(.A1(new_n957), .A2(new_n738), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n669), .A2(new_n606), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n625), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(new_n641), .B2(new_n959), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT108), .ZN(new_n962));
  AOI211_X1 g0762(.A(new_n937), .B(new_n958), .C1(new_n741), .C2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n677), .A2(new_n670), .ZN(new_n965));
  OAI211_X1 g0765(.A(new_n540), .B(new_n543), .C1(new_n517), .C2(new_n669), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n636), .A2(new_n541), .A3(new_n665), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n965), .A2(new_n969), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n970), .B(KEYINPUT44), .Z(new_n971));
  NOR2_X1   g0771(.A1(new_n965), .A2(new_n969), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT45), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(new_n675), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n668), .A2(G330), .ZN(new_n977));
  INV_X1    g0777(.A(new_n674), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n676), .B(new_n978), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n977), .B(new_n979), .Z(new_n980));
  OAI21_X1  g0780(.A(new_n722), .B1(new_n976), .B2(new_n980), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n679), .B(KEYINPUT41), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n728), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n676), .A2(new_n674), .A3(new_n968), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(KEYINPUT42), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n543), .B1(new_n966), .B2(new_n613), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT109), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n987), .A2(new_n988), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n989), .A2(new_n669), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n986), .A2(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n985), .A2(KEYINPUT42), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT43), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n992), .A2(new_n993), .B1(new_n994), .B2(new_n962), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n962), .A2(new_n994), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n995), .B(new_n996), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n675), .A2(new_n969), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n997), .B(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n964), .B1(new_n984), .B2(new_n999), .ZN(G387));
  OAI22_X1  g0800(.A1(new_n730), .A2(new_n680), .B1(G107), .B2(new_n227), .ZN(new_n1001));
  AND2_X1   g0801(.A1(new_n680), .A2(KEYINPUT112), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n680), .A2(KEYINPUT112), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n272), .B1(new_n416), .B2(new_n205), .ZN(new_n1004));
  NOR3_X1   g0804(.A1(new_n1002), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n1005), .A2(KEYINPUT113), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(KEYINPUT113), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n323), .A2(G50), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT50), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1006), .A2(new_n1007), .A3(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n734), .B1(new_n244), .B2(G45), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1001), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(G159), .A2(new_n769), .B1(new_n764), .B2(G77), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n1013), .B1(new_n416), .B2(new_n770), .C1(new_n426), .C2(new_n759), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n757), .A2(new_n368), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n259), .B1(new_n765), .B2(new_n207), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n747), .A2(new_n202), .B1(new_n750), .B2(new_n813), .ZN(new_n1017));
  NOR4_X1   g0817(.A1(new_n1014), .A2(new_n1015), .A3(new_n1016), .A4(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n342), .B1(new_n765), .B2(new_n288), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n788), .A2(G317), .B1(new_n780), .B2(G311), .ZN(new_n1020));
  INV_X1    g0820(.A(G322), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n1020), .B1(new_n262), .B2(new_n770), .C1(new_n774), .C2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT48), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n777), .A2(G283), .B1(new_n764), .B2(G294), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT49), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  AOI211_X1 g0829(.A(new_n1019), .B(new_n1029), .C1(new_n776), .C2(new_n786), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1018), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n729), .B1(new_n744), .B2(new_n1012), .C1(new_n1032), .C2(new_n738), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1033), .B1(new_n978), .B2(new_n741), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n980), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1034), .B1(new_n1035), .B2(new_n728), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n722), .A2(new_n1035), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(new_n724), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n722), .A2(new_n1035), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1036), .B1(new_n1038), .B2(new_n1039), .ZN(G393));
  OAI22_X1  g0840(.A1(new_n254), .A2(new_n734), .B1(new_n207), .B2(new_n227), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n729), .B1(new_n744), .B2(new_n1041), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n757), .A2(new_n205), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n342), .B(new_n1043), .C1(G87), .C2(new_n766), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n747), .A2(new_n751), .B1(new_n768), .B2(new_n813), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT51), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n366), .A2(new_n771), .B1(new_n764), .B2(G68), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(G50), .A2(new_n780), .B1(new_n786), .B2(G143), .ZN(new_n1048));
  NAND4_X1  g0848(.A1(new_n1044), .A2(new_n1046), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(G283), .A2(new_n764), .B1(new_n786), .B2(G322), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n1050), .B(new_n342), .C1(new_n208), .C2(new_n765), .ZN(new_n1051));
  XOR2_X1   g0851(.A(new_n1051), .B(KEYINPUT115), .Z(new_n1052));
  OAI22_X1  g0852(.A1(new_n747), .A2(new_n827), .B1(new_n768), .B2(new_n781), .ZN(new_n1053));
  XOR2_X1   g0853(.A(KEYINPUT114), .B(KEYINPUT52), .Z(new_n1054));
  INV_X1    g0854(.A(new_n1054), .ZN(new_n1055));
  OR2_X1    g0855(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n777), .A2(G116), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(G294), .A2(new_n771), .B1(new_n780), .B2(G303), .ZN(new_n1059));
  NAND4_X1  g0859(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .A4(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1049), .B1(new_n1052), .B2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1042), .B1(new_n1061), .B2(new_n793), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1062), .B1(new_n968), .B2(new_n742), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n724), .B1(new_n976), .B2(new_n1037), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n975), .B1(new_n722), .B2(new_n1035), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1063), .B1(new_n727), .B2(new_n976), .C1(new_n1064), .C2(new_n1065), .ZN(G390));
  AND2_X1   g0866(.A1(new_n805), .A2(G330), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n894), .A2(new_n906), .A3(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1068), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n897), .A2(new_n882), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(new_n881), .B2(new_n888), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n882), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1072), .B1(new_n868), .B2(new_n880), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n695), .A2(new_n700), .A3(new_n804), .ZN(new_n1074));
  AND3_X1   g0874(.A1(new_n1074), .A2(new_n803), .A3(new_n894), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1069), .B1(new_n1071), .B2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1074), .A2(new_n803), .A3(new_n894), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n919), .A2(new_n1072), .A3(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n720), .A2(new_n1067), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n895), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n888), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(new_n919), .B2(new_n837), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n1079), .B(new_n1082), .C1(new_n1084), .C2(new_n1070), .ZN(new_n1085));
  OR3_X1    g0885(.A1(new_n922), .A2(KEYINPUT116), .A3(new_n904), .ZN(new_n1086));
  OAI21_X1  g0886(.A(KEYINPUT116), .B1(new_n922), .B2(new_n904), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n901), .A2(new_n1088), .A3(new_n622), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n895), .A2(new_n1080), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n1090), .A2(new_n1068), .B1(new_n896), .B2(new_n804), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n894), .B1(new_n906), .B2(new_n1067), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n1081), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1074), .A2(new_n803), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1091), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n1089), .A2(new_n1095), .ZN(new_n1096));
  AND3_X1   g0896(.A1(new_n1077), .A2(new_n1085), .A3(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1096), .B1(new_n1077), .B2(new_n1085), .ZN(new_n1098));
  NOR3_X1   g0898(.A1(new_n1097), .A2(new_n1098), .A3(new_n679), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1077), .A2(new_n1085), .A3(new_n728), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n729), .B1(new_n809), .B2(new_n324), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n342), .B1(new_n763), .B2(new_n396), .ZN(new_n1102));
  XOR2_X1   g0902(.A(new_n1102), .B(KEYINPUT120), .Z(new_n1103));
  AOI22_X1  g0903(.A1(new_n788), .A2(G116), .B1(new_n771), .B2(G97), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n769), .A2(G283), .B1(new_n786), .B2(G294), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n759), .A2(new_n208), .B1(new_n765), .B2(new_n416), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1106), .A2(new_n1043), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n1103), .A2(new_n1104), .A3(new_n1105), .A4(new_n1107), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n763), .A2(new_n813), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(new_n1109), .B(KEYINPUT119), .ZN(new_n1110));
  XOR2_X1   g0910(.A(KEYINPUT118), .B(KEYINPUT53), .Z(new_n1111));
  OR2_X1    g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n259), .B1(new_n747), .B2(new_n817), .ZN(new_n1113));
  INV_X1    g0913(.A(G128), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n768), .A2(new_n1114), .B1(new_n765), .B2(new_n202), .ZN(new_n1115));
  AOI211_X1 g0915(.A(new_n1113), .B(new_n1115), .C1(G125), .C2(new_n786), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1112), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(KEYINPUT54), .B(G143), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n812), .A2(new_n759), .B1(new_n770), .B2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1120), .B1(G159), .B2(new_n777), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(new_n1121), .B(KEYINPUT117), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1108), .B1(new_n1118), .B2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1101), .B1(new_n1123), .B2(new_n793), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n1084), .B2(new_n740), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1100), .A2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g0926(.A(KEYINPUT121), .B1(new_n1099), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1077), .A2(new_n1085), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1096), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1077), .A2(new_n1085), .A3(new_n1096), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1130), .A2(new_n724), .A3(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT121), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n1132), .A2(new_n1133), .A3(new_n1100), .A4(new_n1125), .ZN(new_n1134));
  AND2_X1   g0934(.A1(new_n1127), .A2(new_n1134), .ZN(G378));
  INV_X1    g0935(.A(KEYINPUT123), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n617), .A2(new_n356), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n336), .A2(new_n848), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1137), .B(new_n1138), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1136), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1143), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1145), .A2(KEYINPUT123), .A3(new_n1141), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1144), .A2(new_n1146), .A3(new_n739), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n729), .B1(new_n809), .B2(G50), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n747), .A2(new_n1114), .B1(new_n759), .B2(new_n817), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(G125), .A2(new_n769), .B1(new_n771), .B2(G137), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1150), .B1(new_n763), .B2(new_n1119), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n1149), .B(new_n1151), .C1(G150), .C2(new_n777), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT59), .ZN(new_n1153));
  OR2_X1    g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(G33), .A2(G41), .ZN(new_n1156));
  XOR2_X1   g0956(.A(new_n1156), .B(KEYINPUT122), .Z(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(G159), .A2(new_n766), .B1(new_n786), .B2(G124), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1154), .A2(new_n1155), .A3(new_n1158), .A4(new_n1159), .ZN(new_n1160));
  AOI211_X1 g0960(.A(G41), .B(new_n259), .C1(new_n764), .C2(G77), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n369), .A2(new_n771), .B1(new_n786), .B2(G283), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n1161), .B(new_n1162), .C1(new_n416), .C2(new_n757), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n747), .A2(new_n208), .B1(new_n765), .B2(new_n321), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n768), .A2(new_n288), .B1(new_n759), .B2(new_n207), .ZN(new_n1165));
  NOR3_X1   g0965(.A1(new_n1163), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(KEYINPUT58), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1157), .B(new_n202), .C1(G41), .C2(new_n259), .ZN(new_n1168));
  OR2_X1    g0968(.A1(new_n1166), .A2(KEYINPUT58), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n1160), .A2(new_n1167), .A3(new_n1168), .A4(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1148), .B1(new_n1170), .B2(new_n793), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1147), .A2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n900), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n909), .A2(new_n914), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n904), .B1(new_n919), .B2(new_n920), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1176));
  AND3_X1   g0976(.A1(new_n1174), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1145), .A2(new_n1141), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1173), .B1(new_n1177), .B2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1174), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n866), .A2(new_n867), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n880), .B1(new_n1182), .B2(new_n879), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n920), .ZN(new_n1184));
  OAI21_X1  g0984(.A(G330), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(new_n909), .B2(new_n914), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1181), .B(new_n900), .C1(new_n1186), .C2(new_n1178), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1180), .A2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1172), .B1(new_n1188), .B2(new_n727), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  AND2_X1   g0990(.A1(new_n1180), .A2(new_n1187), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1089), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1131), .A2(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(KEYINPUT57), .B1(new_n1191), .B2(new_n1193), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1180), .A2(new_n1187), .A3(KEYINPUT57), .ZN(new_n1195));
  AND2_X1   g0995(.A1(new_n1131), .A2(new_n1192), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n724), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1190), .B1(new_n1194), .B2(new_n1197), .ZN(G375));
  OR2_X1    g0998(.A1(new_n1095), .A2(new_n727), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT124), .ZN(new_n1200));
  OR2_X1    g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n729), .B1(new_n809), .B2(G68), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n768), .A2(new_n817), .B1(new_n750), .B2(new_n1114), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n342), .B(new_n1203), .C1(G58), .C2(new_n766), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n813), .A2(new_n770), .B1(new_n759), .B2(new_n1119), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n747), .A2(new_n812), .B1(new_n763), .B2(new_n751), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1204), .B(new_n1207), .C1(new_n202), .C2(new_n757), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n768), .A2(new_n563), .B1(new_n759), .B2(new_n288), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(G107), .B2(new_n771), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(new_n1210), .B(KEYINPUT125), .ZN(new_n1211));
  NOR3_X1   g1011(.A1(new_n1015), .A2(new_n259), .A3(new_n939), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n788), .A2(G283), .B1(new_n764), .B2(G97), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n1212), .B(new_n1213), .C1(new_n262), .C2(new_n750), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1208), .B1(new_n1211), .B2(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1202), .B1(new_n1215), .B2(new_n793), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1216), .B1(new_n894), .B2(new_n740), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1201), .A2(new_n1217), .A3(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1089), .A2(new_n1095), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1096), .A2(new_n982), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1219), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(new_n1222), .B(KEYINPUT126), .ZN(G381));
  NOR2_X1   g1023(.A1(new_n1099), .A2(new_n1126), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  NOR4_X1   g1025(.A1(G390), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n1226), .B(new_n964), .C1(new_n984), .C2(new_n999), .ZN(new_n1227));
  OR4_X1    g1027(.A1(new_n1225), .A2(new_n1227), .A3(G381), .A4(G375), .ZN(G407));
  AND3_X1   g1028(.A1(new_n1180), .A2(new_n1187), .A3(KEYINPUT57), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n679), .B1(new_n1229), .B2(new_n1193), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT57), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1231), .B1(new_n1196), .B2(new_n1188), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1189), .B1(new_n1230), .B2(new_n1232), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n661), .A2(G343), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1233), .A2(new_n1224), .A3(new_n1234), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(G407), .A2(G213), .A3(new_n1235), .ZN(G409));
  NOR3_X1   g1036(.A1(new_n1196), .A2(new_n1188), .A3(new_n982), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1224), .B1(new_n1237), .B2(new_n1189), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1127), .A2(new_n1134), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1238), .B1(G375), .B2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1234), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1089), .A2(KEYINPUT60), .A3(new_n1095), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(new_n724), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1129), .A2(KEYINPUT60), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1243), .B1(new_n1244), .B2(new_n1220), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1245), .A2(new_n1219), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(G384), .ZN(new_n1247));
  OAI211_X1 g1047(.A(new_n835), .B(new_n808), .C1(new_n1245), .C2(new_n1219), .ZN(new_n1248));
  AND2_X1   g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1240), .A2(new_n1241), .A3(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(KEYINPUT62), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT61), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1234), .A2(G2897), .ZN(new_n1253));
  AND3_X1   g1053(.A1(new_n1247), .A2(new_n1248), .A3(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1253), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1191), .A2(new_n983), .A3(new_n1193), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1190), .A2(new_n1257), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(G378), .A2(new_n1233), .B1(new_n1258), .B2(new_n1224), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1256), .B1(new_n1259), .B2(new_n1234), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT62), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1240), .A2(new_n1261), .A3(new_n1241), .A4(new_n1249), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1251), .A2(new_n1252), .A3(new_n1260), .A4(new_n1262), .ZN(new_n1263));
  XNOR2_X1  g1063(.A(G387), .B(G390), .ZN(new_n1264));
  XNOR2_X1  g1064(.A(G393), .B(G396), .ZN(new_n1265));
  XNOR2_X1  g1065(.A(new_n1264), .B(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1263), .A2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1269));
  AOI21_X1  g1069(.A(KEYINPUT61), .B1(new_n1269), .B2(new_n1256), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT63), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1250), .A2(new_n1271), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1240), .A2(KEYINPUT63), .A3(new_n1241), .A4(new_n1249), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1266), .A2(new_n1270), .A3(new_n1272), .A4(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1268), .A2(new_n1274), .ZN(G405));
  NOR2_X1   g1075(.A1(new_n1233), .A2(new_n1225), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(G375), .A2(new_n1239), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1278), .A2(KEYINPUT127), .A3(new_n1249), .ZN(new_n1279));
  OR2_X1    g1079(.A1(new_n1249), .A2(KEYINPUT127), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1249), .A2(KEYINPUT127), .ZN(new_n1281));
  OAI211_X1 g1081(.A(new_n1280), .B(new_n1281), .C1(new_n1277), .C2(new_n1276), .ZN(new_n1282));
  AND3_X1   g1082(.A1(new_n1266), .A2(new_n1279), .A3(new_n1282), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1266), .B1(new_n1282), .B2(new_n1279), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1283), .A2(new_n1284), .ZN(G402));
endmodule


