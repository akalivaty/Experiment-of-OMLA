//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 1 0 0 0 1 0 1 1 0 0 0 0 0 1 1 0 0 0 1 1 1 0 1 0 0 0 0 0 1 0 0 1 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 0 1 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n737, new_n738, new_n739, new_n741, new_n742, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n855, new_n856,
    new_n858, new_n859, new_n860, new_n861, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1010, new_n1011;
  INV_X1    g000(.A(KEYINPUT83), .ZN(new_n202));
  XNOR2_X1  g001(.A(G15gat), .B(G22gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT16), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n203), .B1(new_n204), .B2(G1gat), .ZN(new_n205));
  INV_X1    g004(.A(G8gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n203), .A2(G1gat), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n202), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(new_n208), .ZN(new_n210));
  NAND4_X1  g009(.A1(new_n210), .A2(KEYINPUT83), .A3(new_n206), .A4(new_n205), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n210), .A2(KEYINPUT82), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT82), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n205), .B1(new_n208), .B2(new_n214), .ZN(new_n215));
  OAI21_X1  g014(.A(G8gat), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n212), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT84), .ZN(new_n218));
  XOR2_X1   g017(.A(G43gat), .B(G50gat), .Z(new_n219));
  INV_X1    g018(.A(KEYINPUT15), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NOR2_X1   g020(.A1(G29gat), .A2(G36gat), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n222), .B(KEYINPUT14), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n219), .A2(new_n220), .ZN(new_n225));
  XNOR2_X1  g024(.A(KEYINPUT79), .B(G29gat), .ZN(new_n226));
  XNOR2_X1  g025(.A(KEYINPUT80), .B(G36gat), .ZN(new_n227));
  OAI21_X1  g026(.A(KEYINPUT81), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n226), .A2(new_n227), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT81), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND4_X1  g030(.A1(new_n224), .A2(new_n225), .A3(new_n228), .A4(new_n231), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n221), .B1(new_n229), .B2(new_n223), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  AND3_X1   g033(.A1(new_n217), .A2(new_n218), .A3(new_n234), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n218), .B1(new_n217), .B2(new_n234), .ZN(new_n236));
  OAI22_X1  g035(.A1(new_n235), .A2(new_n236), .B1(new_n234), .B2(new_n217), .ZN(new_n237));
  NAND2_X1  g036(.A1(G229gat), .A2(G233gat), .ZN(new_n238));
  XOR2_X1   g037(.A(new_n238), .B(KEYINPUT13), .Z(new_n239));
  NAND2_X1  g038(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  AND2_X1   g039(.A1(new_n212), .A2(new_n216), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT17), .ZN(new_n242));
  AND3_X1   g041(.A1(new_n232), .A2(new_n242), .A3(new_n233), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n242), .B1(new_n232), .B2(new_n233), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n241), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  OAI211_X1 g044(.A(new_n245), .B(new_n238), .C1(new_n235), .C2(new_n236), .ZN(new_n246));
  AND3_X1   g045(.A1(new_n246), .A2(KEYINPUT85), .A3(KEYINPUT18), .ZN(new_n247));
  AOI21_X1  g046(.A(KEYINPUT18), .B1(new_n246), .B2(KEYINPUT85), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n240), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(G113gat), .B(G141gat), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n250), .B(G197gat), .ZN(new_n251));
  XOR2_X1   g050(.A(KEYINPUT11), .B(G169gat), .Z(new_n252));
  XNOR2_X1  g051(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XOR2_X1   g052(.A(new_n253), .B(KEYINPUT12), .Z(new_n254));
  NAND2_X1  g053(.A1(new_n249), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n254), .ZN(new_n256));
  OAI211_X1 g055(.A(new_n240), .B(new_n256), .C1(new_n247), .C2(new_n248), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(G141gat), .ZN(new_n260));
  INV_X1    g059(.A(G148gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT2), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(KEYINPUT72), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT72), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(KEYINPUT2), .ZN(new_n266));
  NAND2_X1  g065(.A1(G141gat), .A2(G148gat), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n262), .A2(new_n264), .A3(new_n266), .A4(new_n267), .ZN(new_n268));
  XOR2_X1   g067(.A(G155gat), .B(G162gat), .Z(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(G155gat), .B(G162gat), .ZN(new_n271));
  INV_X1    g070(.A(G155gat), .ZN(new_n272));
  INV_X1    g071(.A(G162gat), .ZN(new_n273));
  OAI21_X1  g072(.A(KEYINPUT2), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n271), .A2(new_n262), .A3(new_n274), .A4(new_n267), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n270), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(KEYINPUT3), .ZN(new_n277));
  XNOR2_X1  g076(.A(KEYINPUT73), .B(KEYINPUT3), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n270), .A2(new_n275), .A3(new_n278), .ZN(new_n279));
  OR2_X1    g078(.A1(KEYINPUT68), .A2(G120gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(KEYINPUT68), .A2(G120gat), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n280), .A2(G113gat), .A3(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(G113gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(G120gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT1), .ZN(new_n286));
  INV_X1    g085(.A(G134gat), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n286), .B1(new_n287), .B2(G127gat), .ZN(new_n288));
  INV_X1    g087(.A(G127gat), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n289), .A2(G134gat), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n285), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n287), .A2(KEYINPUT67), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT67), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(G134gat), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n293), .A2(new_n295), .A3(G127gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n289), .A2(G134gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(G120gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(G113gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(new_n286), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n298), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n292), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n277), .A2(new_n279), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(G225gat), .A2(G233gat), .ZN(new_n306));
  NOR3_X1   g105(.A1(new_n304), .A2(new_n276), .A3(KEYINPUT4), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT4), .ZN(new_n308));
  AOI22_X1  g107(.A1(new_n285), .A2(new_n291), .B1(new_n298), .B2(new_n302), .ZN(new_n309));
  AND2_X1   g108(.A1(new_n270), .A2(new_n275), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n308), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  OAI211_X1 g110(.A(new_n305), .B(new_n306), .C1(new_n307), .C2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT5), .ZN(new_n313));
  AOI211_X1 g112(.A(new_n290), .B(new_n288), .C1(new_n282), .C2(new_n284), .ZN(new_n314));
  AOI22_X1  g113(.A1(new_n296), .A2(new_n297), .B1(new_n301), .B2(new_n286), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n276), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND4_X1  g115(.A1(new_n292), .A2(new_n303), .A3(new_n270), .A4(new_n275), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n306), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n313), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n312), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(KEYINPUT74), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT74), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n312), .A2(new_n320), .A3(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n312), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(new_n313), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n322), .A2(new_n324), .A3(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(G1gat), .B(G29gat), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n328), .B(KEYINPUT0), .ZN(new_n329));
  XNOR2_X1  g128(.A(G57gat), .B(G85gat), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n329), .B(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT6), .ZN(new_n333));
  INV_X1    g132(.A(new_n331), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n322), .A2(new_n326), .A3(new_n334), .A4(new_n324), .ZN(new_n335));
  NAND4_X1  g134(.A1(new_n332), .A2(KEYINPUT78), .A3(new_n333), .A4(new_n335), .ZN(new_n336));
  AOI22_X1  g135(.A1(new_n321), .A2(KEYINPUT74), .B1(new_n325), .B2(new_n313), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n334), .B1(new_n337), .B2(new_n324), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(KEYINPUT6), .ZN(new_n339));
  AND2_X1   g138(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n332), .A2(new_n333), .A3(new_n335), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT78), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g142(.A(KEYINPUT35), .B1(new_n340), .B2(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(KEYINPUT69), .B(KEYINPUT22), .ZN(new_n345));
  INV_X1    g144(.A(G211gat), .ZN(new_n346));
  INV_X1    g145(.A(G218gat), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n345), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(G197gat), .B(G204gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  XOR2_X1   g149(.A(G211gat), .B(G218gat), .Z(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n351), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n348), .A2(new_n353), .A3(new_n349), .ZN(new_n354));
  AND3_X1   g153(.A1(new_n352), .A2(KEYINPUT70), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(KEYINPUT70), .B1(new_n352), .B2(new_n354), .ZN(new_n356));
  OR2_X1    g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(G226gat), .A2(G233gat), .ZN(new_n358));
  XOR2_X1   g157(.A(new_n358), .B(KEYINPUT71), .Z(new_n359));
  XNOR2_X1  g158(.A(KEYINPUT27), .B(G183gat), .ZN(new_n360));
  INV_X1    g159(.A(G190gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT28), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n360), .A2(KEYINPUT28), .A3(new_n361), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(G183gat), .A2(G190gat), .ZN(new_n367));
  OAI21_X1  g166(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(G169gat), .A2(G176gat), .ZN(new_n369));
  NOR2_X1   g168(.A1(G169gat), .A2(G176gat), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT26), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n368), .A2(new_n369), .A3(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n366), .A2(new_n367), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n370), .A2(KEYINPUT23), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT23), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n376), .B1(G169gat), .B2(G176gat), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n375), .B1(new_n377), .B2(new_n370), .ZN(new_n378));
  NOR2_X1   g177(.A1(G183gat), .A2(G190gat), .ZN(new_n379));
  AND2_X1   g178(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n379), .B1(new_n380), .B2(G190gat), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT65), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT24), .ZN(new_n383));
  AND3_X1   g182(.A1(new_n367), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n382), .B1(new_n367), .B2(new_n383), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n381), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n378), .B1(new_n386), .B2(KEYINPUT66), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT66), .ZN(new_n388));
  OAI211_X1 g187(.A(new_n381), .B(new_n388), .C1(new_n384), .C2(new_n385), .ZN(new_n389));
  AOI21_X1  g188(.A(KEYINPUT25), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n391), .B1(G183gat), .B2(G190gat), .ZN(new_n392));
  AOI21_X1  g191(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT25), .ZN(new_n395));
  NOR3_X1   g194(.A1(new_n394), .A2(new_n378), .A3(new_n395), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n374), .B1(new_n390), .B2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT29), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n359), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n378), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n367), .A2(new_n383), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(KEYINPUT65), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n393), .A2(new_n382), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n392), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n400), .B1(new_n404), .B2(new_n388), .ZN(new_n405));
  INV_X1    g204(.A(new_n389), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n395), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n396), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n358), .B1(new_n409), .B2(new_n374), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n357), .B1(new_n399), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n352), .A2(new_n354), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n397), .A2(new_n359), .ZN(new_n413));
  AOI21_X1  g212(.A(KEYINPUT29), .B1(new_n409), .B2(new_n374), .ZN(new_n414));
  INV_X1    g213(.A(new_n358), .ZN(new_n415));
  OAI211_X1 g214(.A(new_n412), .B(new_n413), .C1(new_n414), .C2(new_n415), .ZN(new_n416));
  XNOR2_X1  g215(.A(G8gat), .B(G36gat), .ZN(new_n417));
  XNOR2_X1  g216(.A(G64gat), .B(G92gat), .ZN(new_n418));
  XOR2_X1   g217(.A(new_n417), .B(new_n418), .Z(new_n419));
  NAND3_X1  g218(.A1(new_n411), .A2(new_n416), .A3(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT30), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n411), .A2(new_n416), .ZN(new_n423));
  INV_X1    g222(.A(new_n419), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n411), .A2(new_n416), .A3(KEYINPUT30), .A4(new_n419), .ZN(new_n426));
  AND3_X1   g225(.A1(new_n422), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n386), .A2(KEYINPUT66), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n428), .A2(new_n389), .A3(new_n400), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n396), .B1(new_n429), .B2(new_n395), .ZN(new_n430));
  AND3_X1   g229(.A1(new_n366), .A2(new_n367), .A3(new_n373), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n309), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(G227gat), .A2(G233gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n433), .B(KEYINPUT64), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n374), .B(new_n304), .C1(new_n390), .C2(new_n396), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n432), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(KEYINPUT32), .ZN(new_n437));
  XOR2_X1   g236(.A(G15gat), .B(G43gat), .Z(new_n438));
  XNOR2_X1  g237(.A(G71gat), .B(G99gat), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n438), .B(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT33), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n441), .B1(new_n436), .B2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT34), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n432), .A2(new_n435), .ZN(new_n445));
  INV_X1    g244(.A(new_n434), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n444), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  AOI211_X1 g246(.A(KEYINPUT34), .B(new_n434), .C1(new_n432), .C2(new_n435), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n443), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  NOR3_X1   g249(.A1(new_n443), .A2(new_n447), .A3(new_n448), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n437), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  XNOR2_X1  g251(.A(G78gat), .B(G106gat), .ZN(new_n453));
  XNOR2_X1  g252(.A(KEYINPUT31), .B(G50gat), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n453), .B(new_n454), .ZN(new_n455));
  XOR2_X1   g254(.A(new_n455), .B(KEYINPUT75), .Z(new_n456));
  NAND2_X1  g255(.A1(new_n279), .A2(new_n398), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n457), .B1(new_n355), .B2(new_n356), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n310), .A2(KEYINPUT29), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(new_n412), .ZN(new_n460));
  AND3_X1   g259(.A1(new_n277), .A2(G228gat), .A3(G233gat), .ZN(new_n461));
  AND3_X1   g260(.A1(new_n458), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  XNOR2_X1  g261(.A(KEYINPUT76), .B(G22gat), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n278), .ZN(new_n465));
  AOI22_X1  g264(.A1(new_n459), .A2(new_n412), .B1(new_n276), .B2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n412), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(new_n457), .ZN(new_n468));
  AOI22_X1  g267(.A1(new_n466), .A2(new_n468), .B1(G228gat), .B2(G233gat), .ZN(new_n469));
  NOR3_X1   g268(.A1(new_n462), .A2(new_n464), .A3(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n469), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n458), .A2(new_n460), .A3(new_n461), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n463), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n456), .B1(new_n470), .B2(new_n473), .ZN(new_n474));
  OAI21_X1  g273(.A(G22gat), .B1(new_n462), .B2(new_n469), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n471), .A2(new_n463), .A3(new_n472), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n475), .A2(new_n476), .A3(new_n455), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n436), .A2(new_n442), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(new_n440), .ZN(new_n480));
  INV_X1    g279(.A(new_n447), .ZN(new_n481));
  INV_X1    g280(.A(new_n448), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n480), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n437), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n483), .A2(new_n484), .A3(new_n449), .ZN(new_n485));
  AND4_X1   g284(.A1(new_n427), .A2(new_n452), .A3(new_n478), .A4(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n344), .A2(new_n486), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n452), .A2(new_n427), .A3(new_n478), .A4(new_n485), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n341), .A2(new_n339), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  OAI21_X1  g289(.A(KEYINPUT35), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n487), .A2(new_n491), .ZN(new_n492));
  AND2_X1   g291(.A1(new_n476), .A2(new_n455), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n464), .B1(new_n462), .B2(new_n469), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(new_n476), .ZN(new_n495));
  AOI22_X1  g294(.A1(new_n493), .A2(new_n475), .B1(new_n495), .B2(new_n456), .ZN(new_n496));
  OAI21_X1  g295(.A(KEYINPUT39), .B1(new_n318), .B2(new_n319), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT77), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT77), .ZN(new_n499));
  OAI211_X1 g298(.A(new_n499), .B(KEYINPUT39), .C1(new_n318), .C2(new_n319), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n317), .A2(KEYINPUT4), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n309), .A2(new_n310), .A3(new_n308), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AND2_X1   g302(.A1(new_n503), .A2(new_n305), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n498), .B(new_n500), .C1(new_n504), .C2(new_n306), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n306), .B1(new_n503), .B2(new_n305), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT39), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n331), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  AND3_X1   g307(.A1(new_n505), .A2(KEYINPUT40), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g308(.A(KEYINPUT40), .B1(new_n505), .B2(new_n508), .ZN(new_n510));
  NOR3_X1   g309(.A1(new_n338), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n422), .A2(new_n425), .A3(new_n426), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n496), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n343), .A2(new_n339), .A3(new_n336), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT37), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n419), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n516), .B1(new_n423), .B2(new_n424), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n515), .B1(new_n411), .B2(new_n416), .ZN(new_n518));
  OAI21_X1  g317(.A(KEYINPUT38), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n431), .B1(new_n407), .B2(new_n408), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n358), .B1(new_n520), .B2(KEYINPUT29), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n412), .B1(new_n521), .B2(new_n413), .ZN(new_n522));
  NOR3_X1   g321(.A1(new_n399), .A2(new_n410), .A3(new_n357), .ZN(new_n523));
  OAI21_X1  g322(.A(KEYINPUT37), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT38), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n419), .B1(new_n411), .B2(new_n416), .ZN(new_n526));
  OAI211_X1 g325(.A(new_n524), .B(new_n525), .C1(new_n526), .C2(new_n516), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n519), .A2(new_n420), .A3(new_n527), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n513), .B1(new_n514), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n489), .A2(new_n427), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(new_n496), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT36), .ZN(new_n532));
  AND3_X1   g331(.A1(new_n483), .A2(new_n484), .A3(new_n449), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n484), .B1(new_n483), .B2(new_n449), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n452), .A2(KEYINPUT36), .A3(new_n485), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n529), .A2(new_n531), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n259), .B1(new_n492), .B2(new_n538), .ZN(new_n539));
  AND2_X1   g338(.A1(G71gat), .A2(G78gat), .ZN(new_n540));
  NOR2_X1   g339(.A1(G71gat), .A2(G78gat), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(G57gat), .B(G64gat), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT86), .ZN(new_n544));
  OAI22_X1  g343(.A1(new_n543), .A2(new_n544), .B1(KEYINPUT9), .B2(new_n540), .ZN(new_n545));
  AND2_X1   g344(.A1(new_n543), .A2(new_n544), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n542), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(G57gat), .ZN(new_n548));
  OAI21_X1  g347(.A(KEYINPUT87), .B1(new_n548), .B2(G64gat), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT87), .ZN(new_n550));
  INV_X1    g349(.A(G64gat), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n550), .A2(new_n551), .A3(G57gat), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n548), .A2(G64gat), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n549), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(KEYINPUT88), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n540), .A2(KEYINPUT9), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n542), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT88), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n549), .A2(new_n552), .A3(new_n558), .A4(new_n553), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n555), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(KEYINPUT21), .B1(new_n547), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(G231gat), .A2(G233gat), .ZN(new_n562));
  XOR2_X1   g361(.A(new_n561), .B(new_n562), .Z(new_n563));
  XNOR2_X1  g362(.A(new_n563), .B(new_n289), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n547), .A2(new_n560), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(KEYINPUT89), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT89), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n547), .A2(new_n560), .A3(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n566), .A2(KEYINPUT21), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(new_n241), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n564), .B(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(G155gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(G183gat), .B(G211gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n571), .B(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(G232gat), .ZN(new_n577));
  INV_X1    g376(.A(G233gat), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n579), .A2(KEYINPUT41), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n580), .B(G134gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(new_n273), .ZN(new_n582));
  INV_X1    g381(.A(new_n579), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT41), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n234), .ZN(new_n587));
  XNOR2_X1  g386(.A(G99gat), .B(G106gat), .ZN(new_n588));
  NAND3_X1  g387(.A1(KEYINPUT90), .A2(G85gat), .A3(G92gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(KEYINPUT7), .ZN(new_n590));
  NAND2_X1  g389(.A1(G99gat), .A2(G106gat), .ZN(new_n591));
  INV_X1    g390(.A(G85gat), .ZN(new_n592));
  INV_X1    g391(.A(G92gat), .ZN(new_n593));
  AOI22_X1  g392(.A1(KEYINPUT8), .A2(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n588), .B1(new_n590), .B2(new_n594), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n595), .A2(KEYINPUT91), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  AND3_X1   g396(.A1(new_n590), .A2(new_n588), .A3(new_n594), .ZN(new_n598));
  OAI21_X1  g397(.A(KEYINPUT91), .B1(new_n598), .B2(new_n595), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n586), .B1(new_n587), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(KEYINPUT92), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT91), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n590), .A2(new_n594), .ZN(new_n604));
  INV_X1    g403(.A(new_n588), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n590), .A2(new_n588), .A3(new_n594), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n603), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n608), .A2(new_n596), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n609), .A2(new_n234), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT92), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n610), .A2(new_n611), .A3(new_n586), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n243), .A2(new_n244), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  AOI22_X1  g413(.A1(new_n602), .A2(new_n612), .B1(new_n614), .B2(new_n600), .ZN(new_n615));
  XNOR2_X1  g414(.A(G190gat), .B(G218gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(KEYINPUT93), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT94), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n582), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n602), .A2(new_n612), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n614), .A2(new_n600), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(new_n617), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n615), .A2(new_n618), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n621), .A2(new_n627), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n625), .A2(new_n620), .A3(new_n626), .A4(new_n582), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n576), .A2(new_n630), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n565), .B1(new_n608), .B2(new_n596), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n606), .A2(new_n607), .ZN(new_n633));
  OAI21_X1  g432(.A(KEYINPUT95), .B1(new_n565), .B2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT10), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n598), .A2(new_n595), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT95), .ZN(new_n637));
  NAND4_X1  g436(.A1(new_n636), .A2(new_n637), .A3(new_n547), .A4(new_n560), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n632), .A2(new_n634), .A3(new_n635), .A4(new_n638), .ZN(new_n639));
  NAND4_X1  g438(.A1(new_n609), .A2(KEYINPUT10), .A3(new_n566), .A4(new_n568), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(G230gat), .A2(G233gat), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n632), .A2(new_n638), .A3(new_n634), .ZN(new_n644));
  INV_X1    g443(.A(new_n642), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(G120gat), .B(G148gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(G176gat), .B(G204gat), .ZN(new_n649));
  XOR2_X1   g448(.A(new_n648), .B(new_n649), .Z(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n647), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n647), .A2(new_n651), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n631), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n539), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(KEYINPUT96), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(new_n490), .ZN(new_n659));
  XOR2_X1   g458(.A(KEYINPUT97), .B(G1gat), .Z(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(G1324gat));
  AND2_X1   g460(.A1(new_n657), .A2(KEYINPUT96), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n657), .A2(KEYINPUT96), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n664), .A2(new_n427), .ZN(new_n665));
  XOR2_X1   g464(.A(KEYINPUT16), .B(G8gat), .Z(new_n666));
  AND2_X1   g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  OR2_X1    g466(.A1(new_n667), .A2(KEYINPUT42), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(KEYINPUT42), .ZN(new_n669));
  OAI21_X1  g468(.A(G8gat), .B1(new_n664), .B2(new_n427), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n668), .A2(new_n669), .A3(new_n670), .ZN(G1325gat));
  OAI21_X1  g470(.A(G15gat), .B1(new_n664), .B2(new_n537), .ZN(new_n672));
  INV_X1    g471(.A(G15gat), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n533), .A2(new_n534), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n658), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g475(.A(new_n676), .B(KEYINPUT98), .Z(G1326gat));
  OR3_X1    g476(.A1(new_n664), .A2(KEYINPUT99), .A3(new_n478), .ZN(new_n678));
  OAI21_X1  g477(.A(KEYINPUT99), .B1(new_n664), .B2(new_n478), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g479(.A(KEYINPUT43), .B(G22gat), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n680), .B(new_n681), .ZN(G1327gat));
  AOI21_X1  g481(.A(new_n512), .B1(new_n339), .B2(new_n341), .ZN(new_n683));
  OAI21_X1  g482(.A(KEYINPUT101), .B1(new_n683), .B2(new_n478), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT101), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n530), .A2(new_n685), .A3(new_n496), .ZN(new_n686));
  NAND4_X1  g485(.A1(new_n529), .A2(new_n684), .A3(new_n537), .A4(new_n686), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n630), .B1(new_n492), .B2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n492), .A2(new_n538), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n630), .A2(new_n690), .ZN(new_n692));
  AOI22_X1  g491(.A1(new_n689), .A2(new_n690), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n576), .ZN(new_n694));
  INV_X1    g493(.A(new_n655), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n694), .A2(new_n258), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(KEYINPUT100), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n693), .A2(new_n490), .A3(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT102), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n226), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n700), .B1(new_n699), .B2(new_n698), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n576), .A2(new_n630), .A3(new_n655), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n539), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n704), .A2(new_n490), .A3(new_n226), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT45), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n701), .A2(new_n706), .ZN(G1328gat));
  NAND3_X1  g506(.A1(new_n704), .A2(new_n512), .A3(new_n227), .ZN(new_n708));
  OR2_X1    g507(.A1(new_n708), .A2(KEYINPUT46), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(KEYINPUT46), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n693), .A2(new_n697), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n711), .A2(new_n427), .ZN(new_n712));
  OAI211_X1 g511(.A(new_n709), .B(new_n710), .C1(new_n712), .C2(new_n227), .ZN(G1329gat));
  INV_X1    g512(.A(new_n537), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(G43gat), .ZN(new_n715));
  INV_X1    g514(.A(new_n674), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n703), .A2(new_n716), .ZN(new_n717));
  OAI22_X1  g516(.A1(new_n711), .A2(new_n715), .B1(G43gat), .B2(new_n717), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g518(.A(G50gat), .B1(new_n711), .B2(new_n478), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n478), .A2(G50gat), .ZN(new_n721));
  XOR2_X1   g520(.A(new_n721), .B(KEYINPUT103), .Z(new_n722));
  OAI21_X1  g521(.A(new_n720), .B1(new_n703), .B2(new_n722), .ZN(new_n723));
  XOR2_X1   g522(.A(new_n723), .B(KEYINPUT48), .Z(G1331gat));
  NAND2_X1  g523(.A1(new_n492), .A2(new_n687), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n631), .A2(new_n258), .A3(new_n695), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n727), .A2(new_n489), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(new_n548), .ZN(G1332gat));
  INV_X1    g528(.A(new_n727), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT49), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n512), .B1(new_n731), .B2(new_n551), .ZN(new_n732));
  XOR2_X1   g531(.A(new_n732), .B(KEYINPUT104), .Z(new_n733));
  NAND2_X1  g532(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n731), .A2(new_n551), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n734), .B(new_n735), .ZN(G1333gat));
  NOR3_X1   g535(.A1(new_n727), .A2(G71gat), .A3(new_n716), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n730), .A2(new_n714), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n737), .B1(G71gat), .B2(new_n738), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g539(.A1(new_n727), .A2(new_n478), .ZN(new_n741));
  XNOR2_X1  g540(.A(KEYINPUT105), .B(G78gat), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n741), .B(new_n742), .ZN(G1335gat));
  INV_X1    g542(.A(new_n630), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n576), .A2(new_n258), .ZN(new_n745));
  AND4_X1   g544(.A1(new_n529), .A2(new_n684), .A3(new_n537), .A4(new_n686), .ZN(new_n746));
  NAND4_X1  g545(.A1(new_n674), .A2(new_n489), .A3(new_n427), .A4(new_n478), .ZN(new_n747));
  AOI22_X1  g546(.A1(new_n747), .A2(KEYINPUT35), .B1(new_n344), .B2(new_n486), .ZN(new_n748));
  OAI211_X1 g547(.A(new_n744), .B(new_n745), .C1(new_n746), .C2(new_n748), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n695), .B1(new_n749), .B2(KEYINPUT51), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT51), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n688), .A2(new_n751), .A3(new_n745), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(new_n753), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n754), .A2(new_n592), .A3(new_n490), .ZN(new_n755));
  AND3_X1   g554(.A1(new_n529), .A2(new_n531), .A3(new_n537), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n692), .B1(new_n756), .B2(new_n748), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n576), .A2(new_n258), .A3(new_n695), .ZN(new_n758));
  OAI211_X1 g557(.A(new_n757), .B(new_n758), .C1(new_n688), .C2(KEYINPUT44), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT106), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(new_n420), .ZN(new_n762));
  INV_X1    g561(.A(new_n517), .ZN(new_n763));
  AND2_X1   g562(.A1(new_n397), .A2(new_n359), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n415), .B1(new_n397), .B2(new_n398), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n467), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  OAI22_X1  g565(.A1(new_n414), .A2(new_n359), .B1(new_n520), .B2(new_n358), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n766), .B1(new_n767), .B2(new_n357), .ZN(new_n768));
  AOI21_X1  g567(.A(KEYINPUT38), .B1(new_n768), .B2(KEYINPUT37), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n762), .B1(new_n763), .B2(new_n769), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n340), .A2(new_n343), .A3(new_n770), .A4(new_n519), .ZN(new_n771));
  AOI22_X1  g570(.A1(new_n771), .A2(new_n513), .B1(new_n536), .B2(new_n535), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n685), .B1(new_n530), .B2(new_n496), .ZN(new_n773));
  AOI211_X1 g572(.A(KEYINPUT101), .B(new_n478), .C1(new_n489), .C2(new_n427), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  AOI22_X1  g574(.A1(new_n772), .A2(new_n775), .B1(new_n491), .B2(new_n487), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n690), .B1(new_n776), .B2(new_n630), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n777), .A2(KEYINPUT106), .A3(new_n757), .A4(new_n758), .ZN(new_n778));
  AND2_X1   g577(.A1(new_n761), .A2(new_n778), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n779), .A2(new_n490), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n755), .B1(new_n780), .B2(new_n592), .ZN(G1336gat));
  OAI21_X1  g580(.A(G92gat), .B1(new_n759), .B2(new_n427), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n749), .A2(KEYINPUT51), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n427), .A2(G92gat), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n783), .A2(new_n655), .A3(new_n752), .A4(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT52), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n782), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT107), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n785), .A2(new_n788), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n750), .A2(KEYINPUT107), .A3(new_n752), .A4(new_n784), .ZN(new_n790));
  AND2_X1   g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n761), .A2(new_n778), .A3(new_n512), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(G92gat), .ZN(new_n793));
  AOI211_X1 g592(.A(KEYINPUT108), .B(new_n786), .C1(new_n791), .C2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT108), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n793), .A2(new_n789), .A3(new_n790), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n795), .B1(new_n796), .B2(KEYINPUT52), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n787), .B1(new_n794), .B2(new_n797), .ZN(G1337gat));
  AOI21_X1  g597(.A(G99gat), .B1(new_n754), .B2(new_n674), .ZN(new_n799));
  AND2_X1   g598(.A1(new_n714), .A2(G99gat), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n799), .B1(new_n779), .B2(new_n800), .ZN(G1338gat));
  NOR3_X1   g600(.A1(new_n753), .A2(G106gat), .A3(new_n478), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n802), .A2(KEYINPUT53), .ZN(new_n803));
  OAI21_X1  g602(.A(G106gat), .B1(new_n759), .B2(new_n478), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n779), .A2(new_n496), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n802), .B1(new_n806), .B2(G106gat), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT53), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n805), .B1(new_n807), .B2(new_n808), .ZN(G1339gat));
  NAND3_X1  g608(.A1(new_n639), .A2(new_n640), .A3(new_n645), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(KEYINPUT109), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT109), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n639), .A2(new_n640), .A3(new_n812), .A4(new_n645), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n811), .A2(new_n643), .A3(KEYINPUT54), .A4(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n645), .B1(new_n639), .B2(new_n640), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT54), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n650), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT55), .ZN(new_n819));
  AOI21_X1  g618(.A(KEYINPUT111), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT111), .ZN(new_n821));
  AOI211_X1 g620(.A(new_n821), .B(KEYINPUT55), .C1(new_n814), .C2(new_n817), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n814), .A2(KEYINPUT110), .A3(KEYINPUT55), .A4(new_n817), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n814), .A2(KEYINPUT55), .A3(new_n817), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT110), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n652), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n823), .A2(new_n258), .A3(new_n824), .A4(new_n827), .ZN(new_n828));
  OR2_X1    g627(.A1(new_n235), .A2(new_n236), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n238), .B1(new_n829), .B2(new_n245), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n237), .A2(new_n239), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n253), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n257), .A2(new_n655), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n744), .B1(new_n828), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n821), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n818), .A2(KEYINPUT111), .A3(new_n819), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n836), .A2(new_n827), .A3(new_n824), .A4(new_n837), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n628), .A2(new_n257), .A3(new_n629), .A4(new_n832), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n694), .B1(new_n834), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n656), .A2(new_n259), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n496), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n843), .A2(new_n490), .A3(new_n427), .A4(new_n674), .ZN(new_n844));
  NOR3_X1   g643(.A1(new_n844), .A2(new_n283), .A3(new_n259), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n489), .B1(new_n841), .B2(new_n842), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n846), .A2(new_n486), .ZN(new_n847));
  AOI21_X1  g646(.A(G113gat), .B1(new_n847), .B2(new_n258), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g648(.A(new_n849), .B(KEYINPUT112), .ZN(G1340gat));
  NAND4_X1  g649(.A1(new_n847), .A2(new_n280), .A3(new_n281), .A4(new_n655), .ZN(new_n851));
  OAI21_X1  g650(.A(G120gat), .B1(new_n844), .B2(new_n695), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g652(.A(new_n853), .B(KEYINPUT113), .ZN(G1341gat));
  OAI21_X1  g653(.A(G127gat), .B1(new_n844), .B2(new_n694), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n847), .A2(new_n289), .A3(new_n576), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(G1342gat));
  NAND4_X1  g656(.A1(new_n847), .A2(new_n293), .A3(new_n295), .A4(new_n744), .ZN(new_n858));
  OR2_X1    g657(.A1(new_n858), .A2(KEYINPUT56), .ZN(new_n859));
  OAI21_X1  g658(.A(G134gat), .B1(new_n844), .B2(new_n630), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n858), .A2(KEYINPUT56), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(G1343gat));
  INV_X1    g661(.A(KEYINPUT58), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n714), .A2(new_n478), .ZN(new_n864));
  INV_X1    g663(.A(new_n864), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n865), .A2(new_n512), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n846), .A2(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n258), .A2(new_n260), .ZN(new_n869));
  XNOR2_X1  g668(.A(new_n869), .B(KEYINPUT117), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT116), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n863), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n490), .A2(new_n427), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n714), .A2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(new_n875), .ZN(new_n876));
  NAND4_X1  g675(.A1(new_n258), .A2(new_n824), .A3(new_n827), .A4(new_n835), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(new_n833), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(new_n630), .ZN(new_n879));
  INV_X1    g678(.A(new_n840), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n576), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT115), .ZN(new_n882));
  AOI22_X1  g681(.A1(new_n881), .A2(new_n882), .B1(new_n259), .B2(new_n656), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n744), .B1(new_n877), .B2(new_n833), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n694), .B1(new_n884), .B2(new_n840), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(KEYINPUT115), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT57), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n478), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n833), .B1(new_n838), .B2(new_n259), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n840), .B1(new_n891), .B2(new_n630), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n842), .B1(new_n892), .B2(new_n576), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(new_n496), .ZN(new_n894));
  XNOR2_X1  g693(.A(KEYINPUT114), .B(KEYINPUT57), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n876), .B1(new_n890), .B2(new_n896), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n260), .B1(new_n897), .B2(new_n258), .ZN(new_n898));
  INV_X1    g697(.A(new_n871), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n873), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n894), .A2(new_n895), .ZN(new_n901));
  INV_X1    g700(.A(new_n889), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n902), .B1(new_n883), .B2(new_n886), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n875), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g703(.A(G141gat), .B1(new_n904), .B2(new_n259), .ZN(new_n905));
  OAI211_X1 g704(.A(new_n905), .B(new_n871), .C1(new_n872), .C2(new_n863), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n900), .A2(new_n906), .ZN(G1344gat));
  INV_X1    g706(.A(KEYINPUT59), .ZN(new_n908));
  OAI211_X1 g707(.A(new_n908), .B(G148gat), .C1(new_n904), .C2(new_n695), .ZN(new_n909));
  AOI211_X1 g708(.A(new_n478), .B(new_n895), .C1(new_n841), .C2(new_n842), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n885), .A2(new_n842), .ZN(new_n911));
  AOI21_X1  g710(.A(KEYINPUT57), .B1(new_n911), .B2(new_n496), .ZN(new_n912));
  OAI211_X1 g711(.A(new_n655), .B(new_n875), .C1(new_n910), .C2(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(G148gat), .ZN(new_n914));
  AOI21_X1  g713(.A(KEYINPUT118), .B1(new_n914), .B2(KEYINPUT59), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT118), .ZN(new_n916));
  AOI211_X1 g715(.A(new_n916), .B(new_n908), .C1(new_n913), .C2(G148gat), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n909), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n868), .A2(new_n261), .A3(new_n655), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(G1345gat));
  INV_X1    g719(.A(KEYINPUT119), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n272), .B1(new_n897), .B2(new_n576), .ZN(new_n922));
  NOR3_X1   g721(.A1(new_n867), .A2(G155gat), .A3(new_n694), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n921), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g723(.A(G155gat), .B1(new_n904), .B2(new_n694), .ZN(new_n925));
  INV_X1    g724(.A(new_n923), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n925), .A2(KEYINPUT119), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n924), .A2(new_n927), .ZN(G1346gat));
  AOI21_X1  g727(.A(G162gat), .B1(new_n868), .B2(new_n744), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n630), .A2(new_n273), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n929), .B1(new_n897), .B2(new_n930), .ZN(G1347gat));
  NOR3_X1   g730(.A1(new_n716), .A2(new_n427), .A3(new_n496), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT120), .ZN(new_n933));
  AOI211_X1 g732(.A(new_n933), .B(new_n490), .C1(new_n841), .C2(new_n842), .ZN(new_n934));
  AOI21_X1  g733(.A(KEYINPUT120), .B1(new_n893), .B2(new_n489), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n932), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT121), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OAI211_X1 g737(.A(KEYINPUT121), .B(new_n932), .C1(new_n934), .C2(new_n935), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n259), .A2(G169gat), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT122), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n490), .A2(new_n427), .ZN(new_n944));
  AND2_X1   g743(.A1(new_n944), .A2(new_n674), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n843), .A2(new_n258), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g745(.A(KEYINPUT122), .B1(new_n946), .B2(G169gat), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n943), .B1(new_n941), .B2(new_n947), .ZN(G1348gat));
  NOR2_X1   g747(.A1(new_n695), .A2(G176gat), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n938), .A2(new_n939), .A3(new_n949), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n843), .A2(new_n655), .A3(new_n945), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(G176gat), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n950), .A2(new_n952), .ZN(G1349gat));
  NOR2_X1   g752(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n954));
  INV_X1    g753(.A(new_n954), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n576), .A2(new_n360), .ZN(new_n956));
  OAI21_X1  g755(.A(KEYINPUT123), .B1(new_n936), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n893), .A2(new_n489), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n958), .A2(new_n933), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n893), .A2(KEYINPUT120), .A3(new_n489), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT123), .ZN(new_n962));
  INV_X1    g761(.A(new_n956), .ZN(new_n963));
  NAND4_X1  g762(.A1(new_n961), .A2(new_n962), .A3(new_n932), .A4(new_n963), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n957), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n843), .A2(new_n576), .A3(new_n945), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(G183gat), .ZN(new_n967));
  NAND2_X1  g766(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g768(.A(new_n969), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n955), .B1(new_n965), .B2(new_n970), .ZN(new_n971));
  AOI211_X1 g770(.A(new_n954), .B(new_n969), .C1(new_n957), .C2(new_n964), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n971), .A2(new_n972), .ZN(G1350gat));
  NOR2_X1   g772(.A1(new_n630), .A2(G190gat), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n938), .A2(new_n939), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n975), .A2(KEYINPUT125), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT125), .ZN(new_n977));
  NAND4_X1  g776(.A1(new_n938), .A2(new_n977), .A3(new_n939), .A4(new_n974), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n843), .A2(new_n744), .A3(new_n945), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n980), .A2(G190gat), .ZN(new_n981));
  XNOR2_X1  g780(.A(new_n981), .B(KEYINPUT61), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n979), .A2(new_n982), .ZN(G1351gat));
  INV_X1    g782(.A(KEYINPUT126), .ZN(new_n984));
  NOR4_X1   g783(.A1(new_n714), .A2(new_n984), .A3(new_n490), .A4(new_n427), .ZN(new_n985));
  AOI21_X1  g784(.A(KEYINPUT126), .B1(new_n537), .B2(new_n944), .ZN(new_n986));
  NOR2_X1   g785(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g786(.A(new_n910), .ZN(new_n988));
  INV_X1    g787(.A(new_n912), .ZN(new_n989));
  AOI21_X1  g788(.A(new_n987), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  INV_X1    g789(.A(new_n990), .ZN(new_n991));
  OAI21_X1  g790(.A(G197gat), .B1(new_n991), .B2(new_n259), .ZN(new_n992));
  AOI211_X1 g791(.A(new_n427), .B(new_n865), .C1(new_n959), .C2(new_n960), .ZN(new_n993));
  INV_X1    g792(.A(G197gat), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n993), .A2(new_n994), .A3(new_n258), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n992), .A2(new_n995), .ZN(G1352gat));
  XOR2_X1   g795(.A(KEYINPUT127), .B(G204gat), .Z(new_n997));
  NOR2_X1   g796(.A1(new_n695), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n993), .A2(new_n998), .ZN(new_n999));
  OR2_X1    g798(.A1(new_n999), .A2(KEYINPUT62), .ZN(new_n1000));
  OAI221_X1 g799(.A(new_n655), .B1(new_n985), .B2(new_n986), .C1(new_n910), .C2(new_n912), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n1001), .A2(new_n997), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n999), .A2(KEYINPUT62), .ZN(new_n1003));
  NAND3_X1  g802(.A1(new_n1000), .A2(new_n1002), .A3(new_n1003), .ZN(G1353gat));
  NAND3_X1  g803(.A1(new_n993), .A2(new_n346), .A3(new_n576), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n990), .A2(new_n576), .ZN(new_n1006));
  AND3_X1   g805(.A1(new_n1006), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1007));
  AOI21_X1  g806(.A(KEYINPUT63), .B1(new_n1006), .B2(G211gat), .ZN(new_n1008));
  OAI21_X1  g807(.A(new_n1005), .B1(new_n1007), .B2(new_n1008), .ZN(G1354gat));
  OAI21_X1  g808(.A(G218gat), .B1(new_n991), .B2(new_n630), .ZN(new_n1010));
  NAND3_X1  g809(.A1(new_n993), .A2(new_n347), .A3(new_n744), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n1010), .A2(new_n1011), .ZN(G1355gat));
endmodule


