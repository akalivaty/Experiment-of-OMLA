

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730;

  NAND2_X1 U366 ( .A1(n714), .A2(n705), .ZN(n361) );
  XNOR2_X1 U367 ( .A(n399), .B(n463), .ZN(n701) );
  INV_X1 U368 ( .A(G953), .ZN(n715) );
  NOR2_X2 U369 ( .A1(n532), .A2(n422), .ZN(n424) );
  XNOR2_X2 U370 ( .A(n590), .B(n349), .ZN(n705) );
  XNOR2_X1 U371 ( .A(n383), .B(G122), .ZN(n444) );
  INV_X1 U372 ( .A(G116), .ZN(n383) );
  NAND2_X2 U373 ( .A1(n355), .A2(n354), .ZN(n617) );
  AND2_X1 U374 ( .A1(n580), .A2(n579), .ZN(n589) );
  OR2_X1 U375 ( .A1(n582), .A2(n554), .ZN(n555) );
  XNOR2_X1 U376 ( .A(n384), .B(n496), .ZN(n582) );
  XNOR2_X1 U377 ( .A(n375), .B(KEYINPUT105), .ZN(n724) );
  BUF_X1 U378 ( .A(n559), .Z(n570) );
  XNOR2_X1 U379 ( .A(n524), .B(n416), .ZN(n532) );
  XNOR2_X1 U380 ( .A(n492), .B(KEYINPUT6), .ZN(n558) );
  XNOR2_X1 U381 ( .A(n477), .B(n476), .ZN(n625) );
  XNOR2_X1 U382 ( .A(G146), .B(G125), .ZN(n428) );
  XNOR2_X1 U383 ( .A(n713), .B(n390), .ZN(n478) );
  XNOR2_X1 U384 ( .A(n557), .B(KEYINPUT75), .ZN(n353) );
  XNOR2_X1 U385 ( .A(n424), .B(n348), .ZN(n559) );
  AND2_X1 U386 ( .A1(n553), .A2(n552), .ZN(n714) );
  NAND2_X1 U387 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U388 ( .A(n362), .B(n351), .ZN(n548) );
  NOR2_X1 U389 ( .A1(n729), .A2(n730), .ZN(n362) );
  XNOR2_X1 U390 ( .A(n428), .B(n427), .ZN(n467) );
  INV_X1 U391 ( .A(KEYINPUT85), .ZN(n414) );
  NOR2_X1 U392 ( .A1(n515), .A2(n501), .ZN(n508) );
  XNOR2_X1 U393 ( .A(n465), .B(G469), .ZN(n516) );
  XNOR2_X1 U394 ( .A(n467), .B(n468), .ZN(n712) );
  XNOR2_X1 U395 ( .A(n473), .B(n368), .ZN(n367) );
  XNOR2_X1 U396 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n368) );
  XNOR2_X1 U397 ( .A(G128), .B(G119), .ZN(n471) );
  AND2_X1 U398 ( .A1(n593), .A2(KEYINPUT2), .ZN(n386) );
  INV_X1 U399 ( .A(n361), .ZN(n360) );
  NAND2_X1 U400 ( .A1(n359), .A2(n357), .ZN(n356) );
  NAND2_X1 U401 ( .A1(n358), .A2(n595), .ZN(n357) );
  NAND2_X1 U402 ( .A1(n386), .A2(KEYINPUT77), .ZN(n359) );
  INV_X1 U403 ( .A(n594), .ZN(n358) );
  INV_X1 U404 ( .A(n558), .ZN(n352) );
  INV_X1 U405 ( .A(KEYINPUT39), .ZN(n520) );
  AND2_X1 U406 ( .A1(n372), .A2(n369), .ZN(n521) );
  INV_X1 U407 ( .A(n534), .ZN(n369) );
  INV_X1 U408 ( .A(G472), .ZN(n377) );
  AND2_X1 U409 ( .A1(n596), .A2(n487), .ZN(n378) );
  XNOR2_X1 U410 ( .A(n457), .B(n456), .ZN(n493) );
  INV_X1 U411 ( .A(KEYINPUT80), .ZN(n380) );
  NAND2_X1 U412 ( .A1(n344), .A2(n382), .ZN(n381) );
  NOR2_X1 U413 ( .A1(G953), .A2(G237), .ZN(n479) );
  XNOR2_X1 U414 ( .A(G137), .B(G116), .ZN(n482) );
  XNOR2_X1 U415 ( .A(n460), .B(n459), .ZN(n713) );
  XNOR2_X1 U416 ( .A(n458), .B(KEYINPUT4), .ZN(n459) );
  XNOR2_X1 U417 ( .A(G131), .B(KEYINPUT72), .ZN(n458) );
  XNOR2_X1 U418 ( .A(KEYINPUT3), .B(G119), .ZN(n393) );
  XOR2_X1 U419 ( .A(KEYINPUT89), .B(G110), .Z(n472) );
  XNOR2_X1 U420 ( .A(G113), .B(G143), .ZN(n425) );
  INV_X1 U421 ( .A(KEYINPUT71), .ZN(n402) );
  XNOR2_X1 U422 ( .A(G143), .B(G128), .ZN(n440) );
  NOR2_X1 U423 ( .A1(n535), .A2(n518), .ZN(n372) );
  XNOR2_X1 U424 ( .A(n439), .B(n438), .ZN(n536) );
  XNOR2_X1 U425 ( .A(n437), .B(G475), .ZN(n438) );
  XNOR2_X1 U426 ( .A(n440), .B(G134), .ZN(n460) );
  XNOR2_X1 U427 ( .A(n361), .B(n591), .ZN(n387) );
  NOR2_X1 U428 ( .A1(n662), .A2(n560), .ZN(n561) );
  AND2_X1 U429 ( .A1(n494), .A2(n558), .ZN(n385) );
  XNOR2_X1 U430 ( .A(KEYINPUT91), .B(n569), .ZN(n635) );
  NAND2_X1 U431 ( .A1(n370), .A2(n517), .ZN(n534) );
  XNOR2_X1 U432 ( .A(n567), .B(n371), .ZN(n370) );
  INV_X1 U433 ( .A(KEYINPUT102), .ZN(n371) );
  AND2_X1 U434 ( .A1(n508), .A2(n492), .ZN(n509) );
  XNOR2_X1 U435 ( .A(n366), .B(n365), .ZN(n619) );
  INV_X1 U436 ( .A(n712), .ZN(n365) );
  XNOR2_X1 U437 ( .A(n470), .B(n367), .ZN(n366) );
  NAND2_X1 U438 ( .A1(n361), .A2(n350), .ZN(n354) );
  NAND2_X1 U439 ( .A1(n360), .A2(n356), .ZN(n355) );
  AND2_X1 U440 ( .A1(n599), .A2(G953), .ZN(n700) );
  XNOR2_X1 U441 ( .A(n364), .B(n363), .ZN(n729) );
  INV_X1 U442 ( .A(KEYINPUT40), .ZN(n363) );
  NAND2_X1 U443 ( .A1(n376), .A2(n556), .ZN(n375) );
  XNOR2_X1 U444 ( .A(n527), .B(KEYINPUT36), .ZN(n376) );
  NOR2_X1 U445 ( .A1(n526), .A2(n525), .ZN(n527) );
  OR2_X1 U446 ( .A1(n533), .A2(n532), .ZN(n680) );
  AND2_X1 U447 ( .A1(n493), .A2(n558), .ZN(n577) );
  XNOR2_X1 U448 ( .A(n667), .B(n379), .ZN(G75) );
  INV_X1 U449 ( .A(KEYINPUT53), .ZN(n379) );
  OR2_X1 U450 ( .A1(n361), .A2(n594), .ZN(n344) );
  XOR2_X1 U451 ( .A(n433), .B(n432), .Z(n345) );
  AND2_X1 U452 ( .A1(n353), .A2(n352), .ZN(n346) );
  AND2_X1 U453 ( .A1(n542), .A2(n374), .ZN(n347) );
  XOR2_X1 U454 ( .A(n423), .B(KEYINPUT0), .Z(n348) );
  XOR2_X1 U455 ( .A(KEYINPUT65), .B(KEYINPUT45), .Z(n349) );
  AND2_X1 U456 ( .A1(n386), .A2(n591), .ZN(n350) );
  XNOR2_X1 U457 ( .A(n522), .B(KEYINPUT64), .ZN(n351) );
  NAND2_X1 U458 ( .A1(n353), .A2(n492), .ZN(n569) );
  XNOR2_X2 U459 ( .A(n411), .B(n410), .ZN(n506) );
  NAND2_X1 U460 ( .A1(n550), .A2(n529), .ZN(n364) );
  NOR2_X1 U461 ( .A1(n724), .A2(n373), .ZN(n546) );
  NAND2_X1 U462 ( .A1(n545), .A2(n347), .ZN(n373) );
  AND2_X1 U463 ( .A1(n541), .A2(n543), .ZN(n374) );
  NOR2_X1 U464 ( .A1(n558), .A2(n682), .ZN(n502) );
  XNOR2_X2 U465 ( .A(n378), .B(n377), .ZN(n492) );
  XNOR2_X1 U466 ( .A(n381), .B(n380), .ZN(n666) );
  NAND2_X1 U467 ( .A1(n387), .A2(KEYINPUT2), .ZN(n382) );
  NAND2_X1 U468 ( .A1(n493), .A2(n385), .ZN(n384) );
  XNOR2_X1 U469 ( .A(n478), .B(n389), .ZN(n690) );
  NOR2_X1 U470 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X2 U471 ( .A(n415), .B(n414), .ZN(n524) );
  NAND2_X1 U472 ( .A1(n581), .A2(KEYINPUT44), .ZN(n388) );
  XOR2_X1 U473 ( .A(n464), .B(n463), .Z(n389) );
  XOR2_X1 U474 ( .A(n461), .B(G146), .Z(n390) );
  NAND2_X1 U475 ( .A1(n555), .A2(KEYINPUT84), .ZN(n391) );
  NOR2_X1 U476 ( .A1(n529), .A2(n671), .ZN(n530) );
  XOR2_X1 U477 ( .A(KEYINPUT98), .B(n530), .Z(n573) );
  INV_X1 U478 ( .A(KEYINPUT46), .ZN(n522) );
  INV_X1 U479 ( .A(n727), .ZN(n566) );
  XNOR2_X1 U480 ( .A(n481), .B(n480), .ZN(n484) );
  XNOR2_X1 U481 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U482 ( .A(n486), .B(n485), .ZN(n596) );
  XNOR2_X1 U483 ( .A(KEYINPUT35), .B(KEYINPUT82), .ZN(n564) );
  NAND2_X1 U484 ( .A1(n528), .A2(n537), .ZN(n682) );
  XNOR2_X1 U485 ( .A(n444), .B(KEYINPUT16), .ZN(n394) );
  INV_X1 U486 ( .A(G113), .ZN(n392) );
  XNOR2_X1 U487 ( .A(n393), .B(n392), .ZN(n481) );
  XNOR2_X1 U488 ( .A(n394), .B(n481), .ZN(n399) );
  XNOR2_X1 U489 ( .A(G110), .B(G107), .ZN(n395) );
  XNOR2_X1 U490 ( .A(n395), .B(KEYINPUT87), .ZN(n398) );
  INV_X1 U491 ( .A(KEYINPUT76), .ZN(n396) );
  XNOR2_X1 U492 ( .A(n396), .B(G104), .ZN(n397) );
  XNOR2_X1 U493 ( .A(n398), .B(n397), .ZN(n463) );
  XNOR2_X1 U494 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n400) );
  XNOR2_X1 U495 ( .A(n428), .B(n400), .ZN(n401) );
  XNOR2_X1 U496 ( .A(n401), .B(n440), .ZN(n406) );
  XNOR2_X1 U497 ( .A(n402), .B(G101), .ZN(n461) );
  NAND2_X1 U498 ( .A1(n715), .A2(G224), .ZN(n403) );
  XNOR2_X1 U499 ( .A(n403), .B(KEYINPUT4), .ZN(n404) );
  XNOR2_X1 U500 ( .A(n461), .B(n404), .ZN(n405) );
  XNOR2_X1 U501 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U502 ( .A(n701), .B(n407), .ZN(n611) );
  XNOR2_X1 U503 ( .A(KEYINPUT15), .B(G902), .ZN(n592) );
  INV_X1 U504 ( .A(n592), .ZN(n595) );
  OR2_X2 U505 ( .A1(n611), .A2(n595), .ZN(n411) );
  INV_X1 U506 ( .A(G902), .ZN(n487) );
  INV_X1 U507 ( .A(G237), .ZN(n408) );
  NAND2_X1 U508 ( .A1(n487), .A2(n408), .ZN(n412) );
  NAND2_X1 U509 ( .A1(n412), .A2(G210), .ZN(n409) );
  XNOR2_X1 U510 ( .A(n409), .B(KEYINPUT88), .ZN(n410) );
  NAND2_X1 U511 ( .A1(n412), .A2(G214), .ZN(n638) );
  INV_X1 U512 ( .A(n638), .ZN(n413) );
  NOR2_X2 U513 ( .A1(n506), .A2(n413), .ZN(n415) );
  XNOR2_X1 U514 ( .A(KEYINPUT68), .B(KEYINPUT19), .ZN(n416) );
  NAND2_X1 U515 ( .A1(G234), .A2(G237), .ZN(n417) );
  XNOR2_X1 U516 ( .A(n417), .B(KEYINPUT14), .ZN(n418) );
  XNOR2_X1 U517 ( .A(KEYINPUT74), .B(n418), .ZN(n420) );
  NAND2_X1 U518 ( .A1(G952), .A2(n420), .ZN(n653) );
  NOR2_X1 U519 ( .A1(n653), .A2(G953), .ZN(n656) );
  AND2_X1 U520 ( .A1(G953), .A2(G902), .ZN(n419) );
  NAND2_X1 U521 ( .A1(n420), .A2(n419), .ZN(n497) );
  NOR2_X1 U522 ( .A1(n497), .A2(G898), .ZN(n421) );
  NOR2_X1 U523 ( .A1(n656), .A2(n421), .ZN(n422) );
  INV_X1 U524 ( .A(KEYINPUT70), .ZN(n423) );
  XOR2_X1 U525 ( .A(G122), .B(G104), .Z(n426) );
  XNOR2_X1 U526 ( .A(n426), .B(n425), .ZN(n429) );
  INV_X1 U527 ( .A(KEYINPUT10), .ZN(n427) );
  XOR2_X1 U528 ( .A(n429), .B(n467), .Z(n436) );
  XOR2_X1 U529 ( .A(G140), .B(KEYINPUT12), .Z(n431) );
  NAND2_X1 U530 ( .A1(G214), .A2(n479), .ZN(n430) );
  XNOR2_X1 U531 ( .A(n431), .B(n430), .ZN(n434) );
  XOR2_X1 U532 ( .A(KEYINPUT11), .B(KEYINPUT94), .Z(n433) );
  XNOR2_X1 U533 ( .A(G131), .B(KEYINPUT93), .ZN(n432) );
  XNOR2_X1 U534 ( .A(n434), .B(n345), .ZN(n435) );
  XNOR2_X1 U535 ( .A(n436), .B(n435), .ZN(n604) );
  NOR2_X1 U536 ( .A1(G902), .A2(n604), .ZN(n439) );
  XNOR2_X1 U537 ( .A(KEYINPUT95), .B(KEYINPUT13), .ZN(n437) );
  XOR2_X1 U538 ( .A(KEYINPUT9), .B(KEYINPUT97), .Z(n442) );
  XNOR2_X1 U539 ( .A(G107), .B(KEYINPUT7), .ZN(n441) );
  XNOR2_X1 U540 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U541 ( .A(n460), .B(n443), .ZN(n449) );
  XOR2_X1 U542 ( .A(n444), .B(KEYINPUT96), .Z(n447) );
  NAND2_X1 U543 ( .A1(G234), .A2(n715), .ZN(n445) );
  XOR2_X1 U544 ( .A(KEYINPUT8), .B(n445), .Z(n469) );
  NAND2_X1 U545 ( .A1(G217), .A2(n469), .ZN(n446) );
  XNOR2_X1 U546 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U547 ( .A(n449), .B(n448), .ZN(n696) );
  NOR2_X1 U548 ( .A1(n696), .A2(G902), .ZN(n450) );
  XNOR2_X1 U549 ( .A(n450), .B(G478), .ZN(n537) );
  NAND2_X1 U550 ( .A1(n536), .A2(n537), .ZN(n642) );
  NAND2_X1 U551 ( .A1(n592), .A2(G234), .ZN(n452) );
  XNOR2_X1 U552 ( .A(KEYINPUT90), .B(KEYINPUT20), .ZN(n451) );
  XNOR2_X1 U553 ( .A(n452), .B(n451), .ZN(n474) );
  NAND2_X1 U554 ( .A1(n474), .A2(G221), .ZN(n453) );
  XNOR2_X1 U555 ( .A(n453), .B(KEYINPUT21), .ZN(n626) );
  NOR2_X1 U556 ( .A1(n642), .A2(n626), .ZN(n454) );
  NAND2_X1 U557 ( .A1(n559), .A2(n454), .ZN(n457) );
  INV_X1 U558 ( .A(KEYINPUT66), .ZN(n455) );
  XNOR2_X1 U559 ( .A(n455), .B(KEYINPUT22), .ZN(n456) );
  INV_X1 U560 ( .A(n493), .ZN(n490) );
  XOR2_X1 U561 ( .A(G137), .B(G140), .Z(n468) );
  NAND2_X1 U562 ( .A1(G227), .A2(n715), .ZN(n462) );
  XNOR2_X1 U563 ( .A(n468), .B(n462), .ZN(n464) );
  NOR2_X1 U564 ( .A1(n690), .A2(G902), .ZN(n465) );
  XNOR2_X1 U565 ( .A(KEYINPUT67), .B(KEYINPUT1), .ZN(n466) );
  XNOR2_X2 U566 ( .A(n516), .B(n466), .ZN(n556) );
  NAND2_X1 U567 ( .A1(n469), .A2(G221), .ZN(n470) );
  XNOR2_X1 U568 ( .A(n472), .B(n471), .ZN(n473) );
  NAND2_X1 U569 ( .A1(n619), .A2(n487), .ZN(n477) );
  NAND2_X1 U570 ( .A1(G217), .A2(n474), .ZN(n475) );
  XNOR2_X1 U571 ( .A(n475), .B(KEYINPUT25), .ZN(n476) );
  INV_X1 U572 ( .A(n625), .ZN(n500) );
  OR2_X1 U573 ( .A1(n556), .A2(n500), .ZN(n488) );
  INV_X1 U574 ( .A(n478), .ZN(n486) );
  NAND2_X1 U575 ( .A1(n479), .A2(G210), .ZN(n480) );
  XNOR2_X1 U576 ( .A(n482), .B(KEYINPUT5), .ZN(n483) );
  OR2_X1 U577 ( .A1(n488), .A2(n492), .ZN(n489) );
  OR2_X1 U578 ( .A1(n490), .A2(n489), .ZN(n581) );
  XNOR2_X1 U579 ( .A(G110), .B(KEYINPUT108), .ZN(n491) );
  XNOR2_X1 U580 ( .A(n581), .B(n491), .ZN(G12) );
  AND2_X1 U581 ( .A1(n556), .A2(n625), .ZN(n494) );
  INV_X1 U582 ( .A(KEYINPUT78), .ZN(n495) );
  XNOR2_X1 U583 ( .A(n495), .B(KEYINPUT32), .ZN(n496) );
  XOR2_X1 U584 ( .A(G119), .B(n582), .Z(G21) );
  XOR2_X1 U585 ( .A(KEYINPUT101), .B(KEYINPUT43), .Z(n505) );
  XNOR2_X1 U586 ( .A(KEYINPUT100), .B(n497), .ZN(n498) );
  NOR2_X1 U587 ( .A1(G900), .A2(n498), .ZN(n499) );
  NOR2_X1 U588 ( .A1(n656), .A2(n499), .ZN(n515) );
  OR2_X1 U589 ( .A1(n500), .A2(n626), .ZN(n501) );
  INV_X1 U590 ( .A(n536), .ZN(n528) );
  NAND2_X1 U591 ( .A1(n508), .A2(n502), .ZN(n523) );
  NOR2_X1 U592 ( .A1(n556), .A2(n523), .ZN(n503) );
  NAND2_X1 U593 ( .A1(n638), .A2(n503), .ZN(n504) );
  XNOR2_X1 U594 ( .A(n505), .B(n504), .ZN(n507) );
  NAND2_X1 U595 ( .A1(n507), .A2(n506), .ZN(n551) );
  XNOR2_X1 U596 ( .A(n551), .B(G140), .ZN(G42) );
  XNOR2_X1 U597 ( .A(KEYINPUT28), .B(n509), .ZN(n511) );
  INV_X1 U598 ( .A(n516), .ZN(n510) );
  NAND2_X1 U599 ( .A1(n511), .A2(n510), .ZN(n533) );
  XNOR2_X1 U600 ( .A(n506), .B(KEYINPUT38), .ZN(n639) );
  NAND2_X1 U601 ( .A1(n639), .A2(n638), .ZN(n643) );
  NOR2_X1 U602 ( .A1(n642), .A2(n643), .ZN(n513) );
  XOR2_X1 U603 ( .A(KEYINPUT41), .B(KEYINPUT103), .Z(n512) );
  XNOR2_X1 U604 ( .A(n513), .B(n512), .ZN(n661) );
  NOR2_X1 U605 ( .A1(n533), .A2(n661), .ZN(n514) );
  XNOR2_X1 U606 ( .A(n514), .B(KEYINPUT42), .ZN(n730) );
  INV_X1 U607 ( .A(n515), .ZN(n517) );
  NOR2_X1 U608 ( .A1(n625), .A2(n626), .ZN(n623) );
  NAND2_X1 U609 ( .A1(n623), .A2(n510), .ZN(n567) );
  INV_X1 U610 ( .A(n639), .ZN(n518) );
  NAND2_X1 U611 ( .A1(n492), .A2(n638), .ZN(n519) );
  XNOR2_X1 U612 ( .A(KEYINPUT30), .B(n519), .ZN(n535) );
  XNOR2_X1 U613 ( .A(n521), .B(n520), .ZN(n550) );
  INV_X1 U614 ( .A(n682), .ZN(n529) );
  XNOR2_X1 U615 ( .A(KEYINPUT104), .B(n523), .ZN(n526) );
  INV_X1 U616 ( .A(n524), .ZN(n525) );
  NOR2_X1 U617 ( .A1(n528), .A2(n537), .ZN(n671) );
  INV_X1 U618 ( .A(n573), .ZN(n644) );
  NAND2_X1 U619 ( .A1(n644), .A2(KEYINPUT47), .ZN(n531) );
  XOR2_X1 U620 ( .A(n531), .B(KEYINPUT79), .Z(n543) );
  NAND2_X1 U621 ( .A1(n680), .A2(KEYINPUT47), .ZN(n542) );
  OR2_X1 U622 ( .A1(n535), .A2(n534), .ZN(n540) );
  INV_X1 U623 ( .A(n506), .ZN(n538) );
  NOR2_X1 U624 ( .A1(n537), .A2(n536), .ZN(n562) );
  NAND2_X1 U625 ( .A1(n538), .A2(n562), .ZN(n539) );
  NOR2_X1 U626 ( .A1(n540), .A2(n539), .ZN(n679) );
  INV_X1 U627 ( .A(n679), .ZN(n541) );
  NOR2_X1 U628 ( .A1(n680), .A2(KEYINPUT47), .ZN(n544) );
  NAND2_X1 U629 ( .A1(n573), .A2(n544), .ZN(n545) );
  XNOR2_X1 U630 ( .A(n546), .B(KEYINPUT73), .ZN(n547) );
  XNOR2_X1 U631 ( .A(n549), .B(KEYINPUT48), .ZN(n553) );
  NAND2_X1 U632 ( .A1(n550), .A2(n671), .ZN(n688) );
  AND2_X1 U633 ( .A1(n551), .A2(n688), .ZN(n552) );
  INV_X1 U634 ( .A(KEYINPUT44), .ZN(n585) );
  NAND2_X1 U635 ( .A1(n581), .A2(n585), .ZN(n554) );
  NAND2_X1 U636 ( .A1(n556), .A2(n623), .ZN(n557) );
  XNOR2_X1 U637 ( .A(n346), .B(KEYINPUT33), .ZN(n662) );
  INV_X1 U638 ( .A(n570), .ZN(n560) );
  XNOR2_X1 U639 ( .A(n561), .B(KEYINPUT34), .ZN(n563) );
  NAND2_X1 U640 ( .A1(n563), .A2(n562), .ZN(n565) );
  XNOR2_X2 U641 ( .A(n565), .B(n564), .ZN(n727) );
  NAND2_X1 U642 ( .A1(n391), .A2(n566), .ZN(n580) );
  NOR2_X1 U643 ( .A1(n492), .A2(n567), .ZN(n568) );
  NAND2_X1 U644 ( .A1(n568), .A2(n570), .ZN(n672) );
  NAND2_X1 U645 ( .A1(n635), .A2(n570), .ZN(n572) );
  XOR2_X1 U646 ( .A(KEYINPUT31), .B(KEYINPUT92), .Z(n571) );
  XNOR2_X1 U647 ( .A(n572), .B(n571), .ZN(n686) );
  NAND2_X1 U648 ( .A1(n672), .A2(n686), .ZN(n574) );
  NAND2_X1 U649 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U650 ( .A(n575), .B(KEYINPUT99), .ZN(n578) );
  NOR2_X1 U651 ( .A1(n556), .A2(n625), .ZN(n576) );
  AND2_X1 U652 ( .A1(n577), .A2(n576), .ZN(n668) );
  NOR2_X1 U653 ( .A1(n578), .A2(n668), .ZN(n579) );
  NAND2_X1 U654 ( .A1(n727), .A2(KEYINPUT84), .ZN(n584) );
  NOR2_X1 U655 ( .A1(n582), .A2(n388), .ZN(n583) );
  NAND2_X1 U656 ( .A1(n584), .A2(n583), .ZN(n587) );
  NAND2_X1 U657 ( .A1(n585), .A2(KEYINPUT84), .ZN(n586) );
  NAND2_X1 U658 ( .A1(n587), .A2(n586), .ZN(n588) );
  INV_X1 U659 ( .A(KEYINPUT77), .ZN(n591) );
  XNOR2_X1 U660 ( .A(n592), .B(KEYINPUT81), .ZN(n593) );
  XOR2_X1 U661 ( .A(KEYINPUT77), .B(KEYINPUT2), .Z(n594) );
  NAND2_X1 U662 ( .A1(n617), .A2(G472), .ZN(n598) );
  XOR2_X1 U663 ( .A(KEYINPUT62), .B(n596), .Z(n597) );
  XNOR2_X1 U664 ( .A(n598), .B(n597), .ZN(n600) );
  INV_X1 U665 ( .A(G952), .ZN(n599) );
  NOR2_X2 U666 ( .A1(n600), .A2(n700), .ZN(n603) );
  XNOR2_X1 U667 ( .A(KEYINPUT106), .B(KEYINPUT63), .ZN(n601) );
  XOR2_X1 U668 ( .A(n601), .B(KEYINPUT86), .Z(n602) );
  XNOR2_X1 U669 ( .A(n603), .B(n602), .ZN(G57) );
  NAND2_X1 U670 ( .A1(n617), .A2(G475), .ZN(n606) );
  XOR2_X1 U671 ( .A(KEYINPUT59), .B(n604), .Z(n605) );
  XNOR2_X1 U672 ( .A(n606), .B(n605), .ZN(n607) );
  NOR2_X2 U673 ( .A1(n607), .A2(n700), .ZN(n609) );
  XOR2_X1 U674 ( .A(KEYINPUT69), .B(KEYINPUT60), .Z(n608) );
  XNOR2_X1 U675 ( .A(n609), .B(n608), .ZN(G60) );
  NAND2_X1 U676 ( .A1(n617), .A2(G210), .ZN(n613) );
  XOR2_X1 U677 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n610) );
  XNOR2_X1 U678 ( .A(n611), .B(n610), .ZN(n612) );
  XNOR2_X1 U679 ( .A(n613), .B(n612), .ZN(n614) );
  NOR2_X2 U680 ( .A1(n614), .A2(n700), .ZN(n616) );
  XOR2_X1 U681 ( .A(KEYINPUT83), .B(KEYINPUT56), .Z(n615) );
  XNOR2_X1 U682 ( .A(n616), .B(n615), .ZN(G51) );
  NAND2_X1 U683 ( .A1(n617), .A2(G217), .ZN(n621) );
  XNOR2_X1 U684 ( .A(KEYINPUT122), .B(KEYINPUT123), .ZN(n618) );
  XNOR2_X1 U685 ( .A(n619), .B(n618), .ZN(n620) );
  XNOR2_X1 U686 ( .A(n621), .B(n620), .ZN(n622) );
  NOR2_X1 U687 ( .A1(n622), .A2(n700), .ZN(G66) );
  XNOR2_X1 U688 ( .A(KEYINPUT52), .B(KEYINPUT118), .ZN(n652) );
  NOR2_X1 U689 ( .A1(n623), .A2(n556), .ZN(n624) );
  XNOR2_X1 U690 ( .A(KEYINPUT50), .B(n624), .ZN(n633) );
  XOR2_X1 U691 ( .A(KEYINPUT49), .B(KEYINPUT114), .Z(n628) );
  NAND2_X1 U692 ( .A1(n626), .A2(n625), .ZN(n627) );
  XNOR2_X1 U693 ( .A(n628), .B(n627), .ZN(n629) );
  XNOR2_X1 U694 ( .A(n629), .B(KEYINPUT113), .ZN(n630) );
  NOR2_X1 U695 ( .A1(n492), .A2(n630), .ZN(n631) );
  XNOR2_X1 U696 ( .A(KEYINPUT115), .B(n631), .ZN(n632) );
  NOR2_X1 U697 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U698 ( .A1(n635), .A2(n634), .ZN(n636) );
  XOR2_X1 U699 ( .A(KEYINPUT51), .B(n636), .Z(n637) );
  NOR2_X1 U700 ( .A1(n661), .A2(n637), .ZN(n650) );
  NOR2_X1 U701 ( .A1(n639), .A2(n638), .ZN(n640) );
  XNOR2_X1 U702 ( .A(n640), .B(KEYINPUT116), .ZN(n641) );
  NOR2_X1 U703 ( .A1(n642), .A2(n641), .ZN(n646) );
  NOR2_X1 U704 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U705 ( .A1(n646), .A2(n645), .ZN(n647) );
  XOR2_X1 U706 ( .A(KEYINPUT117), .B(n647), .Z(n648) );
  NOR2_X1 U707 ( .A1(n662), .A2(n648), .ZN(n649) );
  NOR2_X1 U708 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U709 ( .A(n652), .B(n651), .ZN(n658) );
  NOR2_X1 U710 ( .A1(n658), .A2(n653), .ZN(n655) );
  OR2_X1 U711 ( .A1(G953), .A2(KEYINPUT119), .ZN(n654) );
  NOR2_X1 U712 ( .A1(n655), .A2(n654), .ZN(n660) );
  NAND2_X1 U713 ( .A1(n656), .A2(KEYINPUT119), .ZN(n657) );
  NOR2_X1 U714 ( .A1(n658), .A2(n657), .ZN(n659) );
  NOR2_X1 U715 ( .A1(n660), .A2(n659), .ZN(n664) );
  NOR2_X1 U716 ( .A1(n662), .A2(n661), .ZN(n663) );
  NOR2_X1 U717 ( .A1(n664), .A2(n663), .ZN(n665) );
  NAND2_X1 U718 ( .A1(n666), .A2(n665), .ZN(n667) );
  XOR2_X1 U719 ( .A(G101), .B(n668), .Z(G3) );
  NOR2_X1 U720 ( .A1(n682), .A2(n672), .ZN(n670) );
  XNOR2_X1 U721 ( .A(G104), .B(KEYINPUT107), .ZN(n669) );
  XNOR2_X1 U722 ( .A(n670), .B(n669), .ZN(G6) );
  INV_X1 U723 ( .A(n671), .ZN(n685) );
  NOR2_X1 U724 ( .A1(n685), .A2(n672), .ZN(n674) );
  XNOR2_X1 U725 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n673) );
  XNOR2_X1 U726 ( .A(n674), .B(n673), .ZN(n675) );
  XNOR2_X1 U727 ( .A(G107), .B(n675), .ZN(G9) );
  NOR2_X1 U728 ( .A1(n680), .A2(n685), .ZN(n677) );
  XNOR2_X1 U729 ( .A(KEYINPUT109), .B(KEYINPUT29), .ZN(n676) );
  XNOR2_X1 U730 ( .A(n677), .B(n676), .ZN(n678) );
  XOR2_X1 U731 ( .A(G128), .B(n678), .Z(G30) );
  XOR2_X1 U732 ( .A(G143), .B(n679), .Z(G45) );
  NOR2_X1 U733 ( .A1(n680), .A2(n682), .ZN(n681) );
  XOR2_X1 U734 ( .A(G146), .B(n681), .Z(G48) );
  NOR2_X1 U735 ( .A1(n686), .A2(n682), .ZN(n683) );
  XOR2_X1 U736 ( .A(KEYINPUT110), .B(n683), .Z(n684) );
  XNOR2_X1 U737 ( .A(G113), .B(n684), .ZN(G15) );
  NOR2_X1 U738 ( .A1(n686), .A2(n685), .ZN(n687) );
  XOR2_X1 U739 ( .A(G116), .B(n687), .Z(G18) );
  XNOR2_X1 U740 ( .A(G134), .B(KEYINPUT112), .ZN(n689) );
  XNOR2_X1 U741 ( .A(n689), .B(n688), .ZN(G36) );
  NAND2_X1 U742 ( .A1(n617), .A2(G469), .ZN(n694) );
  XOR2_X1 U743 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n692) );
  XNOR2_X1 U744 ( .A(n690), .B(KEYINPUT120), .ZN(n691) );
  XNOR2_X1 U745 ( .A(n692), .B(n691), .ZN(n693) );
  XNOR2_X1 U746 ( .A(n694), .B(n693), .ZN(n695) );
  NOR2_X1 U747 ( .A1(n700), .A2(n695), .ZN(G54) );
  NAND2_X1 U748 ( .A1(n617), .A2(G478), .ZN(n698) );
  XOR2_X1 U749 ( .A(n696), .B(KEYINPUT121), .Z(n697) );
  XNOR2_X1 U750 ( .A(n698), .B(n697), .ZN(n699) );
  NOR2_X1 U751 ( .A1(n700), .A2(n699), .ZN(G63) );
  XNOR2_X1 U752 ( .A(n701), .B(G101), .ZN(n703) );
  NOR2_X1 U753 ( .A1(G898), .A2(n715), .ZN(n702) );
  NOR2_X1 U754 ( .A1(n703), .A2(n702), .ZN(n704) );
  XOR2_X1 U755 ( .A(KEYINPUT124), .B(n704), .Z(n711) );
  NAND2_X1 U756 ( .A1(n705), .A2(n715), .ZN(n709) );
  NAND2_X1 U757 ( .A1(G953), .A2(G224), .ZN(n706) );
  XNOR2_X1 U758 ( .A(KEYINPUT61), .B(n706), .ZN(n707) );
  NAND2_X1 U759 ( .A1(n707), .A2(G898), .ZN(n708) );
  NAND2_X1 U760 ( .A1(n709), .A2(n708), .ZN(n710) );
  XOR2_X1 U761 ( .A(n711), .B(n710), .Z(G69) );
  XNOR2_X1 U762 ( .A(n713), .B(n712), .ZN(n717) );
  XNOR2_X1 U763 ( .A(n714), .B(n717), .ZN(n716) );
  NAND2_X1 U764 ( .A1(n716), .A2(n715), .ZN(n722) );
  XNOR2_X1 U765 ( .A(n717), .B(G227), .ZN(n718) );
  XNOR2_X1 U766 ( .A(n718), .B(KEYINPUT125), .ZN(n719) );
  NAND2_X1 U767 ( .A1(n719), .A2(G900), .ZN(n720) );
  NAND2_X1 U768 ( .A1(G953), .A2(n720), .ZN(n721) );
  NAND2_X1 U769 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U770 ( .A(KEYINPUT126), .B(n723), .ZN(G72) );
  XOR2_X1 U771 ( .A(KEYINPUT37), .B(KEYINPUT111), .Z(n726) );
  XNOR2_X1 U772 ( .A(G125), .B(n724), .ZN(n725) );
  XNOR2_X1 U773 ( .A(n726), .B(n725), .ZN(G27) );
  XNOR2_X1 U774 ( .A(G122), .B(KEYINPUT127), .ZN(n728) );
  XNOR2_X1 U775 ( .A(n728), .B(n727), .ZN(G24) );
  XOR2_X1 U776 ( .A(n729), .B(G131), .Z(G33) );
  XOR2_X1 U777 ( .A(G137), .B(n730), .Z(G39) );
endmodule

