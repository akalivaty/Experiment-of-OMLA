//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 0 1 1 1 1 1 0 1 1 1 0 1 1 1 0 1 1 1 1 0 0 0 0 1 0 0 1 0 1 0 1 1 1 0 1 0 1 1 1 0 0 0 0 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:56 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n448, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n556, new_n558, new_n559, new_n560,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n605, new_n608, new_n610, new_n611, new_n612,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n821, new_n822,
    new_n823, new_n824, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1158, new_n1159, new_n1160,
    new_n1162, new_n1163, new_n1164, new_n1165;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT65), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT66), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT67), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT68), .Z(new_n456));
  NAND2_X1  g031(.A1(new_n454), .A2(new_n456), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(new_n454), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G2106), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT69), .ZN(new_n461));
  INV_X1    g036(.A(new_n456), .ZN(new_n462));
  AOI21_X1  g037(.A(new_n461), .B1(G567), .B2(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  AND2_X1   g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G125), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n464), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(G101), .A2(G2104), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT70), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n474), .B1(new_n465), .B2(KEYINPUT3), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n467), .A2(KEYINPUT70), .A3(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(new_n466), .ZN(new_n478));
  INV_X1    g053(.A(G137), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n473), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n472), .B1(new_n464), .B2(new_n480), .ZN(G160));
  NOR2_X1   g056(.A1(new_n478), .A2(new_n464), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n478), .A2(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n483), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  XNOR2_X1  g063(.A(new_n488), .B(KEYINPUT71), .ZN(G162));
  NAND4_X1  g064(.A1(new_n477), .A2(G126), .A3(G2105), .A4(new_n466), .ZN(new_n490));
  AND2_X1   g065(.A1(KEYINPUT4), .A2(G138), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n477), .A2(new_n464), .A3(new_n466), .A4(new_n491), .ZN(new_n492));
  OR2_X1    g067(.A1(G102), .A2(G2105), .ZN(new_n493));
  XNOR2_X1  g068(.A(KEYINPUT72), .B(G114), .ZN(new_n494));
  OAI211_X1 g069(.A(G2104), .B(new_n493), .C1(new_n494), .C2(new_n464), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n466), .A2(new_n468), .A3(G138), .A4(new_n464), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n490), .A2(new_n492), .A3(new_n495), .A4(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT5), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G62), .ZN(new_n506));
  OR3_X1    g081(.A1(new_n505), .A2(KEYINPUT74), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(G75), .A2(G543), .ZN(new_n508));
  OAI21_X1  g083(.A(KEYINPUT74), .B1(new_n505), .B2(new_n506), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G651), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT6), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G651), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  AND3_X1   g089(.A1(new_n514), .A2(KEYINPUT73), .A3(KEYINPUT6), .ZN(new_n515));
  AOI21_X1  g090(.A(KEYINPUT73), .B1(new_n514), .B2(KEYINPUT6), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n513), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n517), .A2(new_n501), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n517), .A2(new_n505), .ZN(new_n519));
  AOI22_X1  g094(.A1(G50), .A2(new_n518), .B1(new_n519), .B2(G88), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n511), .A2(new_n520), .ZN(G303));
  INV_X1    g096(.A(G303), .ZN(G166));
  NAND2_X1  g097(.A1(G63), .A2(G651), .ZN(new_n523));
  INV_X1    g098(.A(G89), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n523), .B1(new_n517), .B2(new_n524), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n502), .A2(new_n504), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n525), .A2(new_n526), .B1(new_n518), .B2(G51), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT7), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n527), .A2(new_n529), .ZN(G286));
  INV_X1    g105(.A(G286), .ZN(G168));
  AOI22_X1  g106(.A1(new_n526), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n532));
  OR2_X1    g107(.A1(new_n532), .A2(new_n514), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n519), .A2(G90), .ZN(new_n534));
  XNOR2_X1  g109(.A(KEYINPUT75), .B(G52), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n518), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n533), .A2(new_n534), .A3(new_n536), .ZN(G301));
  INV_X1    g112(.A(G301), .ZN(G171));
  AOI22_X1  g113(.A1(new_n526), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n539), .A2(new_n514), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT73), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n541), .B1(new_n512), .B2(G651), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n514), .A2(KEYINPUT73), .A3(KEYINPUT6), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n542), .A2(new_n543), .B1(new_n512), .B2(G651), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n544), .A2(G43), .A3(G543), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n544), .A2(G81), .A3(new_n526), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT76), .ZN(new_n547));
  AND3_X1   g122(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n547), .B1(new_n545), .B2(new_n546), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n540), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT77), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  OAI211_X1 g127(.A(KEYINPUT77), .B(new_n540), .C1(new_n548), .C2(new_n549), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  AND3_X1   g130(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G36), .ZN(G176));
  XOR2_X1   g132(.A(KEYINPUT78), .B(KEYINPUT8), .Z(new_n558));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n558), .B(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n556), .A2(new_n560), .ZN(G188));
  XNOR2_X1  g136(.A(new_n526), .B(KEYINPUT79), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G65), .ZN(new_n563));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G651), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n518), .A2(G53), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT9), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n518), .A2(KEYINPUT9), .A3(G53), .ZN(new_n570));
  AND2_X1   g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n519), .A2(G91), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n566), .A2(new_n571), .A3(new_n572), .ZN(G299));
  NAND2_X1  g148(.A1(new_n518), .A2(G49), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n519), .A2(G87), .ZN(new_n575));
  OAI21_X1  g150(.A(G651), .B1(new_n526), .B2(G74), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(G288));
  AND2_X1   g152(.A1(G48), .A2(G543), .ZN(new_n578));
  OAI211_X1 g153(.A(new_n513), .B(new_n578), .C1(new_n515), .C2(new_n516), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT80), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n544), .A2(KEYINPUT80), .A3(new_n578), .ZN(new_n582));
  AND2_X1   g157(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n526), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n584));
  OR2_X1    g159(.A1(new_n584), .A2(new_n514), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n544), .A2(G86), .A3(new_n526), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n583), .A2(new_n585), .A3(new_n586), .ZN(G305));
  AOI22_X1  g162(.A1(new_n526), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n588));
  OR2_X1    g163(.A1(new_n588), .A2(new_n514), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n519), .A2(G85), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n518), .A2(G47), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(G290));
  NAND2_X1  g167(.A1(G301), .A2(G868), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n562), .A2(G66), .ZN(new_n594));
  NAND2_X1  g169(.A1(G79), .A2(G543), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n596), .A2(G651), .B1(G54), .B2(new_n518), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n519), .A2(G92), .ZN(new_n598));
  XOR2_X1   g173(.A(new_n598), .B(KEYINPUT10), .Z(new_n599));
  NAND2_X1  g174(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n593), .B1(new_n601), .B2(G868), .ZN(G284));
  XNOR2_X1  g177(.A(G284), .B(KEYINPUT81), .ZN(G321));
  NAND2_X1  g178(.A1(G286), .A2(G868), .ZN(new_n604));
  INV_X1    g179(.A(G299), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n605), .B2(G868), .ZN(G297));
  XNOR2_X1  g181(.A(G297), .B(KEYINPUT82), .ZN(G280));
  INV_X1    g182(.A(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n601), .B1(new_n608), .B2(G860), .ZN(G148));
  INV_X1    g184(.A(G868), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n552), .A2(new_n610), .A3(new_n553), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n600), .A2(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n612), .B2(new_n610), .ZN(G323));
  XNOR2_X1  g188(.A(KEYINPUT83), .B(KEYINPUT11), .ZN(new_n614));
  XNOR2_X1  g189(.A(G323), .B(new_n614), .ZN(G282));
  NAND2_X1  g190(.A1(new_n482), .A2(G123), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT85), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n484), .A2(G135), .ZN(new_n619));
  OR2_X1    g194(.A1(G99), .A2(G2105), .ZN(new_n620));
  OAI211_X1 g195(.A(new_n620), .B(G2104), .C1(G111), .C2(new_n464), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n482), .A2(KEYINPUT85), .A3(G123), .ZN(new_n622));
  NAND4_X1  g197(.A1(new_n618), .A2(new_n619), .A3(new_n621), .A4(new_n622), .ZN(new_n623));
  INV_X1    g198(.A(G2096), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g200(.A(KEYINPUT84), .B(KEYINPUT12), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n464), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT13), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(G2100), .Z(new_n630));
  NAND2_X1  g205(.A1(new_n625), .A2(new_n630), .ZN(G156));
  XNOR2_X1  g206(.A(KEYINPUT15), .B(G2430), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2435), .ZN(new_n633));
  XOR2_X1   g208(.A(G2427), .B(G2438), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n635), .A2(KEYINPUT14), .ZN(new_n636));
  XOR2_X1   g211(.A(G2451), .B(G2454), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT16), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n636), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2443), .B(G2446), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(G1341), .B(G1348), .Z(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(KEYINPUT86), .Z(new_n644));
  OAI21_X1  g219(.A(G14), .B1(new_n641), .B2(new_n642), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n644), .A2(new_n645), .ZN(G401));
  XNOR2_X1  g221(.A(G2072), .B(G2078), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT87), .ZN(new_n648));
  XOR2_X1   g223(.A(G2084), .B(G2090), .Z(new_n649));
  XOR2_X1   g224(.A(G2067), .B(G2678), .Z(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n648), .A2(new_n649), .A3(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(KEYINPUT18), .Z(new_n653));
  INV_X1    g228(.A(new_n649), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n654), .A2(new_n650), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n648), .A2(KEYINPUT17), .A3(new_n655), .ZN(new_n656));
  AND2_X1   g231(.A1(new_n655), .A2(KEYINPUT17), .ZN(new_n657));
  OAI221_X1 g232(.A(new_n656), .B1(new_n654), .B2(new_n650), .C1(new_n657), .C2(new_n648), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n653), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(new_n624), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G2100), .ZN(G227));
  XNOR2_X1  g236(.A(G1971), .B(G1976), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT88), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT19), .ZN(new_n664));
  XOR2_X1   g239(.A(G1956), .B(G2474), .Z(new_n665));
  XOR2_X1   g240(.A(G1961), .B(G1966), .Z(new_n666));
  AND2_X1   g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT20), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n665), .A2(new_n666), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n664), .A2(new_n670), .ZN(new_n671));
  OR3_X1    g246(.A1(new_n664), .A2(new_n667), .A3(new_n670), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n669), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(KEYINPUT21), .B(G1986), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G1991), .B(G1996), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT22), .B(G1981), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n677), .B(new_n678), .Z(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(G229));
  NOR2_X1   g255(.A1(G29), .A2(G35), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n681), .B1(G162), .B2(G29), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT29), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n683), .A2(G2090), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(KEYINPUT99), .Z(new_n685));
  INV_X1    g260(.A(G16), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(G19), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n687), .B1(new_n554), .B2(new_n686), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n686), .A2(G22), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n689), .B1(G166), .B2(new_n686), .ZN(new_n690));
  INV_X1    g265(.A(G1971), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  MUX2_X1   g267(.A(G6), .B(G305), .S(G16), .Z(new_n693));
  XOR2_X1   g268(.A(KEYINPUT32), .B(G1981), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  NOR2_X1   g270(.A1(G16), .A2(G23), .ZN(new_n696));
  INV_X1    g271(.A(G288), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n696), .B1(new_n697), .B2(G16), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT33), .B(G1976), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n692), .A2(new_n695), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(KEYINPUT34), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n686), .A2(G24), .ZN(new_n703));
  INV_X1    g278(.A(G290), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n703), .B1(new_n704), .B2(new_n686), .ZN(new_n705));
  MUX2_X1   g280(.A(new_n703), .B(new_n705), .S(KEYINPUT91), .Z(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT92), .B(G1986), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(KEYINPUT34), .ZN(new_n709));
  NAND4_X1  g284(.A1(new_n692), .A2(new_n695), .A3(new_n709), .A4(new_n700), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT89), .ZN(new_n711));
  AND2_X1   g286(.A1(new_n477), .A2(new_n466), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(new_n464), .ZN(new_n713));
  INV_X1    g288(.A(G131), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n711), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n482), .A2(G119), .ZN(new_n716));
  OR2_X1    g291(.A1(G95), .A2(G2105), .ZN(new_n717));
  OAI211_X1 g292(.A(new_n717), .B(G2104), .C1(G107), .C2(new_n464), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n484), .A2(KEYINPUT89), .A3(G131), .ZN(new_n719));
  NAND4_X1  g294(.A1(new_n715), .A2(new_n716), .A3(new_n718), .A4(new_n719), .ZN(new_n720));
  MUX2_X1   g295(.A(G25), .B(new_n720), .S(G29), .Z(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT35), .B(G1991), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(KEYINPUT90), .Z(new_n723));
  XNOR2_X1  g298(.A(new_n721), .B(new_n723), .ZN(new_n724));
  NAND4_X1  g299(.A1(new_n702), .A2(new_n708), .A3(new_n710), .A4(new_n724), .ZN(new_n725));
  AND2_X1   g300(.A1(new_n725), .A2(KEYINPUT36), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n725), .A2(KEYINPUT36), .ZN(new_n727));
  OAI221_X1 g302(.A(new_n685), .B1(G1341), .B2(new_n688), .C1(new_n726), .C2(new_n727), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n686), .A2(KEYINPUT23), .A3(G20), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT23), .ZN(new_n730));
  INV_X1    g305(.A(G20), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n730), .B1(new_n731), .B2(G16), .ZN(new_n732));
  OAI211_X1 g307(.A(new_n729), .B(new_n732), .C1(new_n605), .C2(new_n686), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(G1956), .ZN(new_n734));
  NAND2_X1  g309(.A1(G171), .A2(G16), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G5), .B2(G16), .ZN(new_n736));
  INV_X1    g311(.A(G1961), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(G29), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n623), .A2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT30), .ZN(new_n741));
  AND2_X1   g316(.A1(new_n741), .A2(G28), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n741), .A2(G28), .ZN(new_n743));
  NOR3_X1   g318(.A1(new_n742), .A2(new_n743), .A3(G29), .ZN(new_n744));
  NOR3_X1   g319(.A1(new_n738), .A2(new_n740), .A3(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(G34), .ZN(new_n746));
  AND2_X1   g321(.A1(new_n746), .A2(KEYINPUT24), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n746), .A2(KEYINPUT24), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n739), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G160), .B2(new_n739), .ZN(new_n750));
  INV_X1    g325(.A(G2084), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  XOR2_X1   g327(.A(KEYINPUT31), .B(G11), .Z(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(new_n736), .B2(new_n737), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n745), .A2(new_n752), .A3(new_n754), .ZN(new_n755));
  NOR3_X1   g330(.A1(new_n728), .A2(new_n734), .A3(new_n755), .ZN(new_n756));
  AOI22_X1  g331(.A1(new_n712), .A2(G141), .B1(G105), .B2(G2104), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n757), .A2(G2105), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(G129), .B2(new_n482), .ZN(new_n759));
  XOR2_X1   g334(.A(KEYINPUT96), .B(KEYINPUT26), .Z(new_n760));
  NAND3_X1  g335(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n759), .A2(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n764), .A2(G29), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G29), .B2(G32), .ZN(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT27), .B(G1996), .ZN(new_n767));
  OR2_X1    g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n686), .A2(G21), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G168), .B2(new_n686), .ZN(new_n770));
  INV_X1    g345(.A(G1966), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n739), .A2(G27), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G164), .B2(new_n739), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT98), .Z(new_n775));
  AND2_X1   g350(.A1(new_n775), .A2(G2078), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n775), .A2(G2078), .ZN(new_n777));
  INV_X1    g352(.A(G2072), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n469), .A2(G127), .ZN(new_n779));
  NAND2_X1  g354(.A1(G115), .A2(G2104), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n464), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND3_X1  g356(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT25), .ZN(new_n783));
  INV_X1    g358(.A(G139), .ZN(new_n784));
  OAI21_X1  g359(.A(KEYINPUT95), .B1(new_n713), .B2(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT95), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n484), .A2(new_n786), .A3(G139), .ZN(new_n787));
  AOI211_X1 g362(.A(new_n781), .B(new_n783), .C1(new_n785), .C2(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n788), .A2(new_n739), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(new_n739), .B2(G33), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n777), .B1(new_n778), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(new_n778), .B2(new_n790), .ZN(new_n792));
  AOI211_X1 g367(.A(new_n776), .B(new_n792), .C1(G1341), .C2(new_n688), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n739), .A2(G26), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n482), .A2(G128), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n484), .A2(G140), .ZN(new_n796));
  NOR2_X1   g371(.A1(G104), .A2(G2105), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT93), .Z(new_n798));
  OAI211_X1 g373(.A(new_n798), .B(G2104), .C1(G116), .C2(new_n464), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n795), .A2(new_n796), .A3(new_n799), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n800), .A2(KEYINPUT94), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(KEYINPUT94), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(new_n803), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n794), .B1(new_n804), .B2(new_n739), .ZN(new_n805));
  MUX2_X1   g380(.A(new_n794), .B(new_n805), .S(KEYINPUT28), .Z(new_n806));
  INV_X1    g381(.A(G2067), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n686), .A2(G4), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(new_n601), .B2(new_n686), .ZN(new_n810));
  INV_X1    g385(.A(G1348), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n683), .A2(G2090), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT97), .ZN(new_n814));
  AND3_X1   g389(.A1(new_n766), .A2(new_n814), .A3(new_n767), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n814), .B1(new_n766), .B2(new_n767), .ZN(new_n816));
  NOR3_X1   g391(.A1(new_n813), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  NAND4_X1  g392(.A1(new_n793), .A2(new_n808), .A3(new_n812), .A4(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  NAND4_X1  g394(.A1(new_n756), .A2(new_n768), .A3(new_n772), .A4(new_n819), .ZN(G150));
  NAND2_X1  g395(.A1(G150), .A2(KEYINPUT100), .ZN(new_n821));
  NOR4_X1   g396(.A1(new_n728), .A2(new_n818), .A3(new_n734), .A4(new_n755), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT100), .ZN(new_n823));
  NAND4_X1  g398(.A1(new_n822), .A2(new_n823), .A3(new_n768), .A4(new_n772), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n821), .A2(new_n824), .ZN(G311));
  AOI22_X1  g400(.A1(new_n526), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n826));
  OR2_X1    g401(.A1(new_n826), .A2(new_n514), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n519), .A2(G93), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n518), .A2(G55), .ZN(new_n829));
  AND3_X1   g404(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(G860), .ZN(new_n832));
  XOR2_X1   g407(.A(KEYINPUT104), .B(KEYINPUT37), .Z(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n554), .A2(new_n831), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT102), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n836), .B1(new_n830), .B2(new_n550), .ZN(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n830), .A2(new_n550), .A3(new_n836), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n835), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT103), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n830), .B1(new_n552), .B2(new_n553), .ZN(new_n843));
  INV_X1    g418(.A(new_n839), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n845), .A2(KEYINPUT103), .A3(new_n838), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n842), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n601), .A2(G559), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n847), .B(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT39), .ZN(new_n850));
  XNOR2_X1  g425(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n850), .B(new_n851), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n834), .B1(new_n852), .B2(G860), .ZN(G145));
  XNOR2_X1  g428(.A(new_n623), .B(G160), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n854), .B(G162), .Z(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT106), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n788), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n492), .A2(new_n498), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n490), .A2(new_n495), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(KEYINPUT105), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT105), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n490), .A2(new_n495), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n859), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n858), .B(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n803), .B(new_n720), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n865), .B(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(G142), .ZN(new_n868));
  OR3_X1    g443(.A1(new_n713), .A2(KEYINPUT107), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n482), .A2(G130), .ZN(new_n870));
  OR2_X1    g445(.A1(G106), .A2(G2105), .ZN(new_n871));
  OAI211_X1 g446(.A(new_n871), .B(G2104), .C1(G118), .C2(new_n464), .ZN(new_n872));
  OAI21_X1  g447(.A(KEYINPUT107), .B1(new_n713), .B2(new_n868), .ZN(new_n873));
  NAND4_X1  g448(.A1(new_n869), .A2(new_n870), .A3(new_n872), .A4(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(new_n628), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(new_n763), .ZN(new_n876));
  AND2_X1   g451(.A1(new_n867), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n867), .A2(new_n876), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n856), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(KEYINPUT108), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n877), .A2(new_n878), .ZN(new_n881));
  AOI21_X1  g456(.A(G37), .B1(new_n881), .B2(new_n855), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g459(.A(KEYINPUT112), .ZN(new_n885));
  OR2_X1    g460(.A1(new_n847), .A2(new_n612), .ZN(new_n886));
  AND2_X1   g461(.A1(new_n566), .A2(new_n571), .ZN(new_n887));
  NAND4_X1  g462(.A1(new_n887), .A2(new_n572), .A3(new_n597), .A4(new_n599), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n600), .A2(G299), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NOR3_X1   g465(.A1(new_n890), .A2(KEYINPUT109), .A3(KEYINPUT41), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT41), .ZN(new_n892));
  AND3_X1   g467(.A1(new_n888), .A2(new_n889), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n892), .B1(new_n888), .B2(new_n889), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n891), .B1(new_n895), .B2(KEYINPUT109), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n847), .A2(new_n612), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n886), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT110), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n886), .A2(new_n897), .ZN(new_n901));
  INV_X1    g476(.A(new_n890), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(KEYINPUT110), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n900), .B1(new_n904), .B2(new_n898), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n697), .B(G303), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n906), .B(G305), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n907), .B(G290), .ZN(new_n908));
  XOR2_X1   g483(.A(new_n908), .B(KEYINPUT42), .Z(new_n909));
  OAI21_X1  g484(.A(new_n885), .B1(new_n905), .B2(new_n909), .ZN(new_n910));
  AND3_X1   g485(.A1(new_n886), .A2(new_n896), .A3(new_n897), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(KEYINPUT110), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n899), .B1(new_n901), .B2(new_n902), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n912), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n909), .ZN(new_n915));
  OAI21_X1  g490(.A(KEYINPUT111), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT111), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n905), .A2(new_n917), .A3(new_n909), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n914), .A2(KEYINPUT112), .A3(new_n915), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n910), .A2(new_n916), .A3(new_n918), .A4(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(G868), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n831), .A2(new_n610), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(G295));
  NAND2_X1  g498(.A1(new_n921), .A2(new_n922), .ZN(G331));
  INV_X1    g499(.A(KEYINPUT43), .ZN(new_n925));
  XNOR2_X1  g500(.A(G286), .B(G301), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(KEYINPUT103), .B1(new_n845), .B2(new_n838), .ZN(new_n928));
  NOR4_X1   g503(.A1(new_n843), .A2(new_n844), .A3(new_n841), .A4(new_n837), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n927), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n842), .A2(new_n846), .A3(new_n926), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT113), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n847), .A2(KEYINPUT113), .A3(new_n927), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n896), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n908), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n930), .A2(new_n931), .A3(new_n902), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(G37), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n890), .B1(new_n933), .B2(new_n934), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n895), .B1(new_n930), .B2(new_n931), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n908), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(KEYINPUT114), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT114), .ZN(new_n945));
  OAI211_X1 g520(.A(new_n945), .B(new_n908), .C1(new_n941), .C2(new_n942), .ZN(new_n946));
  AOI211_X1 g521(.A(new_n925), .B(new_n940), .C1(new_n944), .C2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(new_n940), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n935), .A2(new_n937), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(new_n908), .ZN(new_n950));
  AOI21_X1  g525(.A(KEYINPUT43), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g526(.A(KEYINPUT44), .B1(new_n947), .B2(new_n951), .ZN(new_n952));
  AOI211_X1 g527(.A(KEYINPUT43), .B(new_n940), .C1(new_n944), .C2(new_n946), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n925), .B1(new_n948), .B2(new_n950), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n952), .B1(new_n955), .B2(KEYINPUT44), .ZN(G397));
  NAND2_X1  g531(.A1(G160), .A2(G40), .ZN(new_n957));
  OAI21_X1  g532(.A(KEYINPUT118), .B1(new_n864), .B2(G1384), .ZN(new_n958));
  INV_X1    g533(.A(new_n859), .ZN(new_n959));
  AND3_X1   g534(.A1(new_n490), .A2(new_n862), .A3(new_n495), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n862), .B1(new_n490), .B2(new_n495), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n959), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT118), .ZN(new_n963));
  INV_X1    g538(.A(G1384), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n962), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n957), .B1(new_n958), .B2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(G8), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT49), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n581), .A2(new_n586), .A3(new_n582), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(KEYINPUT121), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT121), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n581), .A2(new_n586), .A3(new_n582), .A4(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n971), .A2(new_n585), .A3(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n974), .A2(KEYINPUT122), .A3(G1981), .ZN(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(G1981), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n583), .A2(new_n585), .A3(new_n977), .A4(new_n586), .ZN(new_n978));
  AOI22_X1  g553(.A1(new_n974), .A2(G1981), .B1(new_n978), .B2(KEYINPUT122), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n969), .B1(new_n976), .B2(new_n979), .ZN(new_n980));
  AND2_X1   g555(.A1(new_n974), .A2(G1981), .ZN(new_n981));
  AND2_X1   g556(.A1(new_n978), .A2(KEYINPUT122), .ZN(new_n982));
  OAI211_X1 g557(.A(KEYINPUT49), .B(new_n975), .C1(new_n981), .C2(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n968), .A2(new_n980), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n697), .A2(G1976), .ZN(new_n985));
  XNOR2_X1  g560(.A(KEYINPUT120), .B(G1976), .ZN(new_n986));
  AOI21_X1  g561(.A(KEYINPUT52), .B1(G288), .B2(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n968), .A2(new_n985), .A3(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(new_n957), .ZN(new_n989));
  AND3_X1   g564(.A1(new_n962), .A2(new_n963), .A3(new_n964), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n963), .B1(new_n962), .B2(new_n964), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n989), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n992), .A2(G8), .A3(new_n985), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(KEYINPUT52), .ZN(new_n994));
  AND3_X1   g569(.A1(new_n984), .A2(new_n988), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(G303), .A2(G8), .ZN(new_n996));
  XNOR2_X1  g571(.A(new_n996), .B(KEYINPUT55), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n958), .A2(KEYINPUT50), .A3(new_n965), .ZN(new_n998));
  XOR2_X1   g573(.A(KEYINPUT119), .B(G2090), .Z(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n499), .A2(new_n964), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT50), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n957), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n998), .A2(new_n1000), .A3(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT45), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1001), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n962), .A2(new_n964), .ZN(new_n1008));
  OAI211_X1 g583(.A(new_n989), .B(new_n1007), .C1(new_n1008), .C2(new_n1006), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(new_n691), .ZN(new_n1010));
  AND2_X1   g585(.A1(new_n1005), .A2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n997), .B1(new_n1011), .B2(new_n967), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n958), .A2(new_n1006), .A3(new_n965), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n957), .B1(new_n1002), .B2(KEYINPUT45), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(new_n771), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1003), .B1(new_n990), .B2(new_n991), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n957), .B1(KEYINPUT50), .B2(new_n1001), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1017), .A2(new_n751), .A3(new_n1018), .ZN(new_n1019));
  AOI211_X1 g594(.A(new_n967), .B(G286), .C1(new_n1016), .C2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(new_n997), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1017), .A2(new_n1000), .A3(new_n1018), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1010), .ZN(new_n1024));
  OAI211_X1 g599(.A(G8), .B(new_n1021), .C1(new_n1023), .C2(new_n1024), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n995), .A2(new_n1012), .A3(new_n1020), .A4(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(KEYINPUT123), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n984), .A2(new_n988), .A3(new_n994), .ZN(new_n1028));
  AOI211_X1 g603(.A(new_n967), .B(new_n997), .C1(new_n1022), .C2(new_n1010), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT123), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1030), .A2(new_n1031), .A3(new_n1012), .A4(new_n1020), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT63), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1027), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(G8), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1033), .B1(new_n1035), .B2(new_n997), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1030), .A2(new_n1036), .A3(new_n1020), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1034), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(G1976), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n984), .A2(new_n1039), .A3(new_n697), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(new_n978), .ZN(new_n1041));
  AOI22_X1  g616(.A1(new_n1041), .A2(new_n968), .B1(new_n995), .B2(new_n1029), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1038), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1016), .A2(new_n1019), .ZN(new_n1044));
  OAI21_X1  g619(.A(G8), .B1(new_n1044), .B2(G286), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(KEYINPUT51), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT51), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1047), .B1(new_n1044), .B2(G286), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1046), .B1(new_n1045), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT53), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1050), .B1(new_n1009), .B2(G2078), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT50), .B1(new_n958), .B2(new_n965), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n989), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n737), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1050), .A2(G2078), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1013), .A2(new_n1014), .A3(new_n1055), .ZN(new_n1056));
  AND3_X1   g631(.A1(new_n1054), .A2(KEYINPUT126), .A3(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(KEYINPUT126), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1051), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  XNOR2_X1  g634(.A(G301), .B(KEYINPUT54), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  AND3_X1   g636(.A1(new_n995), .A2(new_n1012), .A3(new_n1025), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1008), .A2(new_n1006), .ZN(new_n1063));
  AOI21_X1  g638(.A(KEYINPUT45), .B1(new_n962), .B2(new_n964), .ZN(new_n1064));
  NOR3_X1   g639(.A1(new_n1063), .A2(new_n957), .A3(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(new_n1055), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1060), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1066), .A2(new_n1054), .A3(new_n1051), .A4(new_n1067), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1049), .A2(new_n1061), .A3(new_n1062), .A4(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n811), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n966), .A2(new_n807), .ZN(new_n1071));
  AND3_X1   g646(.A1(new_n1070), .A2(KEYINPUT125), .A3(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(KEYINPUT125), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT60), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT125), .ZN(new_n1077));
  AOI21_X1  g652(.A(G1348), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n992), .A2(G2067), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1077), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1070), .A2(KEYINPUT125), .A3(new_n1071), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n600), .B1(new_n1082), .B2(KEYINPUT60), .ZN(new_n1083));
  AOI211_X1 g658(.A(new_n1075), .B(new_n601), .C1(new_n1080), .C2(new_n1081), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1076), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT57), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n569), .A2(new_n570), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1086), .B1(new_n1087), .B2(KEYINPUT124), .ZN(new_n1088));
  XNOR2_X1  g663(.A(G299), .B(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(G1956), .B1(new_n998), .B2(new_n1004), .ZN(new_n1090));
  XNOR2_X1  g665(.A(KEYINPUT56), .B(G2072), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1091), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1009), .A2(new_n1092), .ZN(new_n1093));
  NOR3_X1   g668(.A1(new_n1089), .A2(new_n1090), .A3(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1094), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1089), .B1(new_n1090), .B2(new_n1093), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1095), .A2(KEYINPUT61), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT61), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1096), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1098), .B1(new_n1099), .B2(new_n1094), .ZN(new_n1100));
  AND2_X1   g675(.A1(new_n1097), .A2(new_n1100), .ZN(new_n1101));
  XNOR2_X1  g676(.A(KEYINPUT58), .B(G1341), .ZN(new_n1102));
  OAI22_X1  g677(.A1(new_n966), .A2(new_n1102), .B1(new_n1009), .B2(G1996), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(new_n554), .ZN(new_n1104));
  XNOR2_X1  g679(.A(new_n1104), .B(KEYINPUT59), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1085), .A2(new_n1101), .A3(new_n1105), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1094), .A2(new_n600), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1099), .B1(new_n1107), .B2(new_n1074), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1069), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(KEYINPUT127), .B1(new_n1043), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT127), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1042), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1112), .B1(new_n1034), .B2(new_n1037), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1108), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1097), .A2(new_n1100), .ZN(new_n1115));
  OAI21_X1  g690(.A(KEYINPUT60), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(new_n601), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1082), .A2(KEYINPUT60), .A3(new_n600), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1115), .B1(new_n1119), .B2(new_n1076), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1114), .B1(new_n1120), .B2(new_n1105), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n1111), .B(new_n1113), .C1(new_n1121), .C2(new_n1069), .ZN(new_n1122));
  OR2_X1    g697(.A1(new_n1049), .A2(KEYINPUT62), .ZN(new_n1123));
  AOI21_X1  g698(.A(G301), .B1(new_n1049), .B2(KEYINPUT62), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1123), .A2(new_n1124), .A3(new_n1062), .A4(new_n1059), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1110), .A2(new_n1122), .A3(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1064), .A2(new_n989), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1128), .A2(G1996), .A3(new_n763), .ZN(new_n1129));
  XOR2_X1   g704(.A(new_n1129), .B(KEYINPUT117), .Z(new_n1130));
  NOR2_X1   g705(.A1(new_n1127), .A2(G1996), .ZN(new_n1131));
  XNOR2_X1  g706(.A(new_n1131), .B(KEYINPUT116), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1132), .A2(new_n764), .ZN(new_n1133));
  XNOR2_X1  g708(.A(new_n803), .B(new_n807), .ZN(new_n1134));
  OAI211_X1 g709(.A(new_n1130), .B(new_n1133), .C1(new_n1127), .C2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n720), .A2(new_n722), .ZN(new_n1136));
  OR2_X1    g711(.A1(new_n720), .A2(new_n722), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1127), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  OR3_X1    g713(.A1(new_n1127), .A2(G1986), .A3(G290), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1128), .A2(G1986), .A3(G290), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  XNOR2_X1  g716(.A(new_n1141), .B(KEYINPUT115), .ZN(new_n1142));
  NOR3_X1   g717(.A1(new_n1135), .A2(new_n1138), .A3(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1126), .A2(new_n1143), .ZN(new_n1144));
  XOR2_X1   g719(.A(new_n1139), .B(KEYINPUT48), .Z(new_n1145));
  NOR3_X1   g720(.A1(new_n1135), .A2(new_n1138), .A3(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1134), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1128), .B1(new_n1147), .B2(new_n763), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT46), .ZN(new_n1149));
  AND2_X1   g724(.A1(new_n1132), .A2(new_n1149), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1132), .A2(new_n1149), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1148), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  XOR2_X1   g727(.A(new_n1152), .B(KEYINPUT47), .Z(new_n1153));
  OAI22_X1  g728(.A1(new_n1135), .A2(new_n1137), .B1(G2067), .B2(new_n803), .ZN(new_n1154));
  AOI211_X1 g729(.A(new_n1146), .B(new_n1153), .C1(new_n1128), .C2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1144), .A2(new_n1155), .ZN(G329));
  assign    G231 = 1'b0;
  OAI211_X1 g731(.A(G319), .B(new_n679), .C1(new_n953), .C2(new_n954), .ZN(new_n1158));
  NOR2_X1   g732(.A1(G401), .A2(G227), .ZN(new_n1159));
  NAND2_X1  g733(.A1(new_n883), .A2(new_n1159), .ZN(new_n1160));
  NOR2_X1   g734(.A1(new_n1158), .A2(new_n1160), .ZN(G308));
  NAND2_X1  g735(.A1(new_n948), .A2(new_n950), .ZN(new_n1162));
  AOI21_X1  g736(.A(new_n940), .B1(new_n944), .B2(new_n946), .ZN(new_n1163));
  MUX2_X1   g737(.A(new_n1162), .B(new_n1163), .S(new_n925), .Z(new_n1164));
  AND2_X1   g738(.A1(new_n883), .A2(new_n1159), .ZN(new_n1165));
  NAND4_X1  g739(.A1(new_n1164), .A2(new_n1165), .A3(G319), .A4(new_n679), .ZN(G225));
endmodule


