//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 0 1 0 0 0 0 0 1 0 0 1 1 0 1 1 0 0 1 0 0 0 1 0 1 0 1 1 0 0 0 0 0 1 1 1 0 1 0 0 1 0 1 1 1 0 1 1 1 0 0 1 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:57 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT9), .B(G234), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G902), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n187), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  NAND2_X1  g005(.A1(KEYINPUT83), .A2(KEYINPUT3), .ZN(new_n192));
  INV_X1    g006(.A(G107), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n192), .A2(G104), .A3(new_n193), .ZN(new_n194));
  NOR2_X1   g008(.A1(KEYINPUT83), .A2(KEYINPUT3), .ZN(new_n195));
  OAI21_X1  g009(.A(KEYINPUT84), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G104), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n197), .A2(G107), .ZN(new_n198));
  OR2_X1    g012(.A1(KEYINPUT83), .A2(KEYINPUT3), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT84), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n198), .A2(new_n199), .A3(new_n200), .A4(new_n192), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n196), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT82), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n203), .A2(G104), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n197), .A2(KEYINPUT82), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n193), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(KEYINPUT3), .ZN(new_n207));
  XNOR2_X1  g021(.A(KEYINPUT82), .B(G104), .ZN(new_n208));
  AOI21_X1  g022(.A(G101), .B1(new_n208), .B2(G107), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n202), .A2(new_n207), .A3(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT85), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n208), .A2(G107), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n202), .A2(new_n207), .A3(new_n211), .A4(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G101), .ZN(new_n214));
  AOI22_X1  g028(.A1(new_n201), .A2(new_n196), .B1(new_n206), .B2(KEYINPUT3), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n211), .B1(new_n215), .B2(new_n212), .ZN(new_n216));
  OAI211_X1 g030(.A(KEYINPUT4), .B(new_n210), .C1(new_n214), .C2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n215), .A2(new_n212), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(KEYINPUT85), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT4), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n219), .A2(new_n220), .A3(G101), .A4(new_n213), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT65), .ZN(new_n222));
  INV_X1    g036(.A(G146), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n222), .B1(new_n223), .B2(G143), .ZN(new_n224));
  INV_X1    g038(.A(G143), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n225), .A2(KEYINPUT65), .A3(G146), .ZN(new_n226));
  AND3_X1   g040(.A1(new_n223), .A2(KEYINPUT64), .A3(G143), .ZN(new_n227));
  AOI21_X1  g041(.A(KEYINPUT64), .B1(new_n223), .B2(G143), .ZN(new_n228));
  OAI211_X1 g042(.A(new_n224), .B(new_n226), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  AND2_X1   g043(.A1(KEYINPUT0), .A2(G128), .ZN(new_n230));
  NOR2_X1   g044(.A1(KEYINPUT0), .A2(G128), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n225), .A2(G146), .ZN(new_n233));
  OAI21_X1  g047(.A(KEYINPUT66), .B1(new_n223), .B2(G143), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT66), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n235), .A2(new_n225), .A3(G146), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n233), .B1(new_n234), .B2(new_n236), .ZN(new_n237));
  AOI22_X1  g051(.A1(new_n229), .A2(new_n232), .B1(new_n237), .B2(new_n230), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n217), .A2(new_n221), .A3(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT86), .ZN(new_n240));
  INV_X1    g054(.A(G128), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n223), .A2(G143), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n241), .B1(new_n242), .B2(KEYINPUT1), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n229), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n234), .A2(new_n236), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n241), .A2(KEYINPUT1), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n246), .A2(new_n242), .A3(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n245), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(KEYINPUT10), .ZN(new_n250));
  INV_X1    g064(.A(G101), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n197), .A2(G107), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n251), .B1(new_n206), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n210), .A2(new_n254), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n240), .B1(new_n250), .B2(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n253), .B1(new_n215), .B2(new_n209), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n257), .A2(KEYINPUT86), .A3(KEYINPUT10), .A4(new_n249), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT10), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n248), .B1(new_n237), .B2(new_n243), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n210), .A2(new_n254), .A3(new_n260), .ZN(new_n261));
  AOI22_X1  g075(.A1(new_n256), .A2(new_n258), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT11), .ZN(new_n263));
  INV_X1    g077(.A(G134), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n263), .B1(new_n264), .B2(G137), .ZN(new_n265));
  INV_X1    g079(.A(G137), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n266), .A2(KEYINPUT11), .A3(G134), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n264), .A2(G137), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n265), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(G131), .ZN(new_n270));
  INV_X1    g084(.A(G131), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n265), .A2(new_n267), .A3(new_n271), .A4(new_n268), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  XOR2_X1   g087(.A(new_n273), .B(KEYINPUT87), .Z(new_n274));
  NAND3_X1  g088(.A1(new_n239), .A2(new_n262), .A3(new_n274), .ZN(new_n275));
  XNOR2_X1  g089(.A(G110), .B(G140), .ZN(new_n276));
  INV_X1    g090(.A(G953), .ZN(new_n277));
  AND2_X1   g091(.A1(new_n277), .A2(G227), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n276), .B(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n275), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n273), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n239), .A2(new_n262), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT91), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n282), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n239), .A2(new_n262), .A3(KEYINPUT91), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n281), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n261), .B1(new_n257), .B2(new_n249), .ZN(new_n288));
  XNOR2_X1  g102(.A(KEYINPUT88), .B(KEYINPUT12), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n282), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT90), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n282), .B1(new_n288), .B2(KEYINPUT89), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT89), .ZN(new_n294));
  OAI211_X1 g108(.A(new_n261), .B(new_n294), .C1(new_n257), .C2(new_n249), .ZN(new_n295));
  AOI211_X1 g109(.A(new_n292), .B(KEYINPUT12), .C1(new_n293), .C2(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n249), .B1(new_n210), .B2(new_n254), .ZN(new_n297));
  AND3_X1   g111(.A1(new_n210), .A2(new_n254), .A3(new_n260), .ZN(new_n298));
  OAI21_X1  g112(.A(KEYINPUT89), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n299), .A2(new_n273), .A3(new_n295), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT12), .ZN(new_n301));
  AOI21_X1  g115(.A(KEYINPUT90), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n291), .B1(new_n296), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(new_n275), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n287), .B1(new_n304), .B2(new_n279), .ZN(new_n305));
  OAI21_X1  g119(.A(G469), .B1(new_n305), .B2(G902), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT93), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n303), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(new_n281), .ZN(new_n309));
  OAI211_X1 g123(.A(KEYINPUT93), .B(new_n291), .C1(new_n296), .C2(new_n302), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n283), .A2(new_n284), .ZN(new_n312));
  AND3_X1   g126(.A1(new_n312), .A2(new_n273), .A3(new_n286), .ZN(new_n313));
  INV_X1    g127(.A(new_n275), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n279), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  AOI21_X1  g129(.A(G902), .B1(new_n311), .B2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(G469), .ZN(new_n317));
  AOI22_X1  g131(.A1(KEYINPUT92), .A2(new_n306), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT92), .ZN(new_n319));
  OAI211_X1 g133(.A(new_n319), .B(G469), .C1(new_n305), .C2(G902), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n191), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(G116), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n322), .A2(G119), .ZN(new_n323));
  XNOR2_X1  g137(.A(KEYINPUT67), .B(G116), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n323), .B1(new_n324), .B2(G119), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(KEYINPUT5), .ZN(new_n326));
  INV_X1    g140(.A(new_n323), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n326), .B(G113), .C1(KEYINPUT5), .C2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n322), .A2(KEYINPUT67), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT67), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(G116), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n329), .A2(new_n331), .A3(G119), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(new_n327), .ZN(new_n333));
  XOR2_X1   g147(.A(KEYINPUT2), .B(G113), .Z(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(KEYINPUT68), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT68), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n325), .A2(new_n337), .A3(new_n334), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n328), .A2(new_n339), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n340), .A2(new_n255), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n334), .B1(new_n327), .B2(new_n332), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n337), .B1(new_n325), .B2(new_n334), .ZN(new_n345));
  AND4_X1   g159(.A1(new_n337), .A2(new_n334), .A3(new_n332), .A4(new_n327), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n344), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n221), .A2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n217), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n342), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  XNOR2_X1  g164(.A(G110), .B(G122), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n342), .B(new_n351), .C1(new_n348), .C2(new_n349), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n353), .A2(KEYINPUT6), .A3(new_n354), .ZN(new_n355));
  AOI22_X1  g169(.A1(new_n229), .A2(new_n244), .B1(new_n237), .B2(new_n247), .ZN(new_n356));
  INV_X1    g170(.A(G125), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n358), .B1(new_n357), .B2(new_n238), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n277), .A2(G224), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n360), .B(KEYINPUT94), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n359), .B(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT6), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n350), .A2(new_n363), .A3(new_n352), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n355), .A2(new_n362), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n360), .A2(KEYINPUT7), .ZN(new_n366));
  XNOR2_X1  g180(.A(new_n359), .B(new_n366), .ZN(new_n367));
  OR2_X1    g181(.A1(new_n341), .A2(KEYINPUT95), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n340), .A2(new_n255), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n341), .A2(KEYINPUT95), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  XNOR2_X1  g185(.A(new_n351), .B(KEYINPUT8), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n367), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(G902), .B1(new_n373), .B2(new_n354), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n365), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(G210), .B1(G237), .B2(G902), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n365), .A2(new_n374), .A3(new_n376), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(G214), .B1(G237), .B2(G902), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  XNOR2_X1  g196(.A(G125), .B(G140), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(KEYINPUT16), .ZN(new_n384));
  OR3_X1    g198(.A1(new_n357), .A2(KEYINPUT16), .A3(G140), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(new_n223), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n384), .A2(G146), .A3(new_n385), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n387), .A2(KEYINPUT77), .A3(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT77), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n386), .A2(new_n390), .A3(new_n223), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(KEYINPUT97), .ZN(new_n393));
  NOR2_X1   g207(.A1(G237), .A2(G953), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT96), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n395), .A2(new_n225), .ZN(new_n396));
  NOR2_X1   g210(.A1(KEYINPUT96), .A2(G143), .ZN(new_n397));
  OAI211_X1 g211(.A(G214), .B(new_n394), .C1(new_n396), .C2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n394), .A2(G214), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n399), .B1(new_n395), .B2(new_n225), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(G131), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT17), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n401), .B(new_n271), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n404), .B1(new_n405), .B2(new_n403), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT97), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n389), .A2(new_n407), .A3(new_n391), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n393), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  XNOR2_X1  g223(.A(G113), .B(G122), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n410), .B(new_n197), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n383), .B(new_n223), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT18), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n413), .A2(new_n271), .ZN(new_n414));
  OAI221_X1 g228(.A(new_n412), .B1(new_n401), .B2(new_n414), .C1(new_n402), .C2(new_n413), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n409), .A2(new_n411), .A3(new_n415), .ZN(new_n416));
  XOR2_X1   g230(.A(new_n383), .B(KEYINPUT19), .Z(new_n417));
  OAI21_X1  g231(.A(new_n388), .B1(new_n417), .B2(G146), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n415), .B1(new_n405), .B2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(new_n411), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n416), .A2(new_n421), .ZN(new_n422));
  NOR2_X1   g236(.A1(G475), .A2(G902), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(KEYINPUT20), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT20), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n422), .A2(new_n426), .A3(new_n423), .ZN(new_n427));
  INV_X1    g241(.A(new_n416), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n411), .B1(new_n409), .B2(new_n415), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n190), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  AOI22_X1  g244(.A1(new_n425), .A2(new_n427), .B1(new_n430), .B2(G475), .ZN(new_n431));
  NAND2_X1  g245(.A1(G234), .A2(G237), .ZN(new_n432));
  AND3_X1   g246(.A1(new_n432), .A2(G952), .A3(new_n277), .ZN(new_n433));
  AND3_X1   g247(.A1(new_n432), .A2(G902), .A3(G953), .ZN(new_n434));
  XNOR2_X1  g248(.A(KEYINPUT21), .B(G898), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n433), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n324), .A2(G122), .ZN(new_n438));
  AND2_X1   g252(.A1(KEYINPUT98), .A2(G122), .ZN(new_n439));
  NOR2_X1   g253(.A1(KEYINPUT98), .A2(G122), .ZN(new_n440));
  OAI21_X1  g254(.A(G116), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n438), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(G107), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n438), .A2(new_n193), .A3(new_n441), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT99), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n443), .A2(KEYINPUT99), .A3(new_n444), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT100), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n450), .B1(new_n225), .B2(G128), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n241), .A2(KEYINPUT100), .A3(G143), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n225), .A2(G128), .ZN(new_n454));
  AND3_X1   g268(.A1(new_n453), .A2(new_n264), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(KEYINPUT102), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT102), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT13), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n454), .A2(new_n458), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n459), .B(KEYINPUT101), .ZN(new_n460));
  AOI22_X1  g274(.A1(new_n451), .A2(new_n452), .B1(new_n454), .B2(new_n458), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n457), .B1(new_n462), .B2(G134), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n449), .B(new_n456), .C1(new_n455), .C2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n438), .A2(KEYINPUT14), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n441), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n438), .A2(KEYINPUT14), .ZN(new_n467));
  OAI21_X1  g281(.A(G107), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n264), .B1(new_n453), .B2(new_n454), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n468), .B(new_n444), .C1(new_n455), .C2(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n189), .A2(G217), .A3(new_n277), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  AND3_X1   g286(.A1(new_n464), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n472), .B1(new_n464), .B2(new_n470), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n190), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(G478), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n476), .A2(KEYINPUT15), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n477), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n190), .B(new_n479), .C1(new_n473), .C2(new_n474), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n478), .A2(KEYINPUT103), .A3(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(KEYINPUT103), .B1(new_n478), .B2(new_n480), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n431), .B(new_n437), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n382), .A2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT31), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n394), .A2(G210), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n487), .B(KEYINPUT72), .ZN(new_n488));
  XOR2_X1   g302(.A(KEYINPUT26), .B(G101), .Z(new_n489));
  XNOR2_X1  g303(.A(new_n488), .B(new_n489), .ZN(new_n490));
  XNOR2_X1  g304(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n490), .B(new_n491), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n264), .A2(G137), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n266), .A2(G134), .ZN(new_n494));
  OAI21_X1  g308(.A(G131), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n272), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n496), .B1(new_n245), .B2(new_n248), .ZN(new_n497));
  AOI22_X1  g311(.A1(new_n497), .A2(KEYINPUT69), .B1(new_n238), .B2(new_n273), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT70), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n347), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n339), .A2(KEYINPUT70), .A3(new_n344), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT69), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n502), .B1(new_n356), .B2(new_n496), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n498), .A2(new_n500), .A3(new_n501), .A4(new_n503), .ZN(new_n504));
  AND2_X1   g318(.A1(new_n272), .A2(new_n495), .ZN(new_n505));
  AND2_X1   g319(.A1(new_n224), .A2(new_n226), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT64), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n242), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n223), .A2(KEYINPUT64), .A3(G143), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n243), .B1(new_n506), .B2(new_n510), .ZN(new_n511));
  AND3_X1   g325(.A1(new_n246), .A2(new_n242), .A3(new_n247), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n505), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n229), .A2(new_n232), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n237), .A2(new_n230), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n273), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT30), .ZN(new_n517));
  AND3_X1   g331(.A1(new_n513), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  OAI211_X1 g332(.A(KEYINPUT69), .B(new_n505), .C1(new_n511), .C2(new_n512), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n503), .A2(new_n516), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n518), .B1(KEYINPUT30), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n347), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n492), .B(new_n504), .C1(new_n521), .C2(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n486), .B1(new_n523), .B2(KEYINPUT73), .ZN(new_n524));
  AOI21_X1  g338(.A(KEYINPUT70), .B1(new_n339), .B2(new_n344), .ZN(new_n525));
  AOI211_X1 g339(.A(new_n499), .B(new_n343), .C1(new_n336), .C2(new_n338), .ZN(new_n526));
  NOR3_X1   g340(.A1(new_n520), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n520), .A2(KEYINPUT30), .ZN(new_n528));
  INV_X1    g342(.A(new_n518), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n527), .B1(new_n530), .B2(new_n347), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT73), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n531), .A2(new_n532), .A3(KEYINPUT31), .A4(new_n492), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n524), .A2(new_n533), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n492), .B(KEYINPUT74), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT28), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n500), .A2(new_n501), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n513), .A2(new_n516), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n347), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n536), .B1(new_n504), .B2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT75), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n539), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n525), .A2(new_n526), .ZN(new_n544));
  INV_X1    g358(.A(new_n520), .ZN(new_n545));
  AOI22_X1  g359(.A1(new_n544), .A2(new_n545), .B1(new_n347), .B2(new_n538), .ZN(new_n546));
  NOR3_X1   g360(.A1(new_n546), .A2(KEYINPUT75), .A3(new_n536), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n535), .B1(new_n543), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n534), .A2(new_n548), .ZN(new_n549));
  NOR2_X1   g363(.A1(G472), .A2(G902), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n549), .A2(KEYINPUT32), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(KEYINPUT76), .ZN(new_n552));
  INV_X1    g366(.A(new_n550), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n553), .B1(new_n534), .B2(new_n548), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT76), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n554), .A2(new_n555), .A3(KEYINPUT32), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT32), .ZN(new_n557));
  OAI21_X1  g371(.A(KEYINPUT75), .B1(new_n546), .B2(new_n536), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n541), .A2(new_n542), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n558), .A2(new_n559), .A3(new_n539), .ZN(new_n560));
  AOI22_X1  g374(.A1(new_n560), .A2(new_n535), .B1(new_n524), .B2(new_n533), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n557), .B1(new_n561), .B2(new_n553), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n504), .B1(new_n521), .B2(new_n522), .ZN(new_n563));
  INV_X1    g377(.A(new_n492), .ZN(new_n564));
  AOI21_X1  g378(.A(KEYINPUT29), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n565), .B1(new_n560), .B2(new_n535), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n537), .A2(new_n520), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(new_n504), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(KEYINPUT28), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(new_n539), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  AND2_X1   g385(.A1(new_n492), .A2(KEYINPUT29), .ZN(new_n572));
  AOI21_X1  g386(.A(G902), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n566), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(G472), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n552), .A2(new_n556), .A3(new_n562), .A4(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(G234), .ZN(new_n577));
  OAI21_X1  g391(.A(G217), .B1(new_n577), .B2(G902), .ZN(new_n578));
  INV_X1    g392(.A(G119), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(G128), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n241), .A2(KEYINPUT23), .A3(G119), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n579), .A2(G128), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n580), .B(new_n581), .C1(new_n582), .C2(KEYINPUT23), .ZN(new_n583));
  XOR2_X1   g397(.A(KEYINPUT24), .B(G110), .Z(new_n584));
  XNOR2_X1  g398(.A(G119), .B(G128), .ZN(new_n585));
  AOI22_X1  g399(.A1(new_n583), .A2(G110), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n389), .A2(new_n391), .A3(new_n586), .ZN(new_n587));
  XOR2_X1   g401(.A(KEYINPUT78), .B(G110), .Z(new_n588));
  OAI22_X1  g402(.A1(new_n583), .A2(new_n588), .B1(new_n584), .B2(new_n585), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n383), .A2(new_n223), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n589), .A2(new_n388), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(KEYINPUT22), .B(G137), .ZN(new_n593));
  NOR3_X1   g407(.A1(new_n187), .A2(new_n577), .A3(G953), .ZN(new_n594));
  XOR2_X1   g408(.A(new_n593), .B(new_n594), .Z(new_n595));
  XNOR2_X1  g409(.A(new_n592), .B(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT25), .ZN(new_n597));
  AOI21_X1  g411(.A(G902), .B1(new_n597), .B2(KEYINPUT79), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n597), .A2(KEYINPUT79), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n578), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n601), .B1(new_n600), .B2(new_n599), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n578), .A2(new_n190), .ZN(new_n603));
  XOR2_X1   g417(.A(new_n603), .B(KEYINPUT80), .Z(new_n604));
  NAND2_X1  g418(.A1(new_n596), .A2(new_n604), .ZN(new_n605));
  AND2_X1   g419(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  AND3_X1   g420(.A1(new_n576), .A2(KEYINPUT81), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(KEYINPUT81), .B1(new_n576), .B2(new_n606), .ZN(new_n608));
  OAI211_X1 g422(.A(new_n321), .B(new_n485), .C1(new_n607), .C2(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(G101), .ZN(G3));
  INV_X1    g424(.A(new_n321), .ZN(new_n611));
  AOI21_X1  g425(.A(G902), .B1(new_n534), .B2(new_n548), .ZN(new_n612));
  OAI21_X1  g426(.A(G472), .B1(new_n612), .B2(KEYINPUT104), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT104), .ZN(new_n614));
  NOR3_X1   g428(.A1(new_n561), .A2(new_n614), .A3(G902), .ZN(new_n615));
  OAI21_X1  g429(.A(KEYINPUT105), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n549), .A2(new_n190), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(new_n614), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT105), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n612), .A2(KEYINPUT104), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n618), .A2(new_n619), .A3(new_n620), .A4(G472), .ZN(new_n621));
  INV_X1    g435(.A(new_n554), .ZN(new_n622));
  AND3_X1   g436(.A1(new_n616), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n611), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n378), .A2(KEYINPUT106), .A3(new_n379), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT106), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n365), .A2(new_n374), .A3(new_n627), .A4(new_n376), .ZN(new_n628));
  AND2_X1   g442(.A1(new_n628), .A2(new_n381), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n476), .A2(new_n190), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n464), .A2(new_n470), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(new_n471), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n464), .A2(new_n470), .A3(new_n472), .ZN(new_n634));
  AOI21_X1  g448(.A(G902), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n631), .B1(new_n635), .B2(new_n476), .ZN(new_n636));
  OAI21_X1  g450(.A(KEYINPUT33), .B1(new_n473), .B2(new_n474), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT33), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n633), .A2(new_n638), .A3(new_n634), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n637), .A2(new_n639), .A3(G478), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n636), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n641), .A2(new_n431), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NOR3_X1   g457(.A1(new_n630), .A2(new_n436), .A3(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n625), .A2(new_n606), .A3(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT34), .B(G104), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G6));
  INV_X1    g461(.A(new_n483), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n426), .B1(new_n422), .B2(new_n423), .ZN(new_n649));
  AOI22_X1  g463(.A1(KEYINPUT107), .A2(new_n649), .B1(new_n430), .B2(G475), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT107), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n425), .A2(new_n651), .A3(new_n427), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n648), .A2(new_n481), .A3(new_n650), .A4(new_n652), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n630), .A2(new_n436), .A3(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n625), .A2(new_n606), .A3(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT35), .B(G107), .Z(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G9));
  INV_X1    g471(.A(new_n595), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n658), .A2(KEYINPUT36), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n592), .B(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n604), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n602), .A2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  NOR3_X1   g477(.A1(new_n382), .A2(new_n663), .A3(new_n484), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n321), .A2(new_n623), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(KEYINPUT37), .B(G110), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(KEYINPUT108), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n665), .B(new_n667), .ZN(G12));
  NAND2_X1  g482(.A1(new_n576), .A2(new_n662), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n630), .ZN(new_n671));
  INV_X1    g485(.A(G900), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n433), .B1(new_n434), .B2(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n653), .A2(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n321), .A2(new_n670), .A3(new_n671), .A4(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G128), .ZN(G30));
  XNOR2_X1  g490(.A(new_n673), .B(KEYINPUT39), .ZN(new_n677));
  OR2_X1    g491(.A1(new_n611), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(KEYINPUT40), .ZN(new_n679));
  OR3_X1    g493(.A1(new_n611), .A2(KEYINPUT40), .A3(new_n677), .ZN(new_n680));
  XNOR2_X1  g494(.A(KEYINPUT109), .B(KEYINPUT38), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n380), .A2(new_n682), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n681), .B1(new_n378), .B2(new_n379), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n523), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n687), .B1(new_n535), .B2(new_n568), .ZN(new_n688));
  OAI21_X1  g502(.A(G472), .B1(new_n688), .B2(G902), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n552), .A2(new_n556), .A3(new_n562), .A4(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NOR3_X1   g505(.A1(new_n482), .A2(new_n431), .A3(new_n483), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n692), .A2(new_n381), .A3(new_n663), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n686), .A2(new_n691), .A3(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n679), .A2(new_n680), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G143), .ZN(G45));
  NOR3_X1   g510(.A1(new_n641), .A2(new_n431), .A3(new_n673), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n698), .A2(new_n663), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n321), .A2(new_n576), .A3(new_n671), .A4(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G146), .ZN(G48));
  NAND2_X1  g515(.A1(new_n300), .A2(new_n301), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n292), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n300), .A2(KEYINPUT90), .A3(new_n301), .ZN(new_n704));
  AOI22_X1  g518(.A1(new_n703), .A2(new_n704), .B1(new_n288), .B2(new_n290), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n705), .A2(KEYINPUT93), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n310), .A2(new_n309), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n315), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n190), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(G469), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT110), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n708), .A2(new_n317), .A3(new_n190), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n710), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n709), .A2(KEYINPUT110), .A3(G469), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n191), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  AND2_X1   g529(.A1(new_n576), .A2(new_n606), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n715), .A2(new_n716), .A3(new_n644), .ZN(new_n717));
  XNOR2_X1  g531(.A(KEYINPUT41), .B(G113), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n717), .B(new_n718), .ZN(G15));
  NAND2_X1  g533(.A1(new_n713), .A2(new_n714), .ZN(new_n720));
  INV_X1    g534(.A(new_n191), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n720), .A2(new_n716), .A3(new_n654), .A4(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G116), .ZN(G18));
  NOR2_X1   g537(.A1(new_n669), .A2(new_n484), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n715), .A2(new_n671), .A3(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G119), .ZN(G21));
  NAND3_X1  g540(.A1(new_n626), .A2(new_n692), .A3(new_n629), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT111), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n626), .A2(new_n692), .A3(new_n629), .A4(KEYINPUT111), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n617), .A2(G472), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n570), .A2(new_n535), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n534), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(new_n550), .ZN(new_n735));
  AND2_X1   g549(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  AND3_X1   g550(.A1(new_n736), .A2(new_n606), .A3(new_n437), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n715), .A2(new_n731), .A3(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(KEYINPUT112), .B(G122), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n738), .B(new_n739), .ZN(G24));
  AND4_X1   g554(.A1(new_n662), .A2(new_n697), .A3(new_n735), .A4(new_n732), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n715), .A2(new_n671), .A3(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(KEYINPUT113), .B(G125), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n742), .B(new_n743), .ZN(G27));
  INV_X1    g558(.A(KEYINPUT115), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n562), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n746), .A2(new_n551), .A3(new_n575), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n562), .A2(new_n745), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n606), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(new_n697), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n712), .A2(new_n306), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(KEYINPUT114), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT114), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n712), .A2(new_n754), .A3(new_n306), .ZN(new_n755));
  INV_X1    g569(.A(new_n381), .ZN(new_n756));
  NOR3_X1   g570(.A1(new_n380), .A2(new_n756), .A3(new_n191), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n753), .A2(new_n755), .A3(new_n757), .ZN(new_n758));
  OAI21_X1  g572(.A(KEYINPUT42), .B1(new_n751), .B2(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(new_n758), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n698), .A2(KEYINPUT42), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n760), .A2(new_n716), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n759), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(new_n271), .ZN(G33));
  NAND3_X1  g578(.A1(new_n760), .A2(new_n716), .A3(new_n674), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G134), .ZN(G36));
  NOR2_X1   g580(.A1(new_n317), .A2(new_n190), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n279), .B1(new_n705), .B2(new_n314), .ZN(new_n768));
  INV_X1    g582(.A(new_n287), .ZN(new_n769));
  AOI21_X1  g583(.A(KEYINPUT45), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  OAI21_X1  g584(.A(KEYINPUT116), .B1(new_n770), .B2(new_n317), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT116), .ZN(new_n772));
  OAI211_X1 g586(.A(new_n772), .B(G469), .C1(new_n305), .C2(KEYINPUT45), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n305), .A2(KEYINPUT45), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n771), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(KEYINPUT117), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT117), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n771), .A2(new_n774), .A3(new_n777), .A4(new_n773), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n767), .B1(new_n776), .B2(new_n778), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n712), .B1(new_n779), .B2(KEYINPUT46), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT46), .ZN(new_n781));
  AOI211_X1 g595(.A(new_n781), .B(new_n767), .C1(new_n776), .C2(new_n778), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n721), .B1(new_n780), .B2(new_n782), .ZN(new_n783));
  OR2_X1    g597(.A1(new_n783), .A2(new_n677), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n380), .A2(new_n756), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n430), .A2(G475), .ZN(new_n787));
  INV_X1    g601(.A(new_n427), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n787), .B1(new_n788), .B2(new_n649), .ZN(new_n789));
  OAI21_X1  g603(.A(KEYINPUT43), .B1(new_n641), .B2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT43), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n431), .A2(new_n791), .A3(new_n640), .A4(new_n636), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n624), .A2(new_n662), .A3(new_n790), .A4(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT44), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n786), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n795), .B1(new_n794), .B2(new_n793), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n784), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(new_n266), .ZN(G39));
  OR4_X1    g612(.A1(new_n576), .A2(new_n786), .A3(new_n606), .A4(new_n698), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT47), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n783), .A2(new_n800), .ZN(new_n801));
  OAI211_X1 g615(.A(KEYINPUT47), .B(new_n721), .C1(new_n780), .C2(new_n782), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n799), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  XOR2_X1   g617(.A(new_n803), .B(G140), .Z(G42));
  NOR2_X1   g618(.A1(G952), .A2(G953), .ZN(new_n805));
  XOR2_X1   g619(.A(new_n805), .B(KEYINPUT123), .Z(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n725), .A2(new_n738), .A3(new_n717), .A4(new_n722), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n635), .A2(new_n479), .ZN(new_n809));
  INV_X1    g623(.A(new_n480), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n811), .A2(new_n789), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n437), .B1(new_n642), .B2(new_n812), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n813), .A2(new_n382), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n321), .A2(new_n623), .A3(new_n606), .A4(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n609), .A2(new_n815), .A3(new_n665), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(KEYINPUT118), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT118), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n609), .A2(new_n815), .A3(new_n818), .A4(new_n665), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n808), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n318), .A2(new_n320), .ZN(new_n821));
  INV_X1    g635(.A(new_n673), .ZN(new_n822));
  AND4_X1   g636(.A1(new_n811), .A2(new_n650), .A3(new_n652), .A4(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n670), .A2(new_n821), .A3(new_n757), .A4(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n753), .A2(new_n741), .A3(new_n755), .A4(new_n757), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  AND4_X1   g640(.A1(new_n759), .A2(new_n826), .A3(new_n762), .A4(new_n765), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n662), .A2(new_n191), .A3(new_n673), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n753), .A2(new_n755), .A3(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT119), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n753), .A2(KEYINPUT119), .A3(new_n755), .A4(new_n828), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n831), .A2(new_n690), .A3(new_n731), .A4(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n742), .A2(new_n700), .A3(new_n675), .ZN(new_n835));
  OAI21_X1  g649(.A(KEYINPUT52), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n742), .A2(new_n675), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT52), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n837), .A2(new_n838), .A3(new_n833), .A4(new_n700), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n820), .A2(new_n827), .A3(new_n836), .A4(new_n839), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n834), .A2(new_n837), .A3(new_n835), .ZN(new_n841));
  OAI21_X1  g655(.A(KEYINPUT53), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n836), .A2(new_n839), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT53), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n843), .A2(new_n844), .A3(new_n820), .A4(new_n827), .ZN(new_n845));
  AOI21_X1  g659(.A(KEYINPUT54), .B1(new_n842), .B2(new_n845), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n820), .A2(new_n827), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n847), .A2(KEYINPUT120), .A3(new_n843), .A4(KEYINPUT53), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT120), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n849), .B1(new_n840), .B2(new_n844), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n844), .B1(new_n840), .B2(new_n841), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n848), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n846), .B1(KEYINPUT54), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n720), .A2(new_n191), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n801), .A2(new_n802), .A3(new_n854), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n790), .A2(new_n792), .A3(new_n433), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n856), .A2(new_n606), .A3(new_n736), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n857), .A2(new_n786), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n691), .A2(new_n606), .A3(new_n433), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n789), .B1(new_n640), .B2(new_n636), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n860), .A2(new_n715), .A3(new_n785), .A4(new_n861), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n736), .A2(new_n662), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n715), .A2(new_n863), .A3(new_n785), .A4(new_n856), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n857), .A2(new_n685), .A3(new_n381), .ZN(new_n865));
  AND3_X1   g679(.A1(new_n865), .A2(new_n715), .A3(KEYINPUT50), .ZN(new_n866));
  AOI21_X1  g680(.A(KEYINPUT50), .B1(new_n865), .B2(new_n715), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n862), .B(new_n864), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n868), .B(KEYINPUT121), .ZN(new_n869));
  AOI21_X1  g683(.A(KEYINPUT51), .B1(new_n859), .B2(new_n869), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n715), .A2(new_n750), .A3(new_n785), .A4(new_n856), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n871), .B(KEYINPUT48), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n715), .A2(new_n671), .ZN(new_n873));
  OR2_X1    g687(.A1(new_n873), .A2(new_n857), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n860), .A2(new_n715), .A3(new_n642), .A4(new_n785), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n874), .A2(G952), .A3(new_n277), .A4(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT122), .ZN(new_n877));
  AND2_X1   g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n876), .A2(new_n877), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n872), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(new_n868), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(KEYINPUT51), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n882), .B1(new_n855), .B2(new_n858), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n870), .A2(new_n880), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n807), .B1(new_n853), .B2(new_n884), .ZN(new_n885));
  XOR2_X1   g699(.A(new_n720), .B(KEYINPUT49), .Z(new_n886));
  NAND2_X1  g700(.A1(new_n691), .A2(new_n606), .ZN(new_n887));
  NOR4_X1   g701(.A1(new_n641), .A2(new_n789), .A3(new_n756), .A4(new_n191), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n686), .A2(new_n888), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n886), .A2(new_n887), .A3(new_n889), .ZN(new_n890));
  OAI21_X1  g704(.A(KEYINPUT124), .B1(new_n885), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n852), .A2(KEYINPUT54), .ZN(new_n892));
  INV_X1    g706(.A(new_n846), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n892), .A2(new_n884), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(new_n806), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT124), .ZN(new_n896));
  INV_X1    g710(.A(new_n890), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n891), .A2(new_n898), .ZN(G75));
  NOR2_X1   g713(.A1(new_n277), .A2(G952), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n842), .A2(new_n845), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n902), .A2(new_n190), .ZN(new_n903));
  AOI21_X1  g717(.A(KEYINPUT56), .B1(new_n903), .B2(G210), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n355), .A2(new_n364), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n905), .B(new_n362), .Z(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(KEYINPUT55), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n901), .B1(new_n904), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n909), .B1(new_n904), .B2(new_n908), .ZN(G51));
  XNOR2_X1  g724(.A(new_n902), .B(KEYINPUT54), .ZN(new_n911));
  XOR2_X1   g725(.A(new_n767), .B(KEYINPUT57), .Z(new_n912));
  OAI21_X1  g726(.A(new_n708), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n903), .A2(new_n778), .A3(new_n776), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n900), .B1(new_n913), .B2(new_n914), .ZN(G54));
  NAND3_X1  g729(.A1(new_n903), .A2(KEYINPUT58), .A3(G475), .ZN(new_n916));
  INV_X1    g730(.A(new_n422), .ZN(new_n917));
  AND2_X1   g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n916), .A2(new_n917), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n918), .A2(new_n919), .A3(new_n900), .ZN(G60));
  NAND2_X1  g734(.A1(new_n637), .A2(new_n639), .ZN(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n631), .B(KEYINPUT59), .ZN(new_n923));
  OR2_X1    g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n901), .B1(new_n911), .B2(new_n924), .ZN(new_n925));
  OR2_X1    g739(.A1(new_n853), .A2(new_n923), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n925), .B1(new_n922), .B2(new_n926), .ZN(G63));
  INV_X1    g741(.A(new_n902), .ZN(new_n928));
  NAND2_X1  g742(.A1(G217), .A2(G902), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n929), .B(KEYINPUT60), .Z(new_n930));
  NAND2_X1  g744(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(new_n596), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n928), .A2(new_n660), .A3(new_n930), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n933), .A2(new_n901), .A3(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT61), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n933), .A2(KEYINPUT61), .A3(new_n901), .A4(new_n934), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(G66));
  INV_X1    g753(.A(G224), .ZN(new_n940));
  OAI21_X1  g754(.A(G953), .B1(new_n435), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n941), .B1(new_n820), .B2(G953), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n905), .B1(G898), .B2(new_n277), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n942), .B(new_n943), .ZN(G69));
  OR2_X1    g758(.A1(new_n797), .A2(new_n803), .ZN(new_n945));
  AND3_X1   g759(.A1(new_n759), .A2(new_n762), .A3(new_n765), .ZN(new_n946));
  INV_X1    g760(.A(new_n835), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n750), .A2(new_n731), .ZN(new_n948));
  OAI211_X1 g762(.A(new_n946), .B(new_n947), .C1(new_n784), .C2(new_n948), .ZN(new_n949));
  OR3_X1    g763(.A1(new_n945), .A2(G953), .A3(new_n949), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n530), .B(new_n417), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n951), .B1(G900), .B2(G953), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n797), .A2(new_n803), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n607), .A2(new_n608), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n642), .A2(new_n812), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(KEYINPUT126), .ZN(new_n957));
  NOR4_X1   g771(.A1(new_n678), .A2(new_n955), .A3(new_n786), .A4(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n695), .A2(new_n947), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT62), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n695), .A2(KEYINPUT62), .A3(new_n947), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n958), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n954), .A2(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT127), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n954), .A2(KEYINPUT127), .A3(new_n963), .ZN(new_n967));
  AOI21_X1  g781(.A(G953), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n951), .B(KEYINPUT125), .Z(new_n969));
  OAI21_X1  g783(.A(new_n953), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n277), .B1(G227), .B2(G900), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(new_n971), .ZN(new_n973));
  OAI211_X1 g787(.A(new_n953), .B(new_n973), .C1(new_n968), .C2(new_n969), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n972), .A2(new_n974), .ZN(G72));
  INV_X1    g789(.A(new_n820), .ZN(new_n976));
  NOR3_X1   g790(.A1(new_n945), .A2(new_n976), .A3(new_n949), .ZN(new_n977));
  NAND2_X1  g791(.A1(G472), .A2(G902), .ZN(new_n978));
  XOR2_X1   g792(.A(new_n978), .B(KEYINPUT63), .Z(new_n979));
  INV_X1    g793(.A(new_n979), .ZN(new_n980));
  OAI211_X1 g794(.A(new_n564), .B(new_n531), .C1(new_n977), .C2(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(new_n852), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n531), .A2(new_n492), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n979), .B1(new_n983), .B2(new_n687), .ZN(new_n984));
  OAI211_X1 g798(.A(new_n981), .B(new_n901), .C1(new_n982), .C2(new_n984), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n966), .A2(new_n820), .A3(new_n967), .ZN(new_n986));
  AOI211_X1 g800(.A(new_n564), .B(new_n531), .C1(new_n986), .C2(new_n979), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n985), .A2(new_n987), .ZN(G57));
endmodule


