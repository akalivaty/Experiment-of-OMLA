

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X2 U550 ( .A(n641), .ZN(n642) );
  NAND2_X2 U551 ( .A1(G8), .A2(n641), .ZN(n697) );
  XNOR2_X1 U552 ( .A(n595), .B(KEYINPUT91), .ZN(n713) );
  NOR2_X1 U553 ( .A1(n522), .A2(G2105), .ZN(n518) );
  XNOR2_X1 U554 ( .A(n601), .B(n600), .ZN(n602) );
  NOR2_X1 U555 ( .A1(G2105), .A2(G2104), .ZN(n523) );
  NOR2_X1 U556 ( .A1(n593), .A2(n757), .ZN(n515) );
  INV_X1 U557 ( .A(KEYINPUT30), .ZN(n600) );
  INV_X1 U558 ( .A(KEYINPUT98), .ZN(n658) );
  NAND2_X1 U559 ( .A1(G8), .A2(n664), .ZN(n665) );
  INV_X1 U560 ( .A(KEYINPUT65), .ZN(n517) );
  AND2_X1 U561 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U562 ( .A1(G651), .A2(n564), .ZN(n788) );
  XNOR2_X1 U563 ( .A(KEYINPUT40), .B(KEYINPUT103), .ZN(n754) );
  AND2_X1 U564 ( .A1(G2105), .A2(G2104), .ZN(n889) );
  NAND2_X1 U565 ( .A1(n889), .A2(G114), .ZN(n516) );
  XNOR2_X1 U566 ( .A(n516), .B(KEYINPUT90), .ZN(n521) );
  XOR2_X1 U567 ( .A(G2104), .B(KEYINPUT64), .Z(n522) );
  XNOR2_X1 U568 ( .A(n518), .B(n517), .ZN(n587) );
  INV_X1 U569 ( .A(n587), .ZN(n519) );
  INV_X1 U570 ( .A(n519), .ZN(n886) );
  NAND2_X1 U571 ( .A1(G102), .A2(n886), .ZN(n520) );
  NAND2_X1 U572 ( .A1(n521), .A2(n520), .ZN(n527) );
  AND2_X1 U573 ( .A1(G2105), .A2(n522), .ZN(n890) );
  NAND2_X1 U574 ( .A1(G126), .A2(n890), .ZN(n525) );
  XOR2_X1 U575 ( .A(KEYINPUT17), .B(n523), .Z(n885) );
  NAND2_X1 U576 ( .A1(G138), .A2(n885), .ZN(n524) );
  NAND2_X1 U577 ( .A1(n525), .A2(n524), .ZN(n526) );
  NOR2_X1 U578 ( .A1(n527), .A2(n526), .ZN(G164) );
  XOR2_X1 U579 ( .A(G543), .B(KEYINPUT0), .Z(n564) );
  NAND2_X1 U580 ( .A1(G50), .A2(n788), .ZN(n531) );
  INV_X1 U581 ( .A(G651), .ZN(n533) );
  NOR2_X1 U582 ( .A1(G543), .A2(n533), .ZN(n529) );
  XNOR2_X1 U583 ( .A(KEYINPUT1), .B(KEYINPUT67), .ZN(n528) );
  XNOR2_X1 U584 ( .A(n529), .B(n528), .ZN(n789) );
  NAND2_X1 U585 ( .A1(G62), .A2(n789), .ZN(n530) );
  NAND2_X1 U586 ( .A1(n531), .A2(n530), .ZN(n532) );
  XOR2_X1 U587 ( .A(KEYINPUT84), .B(n532), .Z(n537) );
  NOR2_X1 U588 ( .A1(n564), .A2(n533), .ZN(n796) );
  NAND2_X1 U589 ( .A1(n796), .A2(G75), .ZN(n535) );
  NOR2_X1 U590 ( .A1(G651), .A2(G543), .ZN(n793) );
  NAND2_X1 U591 ( .A1(G88), .A2(n793), .ZN(n534) );
  AND2_X1 U592 ( .A1(n535), .A2(n534), .ZN(n536) );
  NAND2_X1 U593 ( .A1(n537), .A2(n536), .ZN(G303) );
  NAND2_X1 U594 ( .A1(n789), .A2(G63), .ZN(n538) );
  XOR2_X1 U595 ( .A(KEYINPUT75), .B(n538), .Z(n540) );
  NAND2_X1 U596 ( .A1(n788), .A2(G51), .ZN(n539) );
  NAND2_X1 U597 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U598 ( .A(KEYINPUT6), .B(n541), .ZN(n548) );
  NAND2_X1 U599 ( .A1(n793), .A2(G89), .ZN(n542) );
  XNOR2_X1 U600 ( .A(n542), .B(KEYINPUT4), .ZN(n544) );
  NAND2_X1 U601 ( .A1(G76), .A2(n796), .ZN(n543) );
  NAND2_X1 U602 ( .A1(n544), .A2(n543), .ZN(n545) );
  XOR2_X1 U603 ( .A(KEYINPUT5), .B(n545), .Z(n546) );
  XNOR2_X1 U604 ( .A(KEYINPUT74), .B(n546), .ZN(n547) );
  NOR2_X1 U605 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U606 ( .A(KEYINPUT7), .B(n549), .Z(G168) );
  NAND2_X1 U607 ( .A1(G77), .A2(n796), .ZN(n551) );
  NAND2_X1 U608 ( .A1(G90), .A2(n793), .ZN(n550) );
  NAND2_X1 U609 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U610 ( .A(KEYINPUT9), .B(n552), .ZN(n556) );
  NAND2_X1 U611 ( .A1(n788), .A2(G52), .ZN(n554) );
  NAND2_X1 U612 ( .A1(G64), .A2(n789), .ZN(n553) );
  AND2_X1 U613 ( .A1(n554), .A2(n553), .ZN(n555) );
  NAND2_X1 U614 ( .A1(n556), .A2(n555), .ZN(G301) );
  NAND2_X1 U615 ( .A1(G78), .A2(n796), .ZN(n558) );
  NAND2_X1 U616 ( .A1(G91), .A2(n793), .ZN(n557) );
  NAND2_X1 U617 ( .A1(n558), .A2(n557), .ZN(n561) );
  NAND2_X1 U618 ( .A1(G53), .A2(n788), .ZN(n559) );
  XNOR2_X1 U619 ( .A(KEYINPUT69), .B(n559), .ZN(n560) );
  NOR2_X1 U620 ( .A1(n561), .A2(n560), .ZN(n563) );
  NAND2_X1 U621 ( .A1(n789), .A2(G65), .ZN(n562) );
  NAND2_X1 U622 ( .A1(n563), .A2(n562), .ZN(G299) );
  XOR2_X1 U623 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U624 ( .A1(G87), .A2(n564), .ZN(n565) );
  XNOR2_X1 U625 ( .A(n565), .B(KEYINPUT82), .ZN(n570) );
  NAND2_X1 U626 ( .A1(G49), .A2(n788), .ZN(n567) );
  NAND2_X1 U627 ( .A1(G74), .A2(G651), .ZN(n566) );
  NAND2_X1 U628 ( .A1(n567), .A2(n566), .ZN(n568) );
  NOR2_X1 U629 ( .A1(n789), .A2(n568), .ZN(n569) );
  NAND2_X1 U630 ( .A1(n570), .A2(n569), .ZN(G288) );
  NAND2_X1 U631 ( .A1(n788), .A2(G48), .ZN(n577) );
  NAND2_X1 U632 ( .A1(G86), .A2(n793), .ZN(n572) );
  NAND2_X1 U633 ( .A1(G61), .A2(n789), .ZN(n571) );
  NAND2_X1 U634 ( .A1(n572), .A2(n571), .ZN(n575) );
  NAND2_X1 U635 ( .A1(n796), .A2(G73), .ZN(n573) );
  XOR2_X1 U636 ( .A(KEYINPUT2), .B(n573), .Z(n574) );
  NOR2_X1 U637 ( .A1(n575), .A2(n574), .ZN(n576) );
  NAND2_X1 U638 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U639 ( .A(KEYINPUT83), .B(n578), .Z(G305) );
  NAND2_X1 U640 ( .A1(G85), .A2(n793), .ZN(n579) );
  XNOR2_X1 U641 ( .A(n579), .B(KEYINPUT66), .ZN(n581) );
  NAND2_X1 U642 ( .A1(n796), .A2(G72), .ZN(n580) );
  NAND2_X1 U643 ( .A1(n581), .A2(n580), .ZN(n584) );
  NAND2_X1 U644 ( .A1(G60), .A2(n789), .ZN(n582) );
  XOR2_X1 U645 ( .A(KEYINPUT68), .B(n582), .Z(n583) );
  NOR2_X1 U646 ( .A1(n584), .A2(n583), .ZN(n586) );
  NAND2_X1 U647 ( .A1(n788), .A2(G47), .ZN(n585) );
  NAND2_X1 U648 ( .A1(n586), .A2(n585), .ZN(G290) );
  NAND2_X1 U649 ( .A1(n587), .A2(G101), .ZN(n588) );
  XOR2_X1 U650 ( .A(KEYINPUT23), .B(n588), .Z(n590) );
  NAND2_X1 U651 ( .A1(n885), .A2(G137), .ZN(n589) );
  NAND2_X1 U652 ( .A1(n590), .A2(n589), .ZN(n756) );
  INV_X1 U653 ( .A(n756), .ZN(n594) );
  INV_X1 U654 ( .A(G40), .ZN(n593) );
  NAND2_X1 U655 ( .A1(G113), .A2(n889), .ZN(n592) );
  NAND2_X1 U656 ( .A1(G125), .A2(n890), .ZN(n591) );
  NAND2_X1 U657 ( .A1(n592), .A2(n591), .ZN(n757) );
  NAND2_X1 U658 ( .A1(n594), .A2(n515), .ZN(n595) );
  NOR2_X1 U659 ( .A1(G164), .A2(G1384), .ZN(n715) );
  NAND2_X2 U660 ( .A1(n713), .A2(n715), .ZN(n641) );
  NOR2_X1 U661 ( .A1(G1971), .A2(n697), .ZN(n597) );
  NOR2_X1 U662 ( .A1(G2090), .A2(n641), .ZN(n596) );
  NOR2_X1 U663 ( .A1(n597), .A2(n596), .ZN(n598) );
  NAND2_X1 U664 ( .A1(n598), .A2(G303), .ZN(n663) );
  NOR2_X1 U665 ( .A1(G1966), .A2(n697), .ZN(n668) );
  NOR2_X1 U666 ( .A1(G2084), .A2(n641), .ZN(n666) );
  NOR2_X1 U667 ( .A1(n668), .A2(n666), .ZN(n599) );
  AND2_X1 U668 ( .A1(n599), .A2(G8), .ZN(n601) );
  XOR2_X1 U669 ( .A(KEYINPUT99), .B(n602), .Z(n603) );
  NOR2_X1 U670 ( .A1(G168), .A2(n603), .ZN(n607) );
  XOR2_X1 U671 ( .A(G2078), .B(KEYINPUT25), .Z(n976) );
  NOR2_X1 U672 ( .A1(n976), .A2(n641), .ZN(n605) );
  NOR2_X1 U673 ( .A1(n642), .A2(G1961), .ZN(n604) );
  NOR2_X1 U674 ( .A1(n605), .A2(n604), .ZN(n655) );
  AND2_X1 U675 ( .A1(G301), .A2(n655), .ZN(n606) );
  NOR2_X1 U676 ( .A1(n607), .A2(n606), .ZN(n609) );
  INV_X1 U677 ( .A(n609), .ZN(n608) );
  NAND2_X1 U678 ( .A1(n608), .A2(KEYINPUT31), .ZN(n612) );
  INV_X1 U679 ( .A(KEYINPUT31), .ZN(n610) );
  NAND2_X1 U680 ( .A1(n610), .A2(n609), .ZN(n611) );
  NAND2_X1 U681 ( .A1(n612), .A2(n611), .ZN(n661) );
  NAND2_X1 U682 ( .A1(n642), .A2(G2072), .ZN(n613) );
  XNOR2_X1 U683 ( .A(n613), .B(KEYINPUT27), .ZN(n615) );
  INV_X1 U684 ( .A(G1956), .ZN(n948) );
  NOR2_X1 U685 ( .A1(n948), .A2(n642), .ZN(n614) );
  NOR2_X1 U686 ( .A1(n615), .A2(n614), .ZN(n618) );
  INV_X1 U687 ( .A(G299), .ZN(n921) );
  NOR2_X1 U688 ( .A1(n618), .A2(n921), .ZN(n617) );
  INV_X1 U689 ( .A(KEYINPUT28), .ZN(n616) );
  XNOR2_X1 U690 ( .A(n617), .B(n616), .ZN(n653) );
  NAND2_X1 U691 ( .A1(n921), .A2(n618), .ZN(n651) );
  NAND2_X1 U692 ( .A1(n642), .A2(G1996), .ZN(n619) );
  XNOR2_X1 U693 ( .A(n619), .B(KEYINPUT26), .ZN(n632) );
  AND2_X1 U694 ( .A1(n641), .A2(G1341), .ZN(n630) );
  NAND2_X1 U695 ( .A1(n793), .A2(G81), .ZN(n620) );
  XNOR2_X1 U696 ( .A(n620), .B(KEYINPUT12), .ZN(n622) );
  NAND2_X1 U697 ( .A1(G68), .A2(n796), .ZN(n621) );
  NAND2_X1 U698 ( .A1(n622), .A2(n621), .ZN(n623) );
  XNOR2_X1 U699 ( .A(KEYINPUT13), .B(n623), .ZN(n629) );
  NAND2_X1 U700 ( .A1(G43), .A2(n788), .ZN(n624) );
  XNOR2_X1 U701 ( .A(n624), .B(KEYINPUT71), .ZN(n627) );
  NAND2_X1 U702 ( .A1(G56), .A2(n789), .ZN(n625) );
  XOR2_X1 U703 ( .A(KEYINPUT14), .B(n625), .Z(n626) );
  NOR2_X1 U704 ( .A1(n627), .A2(n626), .ZN(n628) );
  NAND2_X1 U705 ( .A1(n629), .A2(n628), .ZN(n930) );
  NOR2_X1 U706 ( .A1(n630), .A2(n930), .ZN(n631) );
  AND2_X1 U707 ( .A1(n632), .A2(n631), .ZN(n646) );
  NAND2_X1 U708 ( .A1(G79), .A2(n796), .ZN(n634) );
  NAND2_X1 U709 ( .A1(G54), .A2(n788), .ZN(n633) );
  NAND2_X1 U710 ( .A1(n634), .A2(n633), .ZN(n639) );
  NAND2_X1 U711 ( .A1(G92), .A2(n793), .ZN(n636) );
  NAND2_X1 U712 ( .A1(G66), .A2(n789), .ZN(n635) );
  NAND2_X1 U713 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U714 ( .A(KEYINPUT72), .B(n637), .ZN(n638) );
  NOR2_X1 U715 ( .A1(n639), .A2(n638), .ZN(n640) );
  XNOR2_X1 U716 ( .A(n640), .B(KEYINPUT15), .ZN(n934) );
  NAND2_X1 U717 ( .A1(G1348), .A2(n641), .ZN(n644) );
  NAND2_X1 U718 ( .A1(G2067), .A2(n642), .ZN(n643) );
  NAND2_X1 U719 ( .A1(n644), .A2(n643), .ZN(n647) );
  NOR2_X1 U720 ( .A1(n934), .A2(n647), .ZN(n645) );
  OR2_X1 U721 ( .A1(n646), .A2(n645), .ZN(n649) );
  NAND2_X1 U722 ( .A1(n934), .A2(n647), .ZN(n648) );
  NAND2_X1 U723 ( .A1(n649), .A2(n648), .ZN(n650) );
  NAND2_X1 U724 ( .A1(n651), .A2(n650), .ZN(n652) );
  NAND2_X1 U725 ( .A1(n653), .A2(n652), .ZN(n654) );
  XNOR2_X1 U726 ( .A(n654), .B(KEYINPUT29), .ZN(n657) );
  NOR2_X1 U727 ( .A1(G301), .A2(n655), .ZN(n656) );
  NOR2_X1 U728 ( .A1(n657), .A2(n656), .ZN(n659) );
  XNOR2_X1 U729 ( .A(n659), .B(n658), .ZN(n660) );
  NAND2_X1 U730 ( .A1(n661), .A2(n660), .ZN(n667) );
  NAND2_X1 U731 ( .A1(n667), .A2(G286), .ZN(n662) );
  NAND2_X1 U732 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U733 ( .A(n665), .B(KEYINPUT32), .ZN(n689) );
  NAND2_X1 U734 ( .A1(G8), .A2(n666), .ZN(n671) );
  INV_X1 U735 ( .A(n667), .ZN(n669) );
  NOR2_X1 U736 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U737 ( .A1(n671), .A2(n670), .ZN(n690) );
  NOR2_X1 U738 ( .A1(G1976), .A2(G288), .ZN(n681) );
  INV_X1 U739 ( .A(n697), .ZN(n674) );
  NAND2_X1 U740 ( .A1(n681), .A2(n674), .ZN(n672) );
  NAND2_X1 U741 ( .A1(n672), .A2(KEYINPUT33), .ZN(n682) );
  INV_X1 U742 ( .A(n682), .ZN(n677) );
  NAND2_X1 U743 ( .A1(G1976), .A2(G288), .ZN(n922) );
  INV_X1 U744 ( .A(KEYINPUT33), .ZN(n673) );
  NAND2_X1 U745 ( .A1(n922), .A2(n673), .ZN(n675) );
  NOR2_X1 U746 ( .A1(n675), .A2(n697), .ZN(n676) );
  OR2_X1 U747 ( .A1(n677), .A2(n676), .ZN(n679) );
  AND2_X1 U748 ( .A1(n690), .A2(n679), .ZN(n678) );
  NAND2_X1 U749 ( .A1(n689), .A2(n678), .ZN(n686) );
  INV_X1 U750 ( .A(n679), .ZN(n684) );
  NOR2_X1 U751 ( .A1(G1971), .A2(G303), .ZN(n680) );
  NOR2_X1 U752 ( .A1(n681), .A2(n680), .ZN(n933) );
  AND2_X1 U753 ( .A1(n933), .A2(n682), .ZN(n683) );
  OR2_X1 U754 ( .A1(n684), .A2(n683), .ZN(n685) );
  NAND2_X1 U755 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U756 ( .A(n687), .B(KEYINPUT100), .ZN(n688) );
  XOR2_X1 U757 ( .A(G1981), .B(G305), .Z(n941) );
  NAND2_X1 U758 ( .A1(n688), .A2(n941), .ZN(n701) );
  NAND2_X1 U759 ( .A1(n690), .A2(n689), .ZN(n693) );
  NOR2_X1 U760 ( .A1(G2090), .A2(G303), .ZN(n691) );
  NAND2_X1 U761 ( .A1(G8), .A2(n691), .ZN(n692) );
  NAND2_X1 U762 ( .A1(n693), .A2(n692), .ZN(n694) );
  AND2_X1 U763 ( .A1(n694), .A2(n697), .ZN(n699) );
  NOR2_X1 U764 ( .A1(G1981), .A2(G305), .ZN(n695) );
  XOR2_X1 U765 ( .A(n695), .B(KEYINPUT24), .Z(n696) );
  NOR2_X1 U766 ( .A1(n697), .A2(n696), .ZN(n698) );
  NOR2_X1 U767 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U768 ( .A(n702), .B(KEYINPUT101), .ZN(n716) );
  XNOR2_X1 U769 ( .A(KEYINPUT37), .B(G2067), .ZN(n747) );
  NAND2_X1 U770 ( .A1(n885), .A2(G140), .ZN(n703) );
  XNOR2_X1 U771 ( .A(n703), .B(KEYINPUT92), .ZN(n705) );
  NAND2_X1 U772 ( .A1(G104), .A2(n886), .ZN(n704) );
  NAND2_X1 U773 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U774 ( .A(KEYINPUT34), .B(n706), .ZN(n711) );
  NAND2_X1 U775 ( .A1(G116), .A2(n889), .ZN(n708) );
  NAND2_X1 U776 ( .A1(G128), .A2(n890), .ZN(n707) );
  NAND2_X1 U777 ( .A1(n708), .A2(n707), .ZN(n709) );
  XOR2_X1 U778 ( .A(KEYINPUT35), .B(n709), .Z(n710) );
  NOR2_X1 U779 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U780 ( .A(KEYINPUT36), .B(n712), .ZN(n905) );
  NOR2_X1 U781 ( .A1(n747), .A2(n905), .ZN(n1001) );
  INV_X1 U782 ( .A(n713), .ZN(n714) );
  NOR2_X1 U783 ( .A1(n715), .A2(n714), .ZN(n750) );
  NAND2_X1 U784 ( .A1(n1001), .A2(n750), .ZN(n745) );
  NAND2_X1 U785 ( .A1(n716), .A2(n745), .ZN(n740) );
  INV_X1 U786 ( .A(n750), .ZN(n738) );
  XNOR2_X1 U787 ( .A(G1986), .B(G290), .ZN(n929) );
  NAND2_X1 U788 ( .A1(n886), .A2(G105), .ZN(n717) );
  XNOR2_X1 U789 ( .A(KEYINPUT38), .B(n717), .ZN(n722) );
  NAND2_X1 U790 ( .A1(G117), .A2(n889), .ZN(n719) );
  NAND2_X1 U791 ( .A1(G129), .A2(n890), .ZN(n718) );
  NAND2_X1 U792 ( .A1(n719), .A2(n718), .ZN(n720) );
  XOR2_X1 U793 ( .A(KEYINPUT96), .B(n720), .Z(n721) );
  NAND2_X1 U794 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U795 ( .A(n723), .B(KEYINPUT97), .ZN(n725) );
  NAND2_X1 U796 ( .A1(G141), .A2(n885), .ZN(n724) );
  NAND2_X1 U797 ( .A1(n725), .A2(n724), .ZN(n882) );
  NAND2_X1 U798 ( .A1(G1996), .A2(n882), .ZN(n736) );
  NAND2_X1 U799 ( .A1(n890), .A2(G119), .ZN(n733) );
  NAND2_X1 U800 ( .A1(G131), .A2(n885), .ZN(n727) );
  NAND2_X1 U801 ( .A1(G95), .A2(n886), .ZN(n726) );
  NAND2_X1 U802 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U803 ( .A(KEYINPUT94), .B(n728), .ZN(n731) );
  NAND2_X1 U804 ( .A1(G107), .A2(n889), .ZN(n729) );
  XNOR2_X1 U805 ( .A(KEYINPUT93), .B(n729), .ZN(n730) );
  NOR2_X1 U806 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U807 ( .A1(n733), .A2(n732), .ZN(n734) );
  XOR2_X1 U808 ( .A(KEYINPUT95), .B(n734), .Z(n897) );
  NAND2_X1 U809 ( .A1(G1991), .A2(n897), .ZN(n735) );
  NAND2_X1 U810 ( .A1(n736), .A2(n735), .ZN(n1002) );
  NOR2_X1 U811 ( .A1(n929), .A2(n1002), .ZN(n737) );
  NOR2_X1 U812 ( .A1(n738), .A2(n737), .ZN(n739) );
  NOR2_X1 U813 ( .A1(n740), .A2(n739), .ZN(n753) );
  NOR2_X1 U814 ( .A1(G1996), .A2(n882), .ZN(n1017) );
  NOR2_X1 U815 ( .A1(G1986), .A2(G290), .ZN(n741) );
  NOR2_X1 U816 ( .A1(G1991), .A2(n897), .ZN(n1006) );
  NOR2_X1 U817 ( .A1(n741), .A2(n1006), .ZN(n742) );
  NOR2_X1 U818 ( .A1(n1002), .A2(n742), .ZN(n743) );
  NOR2_X1 U819 ( .A1(n1017), .A2(n743), .ZN(n744) );
  XNOR2_X1 U820 ( .A(n744), .B(KEYINPUT39), .ZN(n746) );
  NAND2_X1 U821 ( .A1(n746), .A2(n745), .ZN(n748) );
  NAND2_X1 U822 ( .A1(n747), .A2(n905), .ZN(n1003) );
  NAND2_X1 U823 ( .A1(n748), .A2(n1003), .ZN(n749) );
  NAND2_X1 U824 ( .A1(n750), .A2(n749), .ZN(n751) );
  XOR2_X1 U825 ( .A(KEYINPUT102), .B(n751), .Z(n752) );
  NOR2_X1 U826 ( .A1(n753), .A2(n752), .ZN(n755) );
  XNOR2_X1 U827 ( .A(n755), .B(n754), .ZN(G329) );
  AND2_X1 U828 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U829 ( .A(G108), .ZN(G238) );
  INV_X1 U830 ( .A(G132), .ZN(G219) );
  INV_X1 U831 ( .A(G82), .ZN(G220) );
  NOR2_X1 U832 ( .A1(n757), .A2(n756), .ZN(G160) );
  NAND2_X1 U833 ( .A1(G7), .A2(G661), .ZN(n758) );
  XNOR2_X1 U834 ( .A(n758), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U835 ( .A(KEYINPUT70), .B(KEYINPUT11), .Z(n760) );
  INV_X1 U836 ( .A(G223), .ZN(n828) );
  NAND2_X1 U837 ( .A1(G567), .A2(n828), .ZN(n759) );
  XNOR2_X1 U838 ( .A(n760), .B(n759), .ZN(G234) );
  INV_X1 U839 ( .A(G860), .ZN(n787) );
  OR2_X1 U840 ( .A1(n930), .A2(n787), .ZN(G153) );
  INV_X1 U841 ( .A(G301), .ZN(G171) );
  NAND2_X1 U842 ( .A1(G868), .A2(G171), .ZN(n762) );
  INV_X1 U843 ( .A(n934), .ZN(n785) );
  INV_X1 U844 ( .A(G868), .ZN(n765) );
  NAND2_X1 U845 ( .A1(n785), .A2(n765), .ZN(n761) );
  NAND2_X1 U846 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U847 ( .A(n763), .B(KEYINPUT73), .ZN(G284) );
  NOR2_X1 U848 ( .A1(G868), .A2(G299), .ZN(n764) );
  XNOR2_X1 U849 ( .A(n764), .B(KEYINPUT76), .ZN(n767) );
  NOR2_X1 U850 ( .A1(n765), .A2(G286), .ZN(n766) );
  NOR2_X1 U851 ( .A1(n767), .A2(n766), .ZN(G297) );
  NAND2_X1 U852 ( .A1(n787), .A2(G559), .ZN(n768) );
  NAND2_X1 U853 ( .A1(n768), .A2(n785), .ZN(n769) );
  XNOR2_X1 U854 ( .A(n769), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U855 ( .A1(G868), .A2(n930), .ZN(n770) );
  XOR2_X1 U856 ( .A(KEYINPUT77), .B(n770), .Z(n773) );
  NAND2_X1 U857 ( .A1(G868), .A2(n785), .ZN(n771) );
  NOR2_X1 U858 ( .A1(G559), .A2(n771), .ZN(n772) );
  NOR2_X1 U859 ( .A1(n773), .A2(n772), .ZN(G282) );
  NAND2_X1 U860 ( .A1(G99), .A2(n886), .ZN(n774) );
  XNOR2_X1 U861 ( .A(n774), .B(KEYINPUT78), .ZN(n781) );
  NAND2_X1 U862 ( .A1(G111), .A2(n889), .ZN(n776) );
  NAND2_X1 U863 ( .A1(G135), .A2(n885), .ZN(n775) );
  NAND2_X1 U864 ( .A1(n776), .A2(n775), .ZN(n779) );
  NAND2_X1 U865 ( .A1(n890), .A2(G123), .ZN(n777) );
  XOR2_X1 U866 ( .A(KEYINPUT18), .B(n777), .Z(n778) );
  NOR2_X1 U867 ( .A1(n779), .A2(n778), .ZN(n780) );
  NAND2_X1 U868 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U869 ( .A(KEYINPUT79), .B(n782), .ZN(n1005) );
  XNOR2_X1 U870 ( .A(n1005), .B(G2096), .ZN(n784) );
  INV_X1 U871 ( .A(G2100), .ZN(n783) );
  NAND2_X1 U872 ( .A1(n784), .A2(n783), .ZN(G156) );
  NAND2_X1 U873 ( .A1(G559), .A2(n785), .ZN(n786) );
  XOR2_X1 U874 ( .A(n930), .B(n786), .Z(n807) );
  NAND2_X1 U875 ( .A1(n787), .A2(n807), .ZN(n800) );
  NAND2_X1 U876 ( .A1(G55), .A2(n788), .ZN(n791) );
  NAND2_X1 U877 ( .A1(G67), .A2(n789), .ZN(n790) );
  NAND2_X1 U878 ( .A1(n791), .A2(n790), .ZN(n792) );
  XNOR2_X1 U879 ( .A(n792), .B(KEYINPUT81), .ZN(n795) );
  NAND2_X1 U880 ( .A1(G93), .A2(n793), .ZN(n794) );
  NAND2_X1 U881 ( .A1(n795), .A2(n794), .ZN(n799) );
  NAND2_X1 U882 ( .A1(n796), .A2(G80), .ZN(n797) );
  XOR2_X1 U883 ( .A(KEYINPUT80), .B(n797), .Z(n798) );
  NOR2_X1 U884 ( .A1(n799), .A2(n798), .ZN(n809) );
  XOR2_X1 U885 ( .A(n800), .B(n809), .Z(G145) );
  INV_X1 U886 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U887 ( .A(G166), .B(n809), .ZN(n806) );
  XNOR2_X1 U888 ( .A(KEYINPUT19), .B(G305), .ZN(n801) );
  XNOR2_X1 U889 ( .A(n801), .B(G288), .ZN(n802) );
  XNOR2_X1 U890 ( .A(KEYINPUT85), .B(n802), .ZN(n804) );
  XNOR2_X1 U891 ( .A(G290), .B(n921), .ZN(n803) );
  XNOR2_X1 U892 ( .A(n804), .B(n803), .ZN(n805) );
  XNOR2_X1 U893 ( .A(n806), .B(n805), .ZN(n910) );
  XNOR2_X1 U894 ( .A(n807), .B(n910), .ZN(n808) );
  NAND2_X1 U895 ( .A1(n808), .A2(G868), .ZN(n811) );
  OR2_X1 U896 ( .A1(G868), .A2(n809), .ZN(n810) );
  NAND2_X1 U897 ( .A1(n811), .A2(n810), .ZN(G295) );
  NAND2_X1 U898 ( .A1(G2084), .A2(G2078), .ZN(n813) );
  XOR2_X1 U899 ( .A(KEYINPUT86), .B(KEYINPUT20), .Z(n812) );
  XNOR2_X1 U900 ( .A(n813), .B(n812), .ZN(n814) );
  NAND2_X1 U901 ( .A1(G2090), .A2(n814), .ZN(n815) );
  XNOR2_X1 U902 ( .A(KEYINPUT21), .B(n815), .ZN(n816) );
  NAND2_X1 U903 ( .A1(n816), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U904 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U905 ( .A1(G220), .A2(G219), .ZN(n817) );
  XNOR2_X1 U906 ( .A(KEYINPUT22), .B(n817), .ZN(n818) );
  NAND2_X1 U907 ( .A1(n818), .A2(G96), .ZN(n819) );
  NOR2_X1 U908 ( .A1(n819), .A2(G218), .ZN(n820) );
  XNOR2_X1 U909 ( .A(n820), .B(KEYINPUT87), .ZN(n832) );
  NAND2_X1 U910 ( .A1(n832), .A2(G2106), .ZN(n826) );
  NAND2_X1 U911 ( .A1(G120), .A2(G69), .ZN(n821) );
  XOR2_X1 U912 ( .A(KEYINPUT88), .B(n821), .Z(n822) );
  NAND2_X1 U913 ( .A1(G57), .A2(n822), .ZN(n823) );
  NOR2_X1 U914 ( .A1(G238), .A2(n823), .ZN(n824) );
  XNOR2_X1 U915 ( .A(KEYINPUT89), .B(n824), .ZN(n833) );
  NAND2_X1 U916 ( .A1(n833), .A2(G567), .ZN(n825) );
  NAND2_X1 U917 ( .A1(n826), .A2(n825), .ZN(n834) );
  NAND2_X1 U918 ( .A1(G483), .A2(G661), .ZN(n827) );
  NOR2_X1 U919 ( .A1(n834), .A2(n827), .ZN(n831) );
  NAND2_X1 U920 ( .A1(n831), .A2(G36), .ZN(G176) );
  NAND2_X1 U921 ( .A1(G2106), .A2(n828), .ZN(G217) );
  AND2_X1 U922 ( .A1(G15), .A2(G2), .ZN(n829) );
  NAND2_X1 U923 ( .A1(G661), .A2(n829), .ZN(G259) );
  NAND2_X1 U924 ( .A1(G3), .A2(G1), .ZN(n830) );
  NAND2_X1 U925 ( .A1(n831), .A2(n830), .ZN(G188) );
  XOR2_X1 U926 ( .A(G96), .B(KEYINPUT106), .Z(G221) );
  XNOR2_X1 U927 ( .A(G69), .B(KEYINPUT107), .ZN(G235) );
  INV_X1 U929 ( .A(G120), .ZN(G236) );
  INV_X1 U930 ( .A(G57), .ZN(G237) );
  NOR2_X1 U931 ( .A1(n833), .A2(n832), .ZN(G325) );
  INV_X1 U932 ( .A(G325), .ZN(G261) );
  INV_X1 U933 ( .A(n834), .ZN(G319) );
  XNOR2_X1 U934 ( .A(G2454), .B(G2427), .ZN(n843) );
  XNOR2_X1 U935 ( .A(G2430), .B(G2451), .ZN(n841) );
  XOR2_X1 U936 ( .A(G2435), .B(KEYINPUT104), .Z(n836) );
  XNOR2_X1 U937 ( .A(G2443), .B(G2438), .ZN(n835) );
  XNOR2_X1 U938 ( .A(n836), .B(n835), .ZN(n837) );
  XOR2_X1 U939 ( .A(n837), .B(G2446), .Z(n839) );
  XNOR2_X1 U940 ( .A(G1341), .B(G1348), .ZN(n838) );
  XNOR2_X1 U941 ( .A(n839), .B(n838), .ZN(n840) );
  XNOR2_X1 U942 ( .A(n841), .B(n840), .ZN(n842) );
  XNOR2_X1 U943 ( .A(n843), .B(n842), .ZN(n844) );
  NAND2_X1 U944 ( .A1(n844), .A2(G14), .ZN(n845) );
  XNOR2_X1 U945 ( .A(KEYINPUT105), .B(n845), .ZN(G401) );
  XOR2_X1 U946 ( .A(KEYINPUT42), .B(KEYINPUT43), .Z(n847) );
  XNOR2_X1 U947 ( .A(G2072), .B(G2678), .ZN(n846) );
  XNOR2_X1 U948 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U949 ( .A(n848), .B(G2100), .Z(n850) );
  XNOR2_X1 U950 ( .A(G2067), .B(G2090), .ZN(n849) );
  XNOR2_X1 U951 ( .A(n850), .B(n849), .ZN(n854) );
  XOR2_X1 U952 ( .A(G2096), .B(KEYINPUT108), .Z(n852) );
  XNOR2_X1 U953 ( .A(G2084), .B(G2078), .ZN(n851) );
  XNOR2_X1 U954 ( .A(n852), .B(n851), .ZN(n853) );
  XNOR2_X1 U955 ( .A(n854), .B(n853), .ZN(G227) );
  XOR2_X1 U956 ( .A(G1976), .B(G1971), .Z(n856) );
  XNOR2_X1 U957 ( .A(G1986), .B(G1961), .ZN(n855) );
  XNOR2_X1 U958 ( .A(n856), .B(n855), .ZN(n857) );
  XOR2_X1 U959 ( .A(n857), .B(G2474), .Z(n859) );
  XNOR2_X1 U960 ( .A(G1991), .B(G1996), .ZN(n858) );
  XNOR2_X1 U961 ( .A(n859), .B(n858), .ZN(n863) );
  XOR2_X1 U962 ( .A(KEYINPUT41), .B(G1981), .Z(n861) );
  XNOR2_X1 U963 ( .A(G1966), .B(G1956), .ZN(n860) );
  XNOR2_X1 U964 ( .A(n861), .B(n860), .ZN(n862) );
  XNOR2_X1 U965 ( .A(n863), .B(n862), .ZN(G229) );
  NAND2_X1 U966 ( .A1(G124), .A2(n890), .ZN(n864) );
  XNOR2_X1 U967 ( .A(n864), .B(KEYINPUT44), .ZN(n869) );
  NAND2_X1 U968 ( .A1(G112), .A2(n889), .ZN(n866) );
  NAND2_X1 U969 ( .A1(G100), .A2(n886), .ZN(n865) );
  NAND2_X1 U970 ( .A1(n866), .A2(n865), .ZN(n867) );
  XOR2_X1 U971 ( .A(KEYINPUT110), .B(n867), .Z(n868) );
  NAND2_X1 U972 ( .A1(n869), .A2(n868), .ZN(n872) );
  NAND2_X1 U973 ( .A1(G136), .A2(n885), .ZN(n870) );
  XNOR2_X1 U974 ( .A(KEYINPUT109), .B(n870), .ZN(n871) );
  NOR2_X1 U975 ( .A1(n872), .A2(n871), .ZN(G162) );
  XNOR2_X1 U976 ( .A(KEYINPUT45), .B(KEYINPUT112), .ZN(n877) );
  NAND2_X1 U977 ( .A1(n886), .A2(G106), .ZN(n875) );
  NAND2_X1 U978 ( .A1(n885), .A2(G142), .ZN(n873) );
  XOR2_X1 U979 ( .A(KEYINPUT111), .B(n873), .Z(n874) );
  NAND2_X1 U980 ( .A1(n875), .A2(n874), .ZN(n876) );
  XOR2_X1 U981 ( .A(n877), .B(n876), .Z(n881) );
  NAND2_X1 U982 ( .A1(G118), .A2(n889), .ZN(n879) );
  NAND2_X1 U983 ( .A1(G130), .A2(n890), .ZN(n878) );
  NAND2_X1 U984 ( .A1(n879), .A2(n878), .ZN(n880) );
  NOR2_X1 U985 ( .A1(n881), .A2(n880), .ZN(n904) );
  XNOR2_X1 U986 ( .A(KEYINPUT48), .B(KEYINPUT113), .ZN(n884) );
  XNOR2_X1 U987 ( .A(n882), .B(KEYINPUT46), .ZN(n883) );
  XNOR2_X1 U988 ( .A(n884), .B(n883), .ZN(n899) );
  NAND2_X1 U989 ( .A1(G139), .A2(n885), .ZN(n888) );
  NAND2_X1 U990 ( .A1(G103), .A2(n886), .ZN(n887) );
  NAND2_X1 U991 ( .A1(n888), .A2(n887), .ZN(n895) );
  NAND2_X1 U992 ( .A1(G115), .A2(n889), .ZN(n892) );
  NAND2_X1 U993 ( .A1(G127), .A2(n890), .ZN(n891) );
  NAND2_X1 U994 ( .A1(n892), .A2(n891), .ZN(n893) );
  XOR2_X1 U995 ( .A(KEYINPUT47), .B(n893), .Z(n894) );
  NOR2_X1 U996 ( .A1(n895), .A2(n894), .ZN(n995) );
  XOR2_X1 U997 ( .A(G160), .B(n995), .Z(n896) );
  XNOR2_X1 U998 ( .A(n897), .B(n896), .ZN(n898) );
  XOR2_X1 U999 ( .A(n899), .B(n898), .Z(n901) );
  XNOR2_X1 U1000 ( .A(G164), .B(G162), .ZN(n900) );
  XNOR2_X1 U1001 ( .A(n901), .B(n900), .ZN(n902) );
  XNOR2_X1 U1002 ( .A(n1005), .B(n902), .ZN(n903) );
  XNOR2_X1 U1003 ( .A(n904), .B(n903), .ZN(n906) );
  XOR2_X1 U1004 ( .A(n906), .B(n905), .Z(n907) );
  NOR2_X1 U1005 ( .A1(G37), .A2(n907), .ZN(G395) );
  XNOR2_X1 U1006 ( .A(KEYINPUT114), .B(G301), .ZN(n908) );
  XNOR2_X1 U1007 ( .A(n908), .B(n930), .ZN(n909) );
  XNOR2_X1 U1008 ( .A(n910), .B(n909), .ZN(n912) );
  XNOR2_X1 U1009 ( .A(n934), .B(G286), .ZN(n911) );
  XNOR2_X1 U1010 ( .A(n912), .B(n911), .ZN(n913) );
  NOR2_X1 U1011 ( .A1(G37), .A2(n913), .ZN(G397) );
  NOR2_X1 U1012 ( .A1(G227), .A2(G229), .ZN(n914) );
  XNOR2_X1 U1013 ( .A(n914), .B(KEYINPUT49), .ZN(n915) );
  NOR2_X1 U1014 ( .A1(G401), .A2(n915), .ZN(n916) );
  NAND2_X1 U1015 ( .A1(G319), .A2(n916), .ZN(n917) );
  XNOR2_X1 U1016 ( .A(KEYINPUT115), .B(n917), .ZN(n919) );
  NOR2_X1 U1017 ( .A1(G395), .A2(G397), .ZN(n918) );
  NAND2_X1 U1018 ( .A1(n919), .A2(n918), .ZN(G225) );
  INV_X1 U1019 ( .A(G225), .ZN(G308) );
  XNOR2_X1 U1020 ( .A(G16), .B(KEYINPUT121), .ZN(n920) );
  XNOR2_X1 U1021 ( .A(n920), .B(KEYINPUT56), .ZN(n947) );
  XNOR2_X1 U1022 ( .A(n921), .B(G1956), .ZN(n923) );
  NAND2_X1 U1023 ( .A1(n923), .A2(n922), .ZN(n925) );
  XNOR2_X1 U1024 ( .A(G1961), .B(G301), .ZN(n924) );
  NOR2_X1 U1025 ( .A1(n925), .A2(n924), .ZN(n927) );
  NAND2_X1 U1026 ( .A1(G1971), .A2(G303), .ZN(n926) );
  NAND2_X1 U1027 ( .A1(n927), .A2(n926), .ZN(n928) );
  NOR2_X1 U1028 ( .A1(n929), .A2(n928), .ZN(n938) );
  XNOR2_X1 U1029 ( .A(G1341), .B(KEYINPUT123), .ZN(n931) );
  XNOR2_X1 U1030 ( .A(n931), .B(n930), .ZN(n932) );
  NAND2_X1 U1031 ( .A1(n933), .A2(n932), .ZN(n936) );
  XNOR2_X1 U1032 ( .A(G1348), .B(n934), .ZN(n935) );
  NOR2_X1 U1033 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1034 ( .A1(n938), .A2(n937), .ZN(n944) );
  XNOR2_X1 U1035 ( .A(G1966), .B(G168), .ZN(n939) );
  XNOR2_X1 U1036 ( .A(n939), .B(KEYINPUT122), .ZN(n940) );
  NAND2_X1 U1037 ( .A1(n941), .A2(n940), .ZN(n942) );
  XOR2_X1 U1038 ( .A(KEYINPUT57), .B(n942), .Z(n943) );
  NOR2_X1 U1039 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1040 ( .A(n945), .B(KEYINPUT124), .ZN(n946) );
  NOR2_X1 U1041 ( .A1(n947), .A2(n946), .ZN(n1028) );
  XNOR2_X1 U1042 ( .A(G16), .B(KEYINPUT125), .ZN(n971) );
  XNOR2_X1 U1043 ( .A(G20), .B(n948), .ZN(n952) );
  XNOR2_X1 U1044 ( .A(G1341), .B(G19), .ZN(n950) );
  XNOR2_X1 U1045 ( .A(G1981), .B(G6), .ZN(n949) );
  NOR2_X1 U1046 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1047 ( .A1(n952), .A2(n951), .ZN(n955) );
  XOR2_X1 U1048 ( .A(KEYINPUT59), .B(G1348), .Z(n953) );
  XNOR2_X1 U1049 ( .A(G4), .B(n953), .ZN(n954) );
  NOR2_X1 U1050 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1051 ( .A(KEYINPUT60), .B(n956), .ZN(n960) );
  XNOR2_X1 U1052 ( .A(G1966), .B(G21), .ZN(n958) );
  XNOR2_X1 U1053 ( .A(G5), .B(G1961), .ZN(n957) );
  NOR2_X1 U1054 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1055 ( .A1(n960), .A2(n959), .ZN(n967) );
  XNOR2_X1 U1056 ( .A(G1986), .B(G24), .ZN(n962) );
  XNOR2_X1 U1057 ( .A(G1971), .B(G22), .ZN(n961) );
  NOR2_X1 U1058 ( .A1(n962), .A2(n961), .ZN(n964) );
  XOR2_X1 U1059 ( .A(G1976), .B(G23), .Z(n963) );
  NAND2_X1 U1060 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1061 ( .A(KEYINPUT58), .B(n965), .ZN(n966) );
  NOR2_X1 U1062 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1063 ( .A(n968), .B(KEYINPUT61), .ZN(n969) );
  XNOR2_X1 U1064 ( .A(n969), .B(KEYINPUT126), .ZN(n970) );
  NAND2_X1 U1065 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1066 ( .A(n972), .B(KEYINPUT127), .ZN(n994) );
  XOR2_X1 U1067 ( .A(G29), .B(KEYINPUT120), .Z(n991) );
  XOR2_X1 U1068 ( .A(G1991), .B(G25), .Z(n973) );
  NAND2_X1 U1069 ( .A1(n973), .A2(G28), .ZN(n982) );
  XNOR2_X1 U1070 ( .A(G1996), .B(G32), .ZN(n975) );
  XNOR2_X1 U1071 ( .A(G33), .B(G2072), .ZN(n974) );
  NOR2_X1 U1072 ( .A1(n975), .A2(n974), .ZN(n980) );
  XNOR2_X1 U1073 ( .A(G2067), .B(G26), .ZN(n978) );
  XNOR2_X1 U1074 ( .A(G27), .B(n976), .ZN(n977) );
  NOR2_X1 U1075 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1076 ( .A1(n980), .A2(n979), .ZN(n981) );
  NOR2_X1 U1077 ( .A1(n982), .A2(n981), .ZN(n983) );
  XOR2_X1 U1078 ( .A(KEYINPUT53), .B(n983), .Z(n986) );
  XOR2_X1 U1079 ( .A(KEYINPUT54), .B(G34), .Z(n984) );
  XNOR2_X1 U1080 ( .A(G2084), .B(n984), .ZN(n985) );
  NAND2_X1 U1081 ( .A1(n986), .A2(n985), .ZN(n988) );
  XNOR2_X1 U1082 ( .A(G35), .B(G2090), .ZN(n987) );
  NOR2_X1 U1083 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1084 ( .A(n989), .B(KEYINPUT55), .ZN(n990) );
  NAND2_X1 U1085 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1086 ( .A1(G11), .A2(n992), .ZN(n993) );
  NOR2_X1 U1087 ( .A1(n994), .A2(n993), .ZN(n1026) );
  XNOR2_X1 U1088 ( .A(G164), .B(G2078), .ZN(n998) );
  XOR2_X1 U1089 ( .A(G2072), .B(n995), .Z(n996) );
  XNOR2_X1 U1090 ( .A(KEYINPUT119), .B(n996), .ZN(n997) );
  NAND2_X1 U1091 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1092 ( .A(n999), .B(KEYINPUT50), .ZN(n1000) );
  NOR2_X1 U1093 ( .A1(n1001), .A2(n1000), .ZN(n1014) );
  INV_X1 U1094 ( .A(n1002), .ZN(n1004) );
  NAND2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1012) );
  NOR2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XOR2_X1 U1097 ( .A(KEYINPUT116), .B(n1007), .Z(n1009) );
  XOR2_X1 U1098 ( .A(G160), .B(G2084), .Z(n1008) );
  NOR2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1100 ( .A(n1010), .B(KEYINPUT117), .ZN(n1011) );
  NOR2_X1 U1101 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1102 ( .A1(n1014), .A2(n1013), .ZN(n1020) );
  XOR2_X1 U1103 ( .A(G2090), .B(G162), .Z(n1015) );
  XNOR2_X1 U1104 ( .A(KEYINPUT118), .B(n1015), .ZN(n1016) );
  NOR2_X1 U1105 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1106 ( .A(KEYINPUT51), .B(n1018), .ZN(n1019) );
  NOR2_X1 U1107 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1108 ( .A(KEYINPUT52), .B(n1021), .ZN(n1023) );
  INV_X1 U1109 ( .A(KEYINPUT55), .ZN(n1022) );
  NAND2_X1 U1110 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1111 ( .A1(n1024), .A2(G29), .ZN(n1025) );
  NAND2_X1 U1112 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NOR2_X1 U1113 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XNOR2_X1 U1114 ( .A(n1029), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1115 ( .A(G311), .ZN(G150) );
endmodule

