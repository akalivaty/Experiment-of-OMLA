

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588;

  XNOR2_X1 U328 ( .A(n361), .B(n360), .ZN(n366) );
  AND2_X1 U329 ( .A1(G232GAT), .A2(G233GAT), .ZN(n296) );
  XOR2_X1 U330 ( .A(G190GAT), .B(G106GAT), .Z(n297) );
  XNOR2_X1 U331 ( .A(n359), .B(n296), .ZN(n360) );
  XNOR2_X1 U332 ( .A(n434), .B(n297), .ZN(n367) );
  XNOR2_X1 U333 ( .A(n368), .B(n367), .ZN(n369) );
  INV_X1 U334 ( .A(G190GAT), .ZN(n452) );
  XOR2_X1 U335 ( .A(n354), .B(n353), .Z(n518) );
  XNOR2_X1 U336 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U337 ( .A(n455), .B(n454), .ZN(G1351GAT) );
  XOR2_X1 U338 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n299) );
  XNOR2_X1 U339 ( .A(G190GAT), .B(KEYINPUT81), .ZN(n298) );
  XNOR2_X1 U340 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U341 ( .A(n300), .B(KEYINPUT19), .Z(n302) );
  XNOR2_X1 U342 ( .A(G169GAT), .B(G183GAT), .ZN(n301) );
  XNOR2_X1 U343 ( .A(n302), .B(n301), .ZN(n443) );
  XOR2_X1 U344 ( .A(G127GAT), .B(KEYINPUT78), .Z(n304) );
  XNOR2_X1 U345 ( .A(KEYINPUT0), .B(KEYINPUT77), .ZN(n303) );
  XNOR2_X1 U346 ( .A(n304), .B(n303), .ZN(n346) );
  XNOR2_X1 U347 ( .A(G99GAT), .B(G71GAT), .ZN(n305) );
  XNOR2_X1 U348 ( .A(n305), .B(G120GAT), .ZN(n415) );
  XNOR2_X1 U349 ( .A(n346), .B(n415), .ZN(n315) );
  XOR2_X1 U350 ( .A(KEYINPUT79), .B(KEYINPUT80), .Z(n307) );
  XNOR2_X1 U351 ( .A(KEYINPUT20), .B(KEYINPUT83), .ZN(n306) );
  XNOR2_X1 U352 ( .A(n307), .B(n306), .ZN(n311) );
  XOR2_X1 U353 ( .A(G176GAT), .B(KEYINPUT82), .Z(n309) );
  XOR2_X1 U354 ( .A(G113GAT), .B(G15GAT), .Z(n391) );
  XOR2_X1 U355 ( .A(G43GAT), .B(G134GAT), .Z(n364) );
  XNOR2_X1 U356 ( .A(n391), .B(n364), .ZN(n308) );
  XNOR2_X1 U357 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U358 ( .A(n311), .B(n310), .Z(n313) );
  NAND2_X1 U359 ( .A1(G227GAT), .A2(G233GAT), .ZN(n312) );
  XNOR2_X1 U360 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U361 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X2 U362 ( .A(n443), .B(n316), .ZN(n532) );
  XOR2_X1 U363 ( .A(KEYINPUT21), .B(KEYINPUT87), .Z(n318) );
  XNOR2_X1 U364 ( .A(KEYINPUT86), .B(G211GAT), .ZN(n317) );
  XNOR2_X1 U365 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U366 ( .A(G197GAT), .B(n319), .Z(n442) );
  XOR2_X1 U367 ( .A(KEYINPUT85), .B(KEYINPUT89), .Z(n321) );
  NAND2_X1 U368 ( .A1(G228GAT), .A2(G233GAT), .ZN(n320) );
  XNOR2_X1 U369 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U370 ( .A(n322), .B(G204GAT), .Z(n327) );
  XNOR2_X1 U371 ( .A(G106GAT), .B(G78GAT), .ZN(n323) );
  XNOR2_X1 U372 ( .A(n323), .B(G148GAT), .ZN(n409) );
  XOR2_X1 U373 ( .A(G155GAT), .B(KEYINPUT2), .Z(n325) );
  XNOR2_X1 U374 ( .A(KEYINPUT3), .B(KEYINPUT88), .ZN(n324) );
  XNOR2_X1 U375 ( .A(n325), .B(n324), .ZN(n350) );
  XNOR2_X1 U376 ( .A(n409), .B(n350), .ZN(n326) );
  XNOR2_X1 U377 ( .A(n327), .B(n326), .ZN(n331) );
  XOR2_X1 U378 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n329) );
  XNOR2_X1 U379 ( .A(G218GAT), .B(KEYINPUT22), .ZN(n328) );
  XNOR2_X1 U380 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U381 ( .A(n331), .B(n330), .Z(n333) );
  XOR2_X1 U382 ( .A(G141GAT), .B(G22GAT), .Z(n392) );
  XOR2_X1 U383 ( .A(G50GAT), .B(G162GAT), .Z(n359) );
  XNOR2_X1 U384 ( .A(n392), .B(n359), .ZN(n332) );
  XNOR2_X1 U385 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U386 ( .A(n442), .B(n334), .ZN(n465) );
  XOR2_X1 U387 ( .A(KEYINPUT6), .B(KEYINPUT4), .Z(n336) );
  XNOR2_X1 U388 ( .A(G1GAT), .B(KEYINPUT90), .ZN(n335) );
  XNOR2_X1 U389 ( .A(n336), .B(n335), .ZN(n354) );
  XOR2_X1 U390 ( .A(G162GAT), .B(G148GAT), .Z(n338) );
  XNOR2_X1 U391 ( .A(G29GAT), .B(G141GAT), .ZN(n337) );
  XNOR2_X1 U392 ( .A(n338), .B(n337), .ZN(n342) );
  XOR2_X1 U393 ( .A(KEYINPUT1), .B(G57GAT), .Z(n340) );
  XNOR2_X1 U394 ( .A(G113GAT), .B(G120GAT), .ZN(n339) );
  XNOR2_X1 U395 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U396 ( .A(n342), .B(n341), .Z(n348) );
  XOR2_X1 U397 ( .A(G85GAT), .B(G134GAT), .Z(n344) );
  NAND2_X1 U398 ( .A1(G225GAT), .A2(G233GAT), .ZN(n343) );
  XNOR2_X1 U399 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U400 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U401 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U402 ( .A(n349), .B(KEYINPUT91), .Z(n352) );
  XNOR2_X1 U403 ( .A(n350), .B(KEYINPUT5), .ZN(n351) );
  XNOR2_X1 U404 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U405 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n356) );
  XNOR2_X1 U406 ( .A(G99GAT), .B(KEYINPUT10), .ZN(n355) );
  XNOR2_X1 U407 ( .A(n356), .B(n355), .ZN(n370) );
  XOR2_X1 U408 ( .A(G85GAT), .B(KEYINPUT71), .Z(n357) );
  XNOR2_X1 U409 ( .A(KEYINPUT70), .B(n357), .ZN(n408) );
  INV_X1 U410 ( .A(n408), .ZN(n358) );
  XOR2_X1 U411 ( .A(G92GAT), .B(n358), .Z(n361) );
  XOR2_X1 U412 ( .A(G29GAT), .B(KEYINPUT8), .Z(n363) );
  XNOR2_X1 U413 ( .A(KEYINPUT7), .B(KEYINPUT67), .ZN(n362) );
  XNOR2_X1 U414 ( .A(n363), .B(n362), .ZN(n395) );
  XNOR2_X1 U415 ( .A(n395), .B(n364), .ZN(n365) );
  XNOR2_X1 U416 ( .A(n366), .B(n365), .ZN(n368) );
  XOR2_X1 U417 ( .A(G36GAT), .B(G218GAT), .Z(n434) );
  XNOR2_X1 U418 ( .A(n370), .B(n369), .ZN(n555) );
  XNOR2_X1 U419 ( .A(KEYINPUT36), .B(n555), .ZN(n584) );
  XOR2_X1 U420 ( .A(G155GAT), .B(G211GAT), .Z(n372) );
  XNOR2_X1 U421 ( .A(G183GAT), .B(G127GAT), .ZN(n371) );
  XNOR2_X1 U422 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U423 ( .A(G57GAT), .B(KEYINPUT13), .Z(n419) );
  XOR2_X1 U424 ( .A(n373), .B(n419), .Z(n375) );
  XNOR2_X1 U425 ( .A(G22GAT), .B(G78GAT), .ZN(n374) );
  XNOR2_X1 U426 ( .A(n375), .B(n374), .ZN(n380) );
  XNOR2_X1 U427 ( .A(G1GAT), .B(KEYINPUT68), .ZN(n376) );
  XNOR2_X1 U428 ( .A(n376), .B(G8GAT), .ZN(n393) );
  XOR2_X1 U429 ( .A(n393), .B(KEYINPUT12), .Z(n378) );
  NAND2_X1 U430 ( .A1(G231GAT), .A2(G233GAT), .ZN(n377) );
  XNOR2_X1 U431 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U432 ( .A(n380), .B(n379), .Z(n388) );
  XOR2_X1 U433 ( .A(KEYINPUT15), .B(KEYINPUT75), .Z(n382) );
  XNOR2_X1 U434 ( .A(G15GAT), .B(G71GAT), .ZN(n381) );
  XNOR2_X1 U435 ( .A(n382), .B(n381), .ZN(n386) );
  XOR2_X1 U436 ( .A(G64GAT), .B(KEYINPUT74), .Z(n384) );
  XNOR2_X1 U437 ( .A(KEYINPUT14), .B(KEYINPUT73), .ZN(n383) );
  XNOR2_X1 U438 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U439 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U440 ( .A(n388), .B(n387), .ZN(n582) );
  NAND2_X1 U441 ( .A1(n584), .A2(n582), .ZN(n390) );
  XOR2_X1 U442 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n389) );
  XNOR2_X1 U443 ( .A(n390), .B(n389), .ZN(n425) );
  XNOR2_X1 U444 ( .A(n392), .B(n391), .ZN(n394) );
  XNOR2_X1 U445 ( .A(n394), .B(n393), .ZN(n399) );
  XOR2_X1 U446 ( .A(n395), .B(KEYINPUT66), .Z(n397) );
  NAND2_X1 U447 ( .A1(G229GAT), .A2(G233GAT), .ZN(n396) );
  XNOR2_X1 U448 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U449 ( .A(n399), .B(n398), .Z(n407) );
  XOR2_X1 U450 ( .A(G197GAT), .B(G36GAT), .Z(n401) );
  XNOR2_X1 U451 ( .A(G43GAT), .B(G50GAT), .ZN(n400) );
  XNOR2_X1 U452 ( .A(n401), .B(n400), .ZN(n405) );
  XOR2_X1 U453 ( .A(KEYINPUT65), .B(KEYINPUT29), .Z(n403) );
  XNOR2_X1 U454 ( .A(G169GAT), .B(KEYINPUT30), .ZN(n402) );
  XNOR2_X1 U455 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U456 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U457 ( .A(n407), .B(n406), .ZN(n558) );
  INV_X1 U458 ( .A(n558), .ZN(n570) );
  XNOR2_X1 U459 ( .A(n409), .B(n408), .ZN(n423) );
  XOR2_X1 U460 ( .A(KEYINPUT33), .B(KEYINPUT72), .Z(n411) );
  NAND2_X1 U461 ( .A1(G230GAT), .A2(G233GAT), .ZN(n410) );
  XNOR2_X1 U462 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U463 ( .A(n412), .B(KEYINPUT69), .Z(n417) );
  XOR2_X1 U464 ( .A(G64GAT), .B(G92GAT), .Z(n414) );
  XNOR2_X1 U465 ( .A(G176GAT), .B(G204GAT), .ZN(n413) );
  XNOR2_X1 U466 ( .A(n414), .B(n413), .ZN(n435) );
  XNOR2_X1 U467 ( .A(n415), .B(n435), .ZN(n416) );
  XNOR2_X1 U468 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U469 ( .A(n418), .B(KEYINPUT32), .Z(n421) );
  XNOR2_X1 U470 ( .A(n419), .B(KEYINPUT31), .ZN(n420) );
  XNOR2_X1 U471 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U472 ( .A(n423), .B(n422), .Z(n576) );
  AND2_X1 U473 ( .A1(n570), .A2(n576), .ZN(n424) );
  NAND2_X1 U474 ( .A1(n425), .A2(n424), .ZN(n432) );
  XOR2_X1 U475 ( .A(KEYINPUT47), .B(KEYINPUT114), .Z(n430) );
  XNOR2_X1 U476 ( .A(n576), .B(KEYINPUT41), .ZN(n548) );
  NAND2_X1 U477 ( .A1(n558), .A2(n548), .ZN(n426) );
  XOR2_X1 U478 ( .A(KEYINPUT46), .B(n426), .Z(n427) );
  NOR2_X1 U479 ( .A1(n582), .A2(n427), .ZN(n428) );
  INV_X1 U480 ( .A(n555), .ZN(n456) );
  NAND2_X1 U481 ( .A1(n428), .A2(n456), .ZN(n429) );
  XNOR2_X1 U482 ( .A(n430), .B(n429), .ZN(n431) );
  NAND2_X1 U483 ( .A1(n432), .A2(n431), .ZN(n433) );
  XNOR2_X1 U484 ( .A(n433), .B(KEYINPUT48), .ZN(n544) );
  XOR2_X1 U485 ( .A(n435), .B(n434), .Z(n437) );
  NAND2_X1 U486 ( .A1(G226GAT), .A2(G233GAT), .ZN(n436) );
  XNOR2_X1 U487 ( .A(n437), .B(n436), .ZN(n441) );
  XOR2_X1 U488 ( .A(KEYINPUT92), .B(KEYINPUT93), .Z(n439) );
  XNOR2_X1 U489 ( .A(G8GAT), .B(KEYINPUT94), .ZN(n438) );
  XNOR2_X1 U490 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U491 ( .A(n441), .B(n440), .Z(n445) );
  XNOR2_X1 U492 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U493 ( .A(n445), .B(n444), .ZN(n504) );
  XOR2_X1 U494 ( .A(KEYINPUT119), .B(n504), .Z(n446) );
  NAND2_X1 U495 ( .A1(n544), .A2(n446), .ZN(n448) );
  XOR2_X1 U496 ( .A(KEYINPUT54), .B(KEYINPUT120), .Z(n447) );
  XNOR2_X1 U497 ( .A(n448), .B(n447), .ZN(n449) );
  NAND2_X1 U498 ( .A1(n518), .A2(n449), .ZN(n569) );
  NOR2_X1 U499 ( .A1(n465), .A2(n569), .ZN(n450) );
  XNOR2_X1 U500 ( .A(n450), .B(KEYINPUT55), .ZN(n451) );
  NOR2_X2 U501 ( .A1(n532), .A2(n451), .ZN(n565) );
  NAND2_X1 U502 ( .A1(n565), .A2(n555), .ZN(n455) );
  XOR2_X1 U503 ( .A(KEYINPUT122), .B(KEYINPUT58), .Z(n453) );
  XNOR2_X1 U504 ( .A(KEYINPUT34), .B(KEYINPUT100), .ZN(n478) );
  NAND2_X1 U505 ( .A1(n558), .A2(n576), .ZN(n490) );
  XOR2_X1 U506 ( .A(KEYINPUT76), .B(KEYINPUT16), .Z(n458) );
  NAND2_X1 U507 ( .A1(n582), .A2(n456), .ZN(n457) );
  XNOR2_X1 U508 ( .A(n458), .B(n457), .ZN(n474) );
  XNOR2_X1 U509 ( .A(n532), .B(KEYINPUT84), .ZN(n460) );
  XNOR2_X1 U510 ( .A(n504), .B(KEYINPUT27), .ZN(n463) );
  XOR2_X1 U511 ( .A(KEYINPUT28), .B(n465), .Z(n526) );
  NAND2_X1 U512 ( .A1(n463), .A2(n526), .ZN(n459) );
  NOR2_X1 U513 ( .A1(n518), .A2(n459), .ZN(n530) );
  NAND2_X1 U514 ( .A1(n460), .A2(n530), .ZN(n473) );
  NAND2_X1 U515 ( .A1(n465), .A2(n532), .ZN(n461) );
  XNOR2_X1 U516 ( .A(n461), .B(KEYINPUT95), .ZN(n462) );
  XNOR2_X1 U517 ( .A(KEYINPUT26), .B(n462), .ZN(n567) );
  NAND2_X1 U518 ( .A1(n463), .A2(n567), .ZN(n546) );
  XNOR2_X1 U519 ( .A(KEYINPUT96), .B(n546), .ZN(n469) );
  INV_X1 U520 ( .A(n504), .ZN(n521) );
  NOR2_X1 U521 ( .A1(n532), .A2(n521), .ZN(n464) );
  NOR2_X1 U522 ( .A1(n465), .A2(n464), .ZN(n466) );
  XOR2_X1 U523 ( .A(n466), .B(KEYINPUT97), .Z(n467) );
  XNOR2_X1 U524 ( .A(KEYINPUT25), .B(n467), .ZN(n468) );
  NAND2_X1 U525 ( .A1(n469), .A2(n468), .ZN(n470) );
  XNOR2_X1 U526 ( .A(KEYINPUT98), .B(n470), .ZN(n471) );
  NAND2_X1 U527 ( .A1(n471), .A2(n518), .ZN(n472) );
  NAND2_X1 U528 ( .A1(n473), .A2(n472), .ZN(n487) );
  NAND2_X1 U529 ( .A1(n474), .A2(n487), .ZN(n501) );
  OR2_X1 U530 ( .A1(n490), .A2(n501), .ZN(n484) );
  NOR2_X1 U531 ( .A1(n518), .A2(n484), .ZN(n476) );
  XNOR2_X1 U532 ( .A(G1GAT), .B(KEYINPUT99), .ZN(n475) );
  XNOR2_X1 U533 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U534 ( .A(n478), .B(n477), .ZN(G1324GAT) );
  NOR2_X1 U535 ( .A1(n521), .A2(n484), .ZN(n479) );
  XOR2_X1 U536 ( .A(G8GAT), .B(n479), .Z(G1325GAT) );
  NOR2_X1 U537 ( .A1(n484), .A2(n532), .ZN(n483) );
  XOR2_X1 U538 ( .A(KEYINPUT101), .B(KEYINPUT35), .Z(n481) );
  XNOR2_X1 U539 ( .A(G15GAT), .B(KEYINPUT102), .ZN(n480) );
  XNOR2_X1 U540 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U541 ( .A(n483), .B(n482), .ZN(G1326GAT) );
  NOR2_X1 U542 ( .A1(n526), .A2(n484), .ZN(n486) );
  XNOR2_X1 U543 ( .A(G22GAT), .B(KEYINPUT103), .ZN(n485) );
  XNOR2_X1 U544 ( .A(n486), .B(n485), .ZN(G1327GAT) );
  NAND2_X1 U545 ( .A1(n584), .A2(n487), .ZN(n488) );
  NOR2_X1 U546 ( .A1(n582), .A2(n488), .ZN(n489) );
  XNOR2_X1 U547 ( .A(KEYINPUT37), .B(n489), .ZN(n515) );
  NOR2_X1 U548 ( .A1(n515), .A2(n490), .ZN(n491) );
  XOR2_X1 U549 ( .A(KEYINPUT38), .B(n491), .Z(n497) );
  NOR2_X1 U550 ( .A1(n497), .A2(n518), .ZN(n492) );
  XNOR2_X1 U551 ( .A(n492), .B(KEYINPUT39), .ZN(n493) );
  XNOR2_X1 U552 ( .A(G29GAT), .B(n493), .ZN(G1328GAT) );
  NOR2_X1 U553 ( .A1(n497), .A2(n521), .ZN(n494) );
  XOR2_X1 U554 ( .A(G36GAT), .B(n494), .Z(G1329GAT) );
  NOR2_X1 U555 ( .A1(n497), .A2(n532), .ZN(n495) );
  XOR2_X1 U556 ( .A(KEYINPUT40), .B(n495), .Z(n496) );
  XNOR2_X1 U557 ( .A(G43GAT), .B(n496), .ZN(G1330GAT) );
  NOR2_X1 U558 ( .A1(n497), .A2(n526), .ZN(n498) );
  XOR2_X1 U559 ( .A(KEYINPUT104), .B(n498), .Z(n499) );
  XNOR2_X1 U560 ( .A(G50GAT), .B(n499), .ZN(G1331GAT) );
  XNOR2_X1 U561 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n503) );
  XOR2_X1 U562 ( .A(KEYINPUT105), .B(n548), .Z(n561) );
  NAND2_X1 U563 ( .A1(n561), .A2(n570), .ZN(n500) );
  XNOR2_X1 U564 ( .A(n500), .B(KEYINPUT106), .ZN(n516) );
  NOR2_X1 U565 ( .A1(n516), .A2(n501), .ZN(n510) );
  INV_X1 U566 ( .A(n518), .ZN(n543) );
  NAND2_X1 U567 ( .A1(n510), .A2(n543), .ZN(n502) );
  XNOR2_X1 U568 ( .A(n503), .B(n502), .ZN(G1332GAT) );
  XOR2_X1 U569 ( .A(G64GAT), .B(KEYINPUT107), .Z(n506) );
  NAND2_X1 U570 ( .A1(n510), .A2(n504), .ZN(n505) );
  XNOR2_X1 U571 ( .A(n506), .B(n505), .ZN(G1333GAT) );
  INV_X1 U572 ( .A(n532), .ZN(n507) );
  NAND2_X1 U573 ( .A1(n507), .A2(n510), .ZN(n508) );
  XNOR2_X1 U574 ( .A(G71GAT), .B(n508), .ZN(G1334GAT) );
  XOR2_X1 U575 ( .A(G78GAT), .B(KEYINPUT108), .Z(n512) );
  INV_X1 U576 ( .A(n526), .ZN(n509) );
  NAND2_X1 U577 ( .A1(n510), .A2(n509), .ZN(n511) );
  XNOR2_X1 U578 ( .A(n512), .B(n511), .ZN(n514) );
  XOR2_X1 U579 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n513) );
  XNOR2_X1 U580 ( .A(n514), .B(n513), .ZN(G1335GAT) );
  XNOR2_X1 U581 ( .A(G85GAT), .B(KEYINPUT111), .ZN(n520) );
  NOR2_X1 U582 ( .A1(n516), .A2(n515), .ZN(n517) );
  XOR2_X1 U583 ( .A(KEYINPUT110), .B(n517), .Z(n527) );
  NOR2_X1 U584 ( .A1(n518), .A2(n527), .ZN(n519) );
  XNOR2_X1 U585 ( .A(n520), .B(n519), .ZN(G1336GAT) );
  NOR2_X1 U586 ( .A1(n527), .A2(n521), .ZN(n522) );
  XOR2_X1 U587 ( .A(KEYINPUT112), .B(n522), .Z(n523) );
  XNOR2_X1 U588 ( .A(G92GAT), .B(n523), .ZN(G1337GAT) );
  NOR2_X1 U589 ( .A1(n527), .A2(n532), .ZN(n525) );
  XNOR2_X1 U590 ( .A(G99GAT), .B(KEYINPUT113), .ZN(n524) );
  XNOR2_X1 U591 ( .A(n525), .B(n524), .ZN(G1338GAT) );
  NOR2_X1 U592 ( .A1(n527), .A2(n526), .ZN(n528) );
  XOR2_X1 U593 ( .A(KEYINPUT44), .B(n528), .Z(n529) );
  XNOR2_X1 U594 ( .A(G106GAT), .B(n529), .ZN(G1339GAT) );
  NAND2_X1 U595 ( .A1(n544), .A2(n530), .ZN(n531) );
  NOR2_X1 U596 ( .A1(n532), .A2(n531), .ZN(n539) );
  NAND2_X1 U597 ( .A1(n539), .A2(n558), .ZN(n533) );
  XNOR2_X1 U598 ( .A(n533), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U599 ( .A(G120GAT), .B(KEYINPUT49), .Z(n535) );
  NAND2_X1 U600 ( .A1(n539), .A2(n561), .ZN(n534) );
  XNOR2_X1 U601 ( .A(n535), .B(n534), .ZN(G1341GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT50), .B(KEYINPUT115), .Z(n537) );
  NAND2_X1 U603 ( .A1(n539), .A2(n582), .ZN(n536) );
  XNOR2_X1 U604 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U605 ( .A(G127GAT), .B(n538), .ZN(G1342GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT116), .B(KEYINPUT51), .Z(n541) );
  NAND2_X1 U607 ( .A1(n539), .A2(n555), .ZN(n540) );
  XNOR2_X1 U608 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U609 ( .A(G134GAT), .B(n542), .ZN(G1343GAT) );
  NAND2_X1 U610 ( .A1(n544), .A2(n543), .ZN(n545) );
  NOR2_X1 U611 ( .A1(n546), .A2(n545), .ZN(n554) );
  NAND2_X1 U612 ( .A1(n554), .A2(n558), .ZN(n547) );
  XNOR2_X1 U613 ( .A(n547), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n550) );
  NAND2_X1 U615 ( .A1(n554), .A2(n548), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U617 ( .A(G148GAT), .B(n551), .ZN(G1345GAT) );
  XOR2_X1 U618 ( .A(G155GAT), .B(KEYINPUT117), .Z(n553) );
  NAND2_X1 U619 ( .A1(n554), .A2(n582), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(G1346GAT) );
  NAND2_X1 U621 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n556), .B(KEYINPUT118), .ZN(n557) );
  XNOR2_X1 U623 ( .A(G162GAT), .B(n557), .ZN(G1347GAT) );
  NAND2_X1 U624 ( .A1(n565), .A2(n558), .ZN(n559) );
  XOR2_X1 U625 ( .A(KEYINPUT121), .B(n559), .Z(n560) );
  XNOR2_X1 U626 ( .A(G169GAT), .B(n560), .ZN(G1348GAT) );
  XOR2_X1 U627 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n563) );
  NAND2_X1 U628 ( .A1(n565), .A2(n561), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U630 ( .A(G176GAT), .B(n564), .ZN(G1349GAT) );
  NAND2_X1 U631 ( .A1(n565), .A2(n582), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n566), .B(G183GAT), .ZN(G1350GAT) );
  INV_X1 U633 ( .A(n567), .ZN(n568) );
  NOR2_X1 U634 ( .A1(n569), .A2(n568), .ZN(n585) );
  INV_X1 U635 ( .A(n585), .ZN(n577) );
  NOR2_X1 U636 ( .A1(n570), .A2(n577), .ZN(n575) );
  XOR2_X1 U637 ( .A(KEYINPUT60), .B(KEYINPUT124), .Z(n572) );
  XNOR2_X1 U638 ( .A(G197GAT), .B(KEYINPUT123), .ZN(n571) );
  XNOR2_X1 U639 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U640 ( .A(KEYINPUT59), .B(n573), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(G1352GAT) );
  NOR2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n581) );
  XOR2_X1 U643 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n579) );
  XNOR2_X1 U644 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1353GAT) );
  AND2_X1 U647 ( .A1(n582), .A2(n585), .ZN(n583) );
  XOR2_X1 U648 ( .A(G211GAT), .B(n583), .Z(G1354GAT) );
  XOR2_X1 U649 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n587) );
  NAND2_X1 U650 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n587), .B(n586), .ZN(n588) );
  XNOR2_X1 U652 ( .A(G218GAT), .B(n588), .ZN(G1355GAT) );
endmodule

