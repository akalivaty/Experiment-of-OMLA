//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 0 0 1 1 1 0 1 0 1 0 0 0 0 0 0 0 1 0 1 1 1 0 1 1 1 0 1 0 0 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 0 1 0 0 1 0 0 1 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:01 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1287, new_n1288, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(KEYINPUT64), .B(KEYINPUT0), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n210), .B(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n213));
  INV_X1    g0013(.A(G68), .ZN(new_n214));
  INV_X1    g0014(.A(G238), .ZN(new_n215));
  INV_X1    g0015(.A(G87), .ZN(new_n216));
  INV_X1    g0016(.A(G250), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n219));
  INV_X1    g0019(.A(G77), .ZN(new_n220));
  INV_X1    g0020(.A(G244), .ZN(new_n221));
  INV_X1    g0021(.A(G107), .ZN(new_n222));
  INV_X1    g0022(.A(G264), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n208), .B1(new_n218), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT1), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n227), .A2(new_n206), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n202), .A2(G50), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  AOI211_X1 g0030(.A(new_n212), .B(new_n226), .C1(new_n228), .C2(new_n230), .ZN(G361));
  XOR2_X1   g0031(.A(G238), .B(G244), .Z(new_n232));
  XNOR2_X1  g0032(.A(G226), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G58), .B(G77), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n241), .B(new_n242), .Z(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  AOI21_X1  g0047(.A(new_n227), .B1(G33), .B2(G41), .ZN(new_n248));
  INV_X1    g0048(.A(G274), .ZN(new_n249));
  OAI21_X1  g0049(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n250));
  NOR3_X1   g0050(.A1(new_n248), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(G33), .A2(G41), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n252), .A2(G1), .A3(G13), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(new_n250), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n251), .B1(G232), .B2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(KEYINPUT3), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  XNOR2_X1  g0059(.A(KEYINPUT74), .B(KEYINPUT3), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n259), .B1(new_n260), .B2(G33), .ZN(new_n261));
  NOR2_X1   g0061(.A1(G223), .A2(G1698), .ZN(new_n262));
  INV_X1    g0062(.A(G226), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n262), .B1(new_n263), .B2(G1698), .ZN(new_n264));
  AOI22_X1  g0064(.A1(new_n261), .A2(new_n264), .B1(G33), .B2(G87), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n256), .B1(new_n253), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G169), .ZN(new_n267));
  OAI211_X1 g0067(.A(new_n256), .B(G179), .C1(new_n253), .C2(new_n265), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g0069(.A(G58), .B(G68), .ZN(new_n270));
  NOR2_X1   g0070(.A1(G20), .A2(G33), .ZN(new_n271));
  AOI22_X1  g0071(.A1(new_n270), .A2(G20), .B1(G159), .B2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT3), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(KEYINPUT74), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT74), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(KEYINPUT3), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n274), .A2(new_n276), .A3(G33), .ZN(new_n277));
  AOI21_X1  g0077(.A(G20), .B1(new_n277), .B2(new_n258), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT7), .ZN(new_n279));
  OAI21_X1  g0079(.A(G68), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  XNOR2_X1  g0080(.A(KEYINPUT75), .B(KEYINPUT7), .ZN(new_n281));
  AOI211_X1 g0081(.A(G20), .B(new_n281), .C1(new_n277), .C2(new_n258), .ZN(new_n282));
  OAI211_X1 g0082(.A(KEYINPUT16), .B(new_n272), .C1(new_n280), .C2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n227), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT16), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n273), .A2(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n258), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n281), .B1(new_n206), .B2(new_n289), .ZN(new_n290));
  OAI21_X1  g0090(.A(KEYINPUT76), .B1(new_n260), .B2(G33), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT76), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n275), .A2(KEYINPUT3), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n273), .A2(KEYINPUT74), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n292), .B(new_n257), .C1(new_n293), .C2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT77), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n296), .B1(new_n257), .B2(KEYINPUT3), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n273), .A2(KEYINPUT77), .A3(G33), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n291), .A2(new_n295), .A3(new_n297), .A4(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n206), .A2(KEYINPUT7), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n290), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n272), .B1(new_n302), .B2(new_n214), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n286), .B1(new_n287), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G13), .ZN(new_n305));
  NOR3_X1   g0105(.A1(new_n305), .A2(new_n206), .A3(G1), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n306), .A2(new_n285), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  XNOR2_X1  g0108(.A(KEYINPUT8), .B(G58), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT68), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n311), .B1(new_n206), .B2(G1), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n205), .A2(KEYINPUT68), .A3(G20), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n310), .A2(new_n314), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n305), .A2(G1), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(G20), .ZN(new_n317));
  OAI22_X1  g0117(.A1(new_n308), .A2(new_n315), .B1(new_n317), .B2(new_n310), .ZN(new_n318));
  OAI211_X1 g0118(.A(KEYINPUT18), .B(new_n269), .C1(new_n304), .C2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(KEYINPUT78), .ZN(new_n320));
  INV_X1    g0120(.A(new_n318), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n297), .A2(new_n298), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n257), .B1(new_n293), .B2(new_n294), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n322), .B1(new_n323), .B2(KEYINPUT76), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n300), .B1(new_n324), .B2(new_n295), .ZN(new_n325));
  OAI21_X1  g0125(.A(G68), .B1(new_n325), .B2(new_n290), .ZN(new_n326));
  AOI21_X1  g0126(.A(KEYINPUT16), .B1(new_n326), .B2(new_n272), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n321), .B1(new_n327), .B2(new_n286), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT78), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n328), .A2(new_n329), .A3(KEYINPUT18), .A4(new_n269), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(new_n269), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT18), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n320), .A2(new_n330), .A3(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(G200), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n266), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(G190), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n256), .B(new_n337), .C1(new_n253), .C2(new_n265), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n321), .B(new_n339), .C1(new_n327), .C2(new_n286), .ZN(new_n340));
  XNOR2_X1  g0140(.A(new_n340), .B(KEYINPUT17), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n334), .A2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(G50), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n344), .B1(new_n312), .B2(new_n313), .ZN(new_n345));
  AOI22_X1  g0145(.A1(new_n307), .A2(new_n345), .B1(new_n344), .B2(new_n306), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n206), .B1(new_n201), .B2(new_n344), .ZN(new_n347));
  XNOR2_X1  g0147(.A(new_n347), .B(KEYINPUT67), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n206), .A2(G33), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  AOI22_X1  g0150(.A1(new_n310), .A2(new_n350), .B1(G150), .B2(new_n271), .ZN(new_n351));
  AND2_X1   g0151(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n285), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n346), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  XNOR2_X1  g0154(.A(new_n354), .B(KEYINPUT9), .ZN(new_n355));
  MUX2_X1   g0155(.A(G222), .B(G223), .S(G1698), .Z(new_n356));
  XNOR2_X1  g0156(.A(KEYINPUT3), .B(G33), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n358), .B1(new_n220), .B2(new_n357), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT66), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n253), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n361), .B1(new_n360), .B2(new_n359), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n251), .B1(G226), .B2(new_n255), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT71), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n364), .A2(G200), .B1(new_n365), .B2(KEYINPUT10), .ZN(new_n366));
  AND2_X1   g0166(.A1(new_n362), .A2(new_n363), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(G190), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n355), .A2(new_n366), .A3(new_n368), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n365), .A2(KEYINPUT10), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n370), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n355), .A2(new_n366), .A3(new_n368), .A4(new_n372), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n354), .B1(new_n367), .B2(G169), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n364), .A2(G179), .ZN(new_n375));
  OR2_X1    g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n371), .A2(new_n373), .A3(new_n376), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n310), .A2(new_n271), .B1(G20), .B2(G77), .ZN(new_n378));
  XNOR2_X1  g0178(.A(KEYINPUT15), .B(G87), .ZN(new_n379));
  OR2_X1    g0179(.A1(new_n379), .A2(new_n349), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n353), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n307), .A2(G77), .A3(new_n314), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n382), .B1(G77), .B2(new_n317), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n357), .A2(G238), .A3(G1698), .ZN(new_n385));
  INV_X1    g0185(.A(G1698), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n357), .A2(G232), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n222), .A2(KEYINPUT69), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT69), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(G107), .ZN(new_n390));
  AND2_X1   g0190(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  OAI211_X1 g0191(.A(new_n385), .B(new_n387), .C1(new_n391), .C2(new_n357), .ZN(new_n392));
  OR2_X1    g0192(.A1(new_n392), .A2(KEYINPUT70), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n253), .B1(new_n392), .B2(KEYINPUT70), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n251), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n396), .B1(new_n221), .B2(new_n254), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n395), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(G169), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n384), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n397), .B1(new_n393), .B2(new_n394), .ZN(new_n402));
  INV_X1    g0202(.A(G179), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n402), .A2(G190), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n406), .B(new_n384), .C1(new_n335), .C2(new_n402), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n377), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n306), .A2(new_n214), .ZN(new_n410));
  XNOR2_X1  g0210(.A(new_n410), .B(KEYINPUT12), .ZN(new_n411));
  AOI22_X1  g0211(.A1(new_n271), .A2(G50), .B1(G20), .B2(new_n214), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n412), .B1(new_n220), .B2(new_n349), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n413), .A2(KEYINPUT11), .A3(new_n285), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n307), .A2(G68), .A3(new_n314), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n411), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(KEYINPUT11), .B1(new_n413), .B2(new_n285), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT14), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n263), .A2(new_n386), .ZN(new_n421));
  OR2_X1    g0221(.A1(new_n386), .A2(G232), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n357), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(G33), .A2(G97), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n423), .A2(KEYINPUT72), .A3(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(KEYINPUT72), .B1(new_n423), .B2(new_n424), .ZN(new_n427));
  NOR3_X1   g0227(.A1(new_n426), .A2(new_n427), .A3(new_n253), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n251), .B1(G238), .B2(new_n255), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  NOR3_X1   g0230(.A1(new_n428), .A2(KEYINPUT13), .A3(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT13), .ZN(new_n432));
  INV_X1    g0232(.A(new_n427), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n433), .A2(new_n248), .A3(new_n425), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n432), .B1(new_n434), .B2(new_n429), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n420), .B(G169), .C1(new_n431), .C2(new_n435), .ZN(new_n436));
  OAI21_X1  g0236(.A(KEYINPUT13), .B1(new_n428), .B2(new_n430), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n434), .A2(new_n432), .A3(new_n429), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n437), .A2(new_n438), .A3(G179), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n437), .A2(new_n438), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n420), .B1(new_n441), .B2(G169), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n419), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n441), .A2(G200), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n437), .A2(new_n438), .A3(G190), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n444), .A2(new_n418), .A3(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(KEYINPUT73), .B1(new_n443), .B2(new_n446), .ZN(new_n447));
  AND3_X1   g0247(.A1(new_n443), .A2(KEYINPUT73), .A3(new_n446), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n343), .B(new_n409), .C1(new_n447), .C2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT86), .ZN(new_n451));
  INV_X1    g0251(.A(G257), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n452), .A2(new_n386), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n277), .A2(new_n451), .A3(new_n258), .A4(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(G33), .A2(G294), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n217), .A2(G1698), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n277), .A2(new_n258), .A3(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n454), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n451), .B1(new_n261), .B2(new_n453), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n248), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT87), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n277), .A2(new_n258), .A3(new_n453), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(KEYINPUT86), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n464), .A2(new_n454), .A3(new_n455), .A4(new_n457), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n465), .A2(KEYINPUT87), .A3(new_n248), .ZN(new_n466));
  XNOR2_X1  g0266(.A(KEYINPUT5), .B(G41), .ZN(new_n467));
  INV_X1    g0267(.A(G45), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n468), .A2(G1), .ZN(new_n469));
  AND2_X1   g0269(.A1(G1), .A2(G13), .ZN(new_n470));
  AOI22_X1  g0270(.A1(new_n467), .A2(new_n469), .B1(new_n470), .B2(new_n252), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(G264), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n205), .A2(G45), .ZN(new_n473));
  OR2_X1    g0273(.A1(KEYINPUT5), .A2(G41), .ZN(new_n474));
  NAND2_X1  g0274(.A1(KEYINPUT5), .A2(G41), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n249), .B1(new_n470), .B2(new_n252), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n472), .A2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n462), .A2(new_n337), .A3(new_n466), .A4(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n460), .A2(new_n480), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n335), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT83), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n388), .A2(new_n390), .A3(G20), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n485), .B1(new_n486), .B2(KEYINPUT23), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n216), .A2(G20), .ZN(new_n488));
  AOI21_X1  g0288(.A(KEYINPUT22), .B1(new_n357), .B2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT23), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n490), .A2(new_n222), .A3(G20), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n206), .A2(G33), .A3(G116), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NOR3_X1   g0293(.A1(new_n487), .A2(new_n489), .A3(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT24), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT22), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n496), .A2(new_n216), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n277), .A2(new_n206), .A3(new_n258), .A4(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n486), .A2(new_n485), .A3(KEYINPUT23), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n494), .A2(new_n495), .A3(new_n498), .A4(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n486), .A2(KEYINPUT23), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(KEYINPUT83), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n488), .A2(new_n258), .A3(new_n288), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n493), .B1(new_n496), .B2(new_n503), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n502), .A2(new_n504), .A3(new_n498), .A4(new_n499), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(KEYINPUT24), .ZN(new_n506));
  AND2_X1   g0306(.A1(new_n500), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g0307(.A(KEYINPUT84), .B1(new_n507), .B2(new_n353), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT25), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n316), .A2(new_n509), .A3(G20), .A4(new_n222), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n316), .A2(G20), .A3(new_n222), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(KEYINPUT25), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n205), .A2(G33), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n353), .A2(new_n317), .A3(new_n513), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n510), .B(new_n512), .C1(new_n514), .C2(new_n222), .ZN(new_n515));
  XNOR2_X1  g0315(.A(new_n515), .B(KEYINPUT85), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n353), .B1(new_n500), .B2(new_n506), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT84), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  AND3_X1   g0319(.A1(new_n484), .A2(new_n508), .A3(new_n519), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n480), .B1(new_n460), .B2(new_n461), .ZN(new_n521));
  AOI21_X1  g0321(.A(KEYINPUT87), .B1(new_n465), .B2(new_n248), .ZN(new_n522));
  OAI21_X1  g0322(.A(G169), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n479), .B1(new_n465), .B2(new_n248), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(G179), .ZN(new_n525));
  AOI22_X1  g0325(.A1(new_n508), .A2(new_n519), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  OAI21_X1  g0326(.A(KEYINPUT88), .B1(new_n520), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n508), .A2(new_n519), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n523), .A2(new_n525), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT88), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n484), .A2(new_n508), .A3(new_n519), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT21), .ZN(new_n534));
  NAND2_X1  g0334(.A1(G33), .A2(G283), .ZN(new_n535));
  INV_X1    g0335(.A(G97), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n535), .B(new_n206), .C1(G33), .C2(new_n536), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n537), .B(new_n285), .C1(new_n206), .C2(G116), .ZN(new_n538));
  XNOR2_X1  g0338(.A(new_n538), .B(KEYINPUT20), .ZN(new_n539));
  INV_X1    g0339(.A(G116), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n306), .A2(new_n540), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n541), .B1(new_n514), .B2(new_n540), .ZN(new_n542));
  OAI21_X1  g0342(.A(G169), .B1(new_n539), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g0343(.A1(G257), .A2(G1698), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n544), .B1(new_n223), .B2(G1698), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n545), .A2(new_n277), .A3(new_n258), .ZN(new_n546));
  INV_X1    g0346(.A(G303), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(KEYINPUT82), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT82), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(G303), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n289), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n253), .B1(new_n546), .B2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(new_n475), .ZN(new_n554));
  NOR2_X1   g0354(.A1(KEYINPUT5), .A2(G41), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n469), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n253), .ZN(new_n557));
  INV_X1    g0357(.A(G270), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n478), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n553), .A2(new_n559), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n534), .B1(new_n543), .B2(new_n560), .ZN(new_n561));
  OR2_X1    g0361(.A1(new_n539), .A2(new_n542), .ZN(new_n562));
  AOI22_X1  g0362(.A1(new_n471), .A2(G270), .B1(new_n476), .B2(new_n477), .ZN(new_n563));
  AOI22_X1  g0363(.A1(new_n258), .A2(new_n288), .B1(new_n548), .B2(new_n550), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n564), .B1(new_n261), .B2(new_n545), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n563), .B1(new_n565), .B2(new_n253), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n562), .A2(KEYINPUT21), .A3(G169), .A4(new_n566), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n539), .A2(new_n542), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n563), .B(G179), .C1(new_n565), .C2(new_n253), .ZN(new_n569));
  OR2_X1    g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n560), .A2(G190), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n571), .B(new_n568), .C1(new_n335), .C2(new_n560), .ZN(new_n572));
  AND4_X1   g0372(.A1(new_n561), .A2(new_n567), .A3(new_n570), .A4(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n514), .A2(G97), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n317), .A2(new_n536), .ZN(new_n575));
  AND3_X1   g0375(.A1(new_n574), .A2(KEYINPUT79), .A3(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(KEYINPUT79), .B1(new_n574), .B2(new_n575), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n222), .A2(KEYINPUT6), .A3(G97), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n536), .A2(new_n222), .ZN(new_n580));
  NOR2_X1   g0380(.A1(G97), .A2(G107), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n579), .B1(new_n582), .B2(KEYINPUT6), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n583), .A2(G20), .B1(G77), .B2(new_n271), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n584), .B1(new_n302), .B2(new_n391), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n578), .B1(new_n585), .B2(new_n285), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n221), .A2(G1698), .ZN(new_n587));
  AOI21_X1  g0387(.A(KEYINPUT4), .B1(new_n261), .B2(new_n587), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n258), .A2(new_n288), .A3(G250), .A4(G1698), .ZN(new_n589));
  AND2_X1   g0389(.A1(KEYINPUT4), .A2(G244), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n258), .A2(new_n288), .A3(new_n590), .A4(new_n386), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n589), .A2(new_n591), .A3(new_n535), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n248), .B1(new_n588), .B2(new_n592), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n478), .B1(new_n557), .B2(new_n452), .ZN(new_n594));
  INV_X1    g0394(.A(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n593), .A2(new_n403), .A3(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT4), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n277), .A2(new_n258), .ZN(new_n598));
  INV_X1    g0398(.A(new_n587), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n597), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(new_n592), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n594), .B1(new_n602), .B2(new_n248), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n596), .B1(new_n603), .B2(G169), .ZN(new_n604));
  OR2_X1    g0404(.A1(new_n586), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n603), .A2(new_n337), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n606), .B1(G200), .B2(new_n603), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n586), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n277), .A2(new_n206), .A3(G68), .A4(new_n258), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT19), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n388), .A2(new_n390), .A3(new_n216), .A4(new_n536), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n424), .A2(new_n206), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NOR3_X1   g0413(.A1(new_n349), .A2(KEYINPUT19), .A3(new_n536), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n609), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n285), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n379), .A2(new_n306), .ZN(new_n617));
  XNOR2_X1  g0417(.A(new_n379), .B(KEYINPUT81), .ZN(new_n618));
  INV_X1    g0418(.A(new_n514), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n616), .A2(new_n617), .A3(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n253), .A2(G250), .A3(new_n473), .ZN(new_n622));
  INV_X1    g0422(.A(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n253), .A2(G274), .A3(new_n469), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT80), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n477), .A2(KEYINPUT80), .A3(new_n469), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n623), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NOR2_X1   g0428(.A1(G238), .A2(G1698), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n629), .B1(new_n221), .B2(G1698), .ZN(new_n630));
  AOI22_X1  g0430(.A1(new_n261), .A2(new_n630), .B1(G33), .B2(G116), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n628), .B1(new_n631), .B2(new_n253), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n400), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n628), .B(new_n403), .C1(new_n631), .C2(new_n253), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n621), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  AOI22_X1  g0435(.A1(new_n615), .A2(new_n285), .B1(new_n306), .B2(new_n379), .ZN(new_n636));
  AOI21_X1  g0436(.A(KEYINPUT80), .B1(new_n477), .B2(new_n469), .ZN(new_n637));
  AND4_X1   g0437(.A1(KEYINPUT80), .A2(new_n253), .A3(G274), .A4(new_n469), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n622), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n630), .A2(new_n277), .A3(new_n258), .ZN(new_n640));
  NAND2_X1  g0440(.A1(G33), .A2(G116), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n253), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(G200), .B1(new_n639), .B2(new_n642), .ZN(new_n643));
  OAI211_X1 g0443(.A(new_n628), .B(G190), .C1(new_n631), .C2(new_n253), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n619), .A2(G87), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n636), .A2(new_n643), .A3(new_n644), .A4(new_n645), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n635), .A2(new_n646), .ZN(new_n647));
  AND4_X1   g0447(.A1(new_n573), .A2(new_n605), .A3(new_n608), .A4(new_n647), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n450), .A2(new_n527), .A3(new_n533), .A4(new_n648), .ZN(new_n649));
  XOR2_X1   g0449(.A(new_n649), .B(KEYINPUT89), .Z(G372));
  NAND2_X1  g0450(.A1(new_n371), .A2(new_n373), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n446), .A2(new_n404), .A3(new_n401), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n443), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(new_n341), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n333), .A2(new_n319), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT91), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n651), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n654), .A2(KEYINPUT91), .A3(new_n655), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n660), .A2(new_n376), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n567), .A2(new_n561), .A3(new_n570), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n530), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n586), .A2(new_n604), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n665), .B1(new_n586), .B2(new_n607), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n664), .A2(new_n532), .A3(new_n666), .A4(new_n647), .ZN(new_n667));
  XNOR2_X1  g0467(.A(new_n635), .B(KEYINPUT90), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT26), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n635), .A2(new_n646), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n669), .B1(new_n605), .B2(new_n670), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n665), .A2(new_n647), .A3(KEYINPUT26), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n668), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n667), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n661), .B1(new_n449), .B2(new_n675), .ZN(G369));
  NAND2_X1  g0476(.A1(new_n316), .A2(new_n206), .ZN(new_n677));
  OR2_X1    g0477(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n678), .A2(G213), .A3(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(G343), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n528), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n527), .A2(new_n533), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(KEYINPUT92), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT92), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n527), .A2(new_n533), .A3(new_n686), .A4(new_n683), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n682), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n688), .B1(new_n530), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n562), .A2(new_n682), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n573), .A2(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n692), .B1(new_n663), .B2(new_n691), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(G330), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n690), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n663), .A2(new_n682), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n685), .A2(new_n687), .A3(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT94), .ZN(new_n699));
  XOR2_X1   g0499(.A(new_n682), .B(KEYINPUT93), .Z(new_n700));
  NAND2_X1  g0500(.A1(new_n526), .A2(new_n700), .ZN(new_n701));
  AND3_X1   g0501(.A1(new_n698), .A2(new_n699), .A3(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n699), .B1(new_n698), .B2(new_n701), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n696), .B1(new_n702), .B2(new_n703), .ZN(G399));
  INV_X1    g0504(.A(new_n209), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(G41), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n611), .A2(G116), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NOR3_X1   g0508(.A1(new_n706), .A2(new_n205), .A3(new_n708), .ZN(new_n709));
  AOI22_X1  g0509(.A1(new_n709), .A2(KEYINPUT95), .B1(new_n230), .B2(new_n706), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n710), .B1(KEYINPUT95), .B2(new_n709), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n711), .B(KEYINPUT28), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n682), .B1(new_n667), .B2(new_n673), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(KEYINPUT29), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n532), .A2(new_n605), .A3(new_n608), .A4(new_n647), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n662), .B1(new_n528), .B2(new_n529), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n668), .ZN(new_n718));
  AOI21_X1  g0518(.A(KEYINPUT26), .B1(new_n665), .B2(new_n647), .ZN(new_n719));
  NOR4_X1   g0519(.A1(new_n670), .A2(new_n586), .A3(new_n604), .A4(new_n669), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n718), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n700), .B1(new_n717), .B2(new_n721), .ZN(new_n722));
  XNOR2_X1  g0522(.A(KEYINPUT97), .B(KEYINPUT29), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n714), .A2(new_n724), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n648), .A2(new_n527), .A3(new_n533), .A4(new_n700), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT31), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n632), .A2(new_n566), .A3(new_n403), .ZN(new_n728));
  NOR3_X1   g0528(.A1(new_n728), .A2(new_n524), .A3(new_n603), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n639), .A2(new_n642), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n730), .A2(new_n560), .A3(G179), .A4(new_n472), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n460), .A2(new_n593), .A3(new_n595), .ZN(new_n732));
  OAI21_X1  g0532(.A(KEYINPUT30), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  AND3_X1   g0533(.A1(new_n460), .A2(new_n593), .A3(new_n595), .ZN(new_n734));
  OAI211_X1 g0534(.A(new_n628), .B(new_n472), .C1(new_n631), .C2(new_n253), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(new_n569), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT30), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n734), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n729), .B1(new_n733), .B2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT96), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n682), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n403), .B1(new_n553), .B2(new_n559), .ZN(new_n742));
  NOR3_X1   g0542(.A1(new_n603), .A2(new_n730), .A3(new_n742), .ZN(new_n743));
  AOI221_X4 g0543(.A(KEYINPUT96), .B1(new_n743), .B2(new_n482), .C1(new_n738), .C2(new_n733), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n727), .B1(new_n741), .B2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n739), .ZN(new_n746));
  INV_X1    g0546(.A(new_n700), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n746), .A2(KEYINPUT31), .A3(new_n747), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n726), .A2(new_n745), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(G330), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n725), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n712), .B1(new_n752), .B2(G1), .ZN(G364));
  NOR2_X1   g0553(.A1(new_n305), .A2(G20), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n205), .B1(new_n754), .B2(G45), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n706), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n695), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n758), .B1(G330), .B2(new_n693), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n227), .B1(G20), .B2(new_n400), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n206), .A2(G179), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n762), .A2(G190), .A3(G200), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(new_n216), .ZN(new_n764));
  NOR2_X1   g0564(.A1(G190), .A2(G200), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(G159), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(KEYINPUT32), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n206), .A2(new_n403), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G200), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(G190), .ZN(new_n772));
  AOI211_X1 g0572(.A(new_n764), .B(new_n769), .C1(G68), .C2(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n770), .A2(new_n765), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n357), .B1(new_n774), .B2(new_n220), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n770), .A2(G190), .A3(new_n335), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n775), .B1(G58), .B2(new_n777), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n762), .A2(new_n337), .A3(G200), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(new_n222), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n780), .B1(new_n768), .B2(KEYINPUT32), .ZN(new_n781));
  NOR3_X1   g0581(.A1(new_n337), .A2(G179), .A3(G200), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(new_n206), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n771), .A2(new_n337), .ZN(new_n785));
  AOI22_X1  g0585(.A1(G97), .A2(new_n784), .B1(new_n785), .B2(G50), .ZN(new_n786));
  NAND4_X1  g0586(.A1(new_n773), .A2(new_n778), .A3(new_n781), .A4(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(G322), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n776), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(G311), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n289), .B1(new_n774), .B2(new_n790), .ZN(new_n791));
  AOI211_X1 g0591(.A(new_n789), .B(new_n791), .C1(G329), .C2(new_n767), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n785), .A2(G326), .ZN(new_n793));
  XNOR2_X1  g0593(.A(KEYINPUT33), .B(G317), .ZN(new_n794));
  INV_X1    g0594(.A(new_n763), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n772), .A2(new_n794), .B1(new_n795), .B2(G303), .ZN(new_n796));
  INV_X1    g0596(.A(new_n779), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n784), .A2(G294), .B1(new_n797), .B2(G283), .ZN(new_n798));
  NAND4_X1  g0598(.A1(new_n792), .A2(new_n793), .A3(new_n796), .A4(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n761), .B1(new_n787), .B2(new_n799), .ZN(new_n800));
  XNOR2_X1  g0600(.A(new_n757), .B(KEYINPUT98), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n209), .A2(new_n357), .ZN(new_n802));
  INV_X1    g0602(.A(G355), .ZN(new_n803));
  OAI22_X1  g0603(.A1(new_n802), .A2(new_n803), .B1(G116), .B2(new_n209), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n705), .A2(new_n261), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n806), .B1(new_n468), .B2(new_n230), .ZN(new_n807));
  OR2_X1    g0607(.A1(new_n243), .A2(new_n468), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n804), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(G13), .A2(G33), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n811), .A2(G20), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n812), .A2(new_n760), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n801), .B1(new_n809), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n800), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n812), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n816), .B1(new_n693), .B2(new_n817), .ZN(new_n818));
  AND2_X1   g0618(.A1(new_n759), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(G396));
  INV_X1    g0620(.A(new_n785), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n821), .A2(new_n547), .B1(new_n763), .B2(new_n222), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n822), .B1(G87), .B2(new_n797), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n357), .B1(new_n777), .B2(G294), .ZN(new_n824));
  INV_X1    g0624(.A(new_n774), .ZN(new_n825));
  AOI22_X1  g0625(.A1(G116), .A2(new_n825), .B1(new_n767), .B2(G311), .ZN(new_n826));
  AOI22_X1  g0626(.A1(G97), .A2(new_n784), .B1(new_n772), .B2(G283), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n823), .A2(new_n824), .A3(new_n826), .A4(new_n827), .ZN(new_n828));
  XOR2_X1   g0628(.A(KEYINPUT99), .B(G143), .Z(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n777), .A2(new_n830), .B1(new_n825), .B2(G159), .ZN(new_n831));
  INV_X1    g0631(.A(new_n772), .ZN(new_n832));
  INV_X1    g0632(.A(G150), .ZN(new_n833));
  INV_X1    g0633(.A(G137), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n831), .B1(new_n832), .B2(new_n833), .C1(new_n834), .C2(new_n821), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT34), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(G58), .ZN(new_n838));
  OAI22_X1  g0638(.A1(new_n783), .A2(new_n838), .B1(new_n779), .B2(new_n214), .ZN(new_n839));
  INV_X1    g0639(.A(G132), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n261), .B1(new_n840), .B2(new_n766), .ZN(new_n841));
  AOI211_X1 g0641(.A(new_n839), .B(new_n841), .C1(G50), .C2(new_n795), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n837), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n835), .A2(new_n836), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n828), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(new_n760), .ZN(new_n846));
  INV_X1    g0646(.A(new_n801), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n760), .A2(new_n810), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n847), .B1(new_n220), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n405), .A2(new_n682), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n407), .B1(new_n384), .B2(new_n689), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n850), .B1(new_n405), .B2(new_n851), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n846), .B(new_n849), .C1(new_n852), .C2(new_n811), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n851), .A2(new_n405), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n854), .B1(new_n405), .B2(new_n682), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n722), .A2(new_n855), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n700), .B(new_n852), .C1(new_n717), .C2(new_n721), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  OR2_X1    g0658(.A1(new_n858), .A2(new_n750), .ZN(new_n859));
  INV_X1    g0659(.A(new_n757), .ZN(new_n860));
  AND2_X1   g0660(.A1(new_n858), .A2(new_n750), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT100), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n859), .B(new_n860), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n861), .A2(new_n862), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n853), .B1(new_n863), .B2(new_n865), .ZN(G384));
  OR2_X1    g0666(.A1(new_n583), .A2(KEYINPUT35), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n583), .A2(KEYINPUT35), .ZN(new_n868));
  NAND4_X1  g0668(.A1(new_n867), .A2(G116), .A3(new_n228), .A4(new_n868), .ZN(new_n869));
  XOR2_X1   g0669(.A(new_n869), .B(KEYINPUT36), .Z(new_n870));
  OAI211_X1 g0670(.A(new_n230), .B(G77), .C1(new_n838), .C2(new_n214), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n344), .A2(G68), .ZN(new_n872));
  AOI211_X1 g0672(.A(new_n205), .B(G13), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n870), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(G169), .B1(new_n431), .B2(new_n435), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(KEYINPUT14), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n876), .A2(new_n439), .A3(new_n436), .ZN(new_n877));
  AND3_X1   g0677(.A1(new_n444), .A2(new_n418), .A3(new_n445), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n419), .B(new_n682), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n418), .A2(new_n689), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n443), .A2(new_n446), .A3(new_n881), .ZN(new_n882));
  AND2_X1   g0682(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  XOR2_X1   g0683(.A(new_n850), .B(KEYINPUT101), .Z(new_n884));
  AOI21_X1  g0684(.A(new_n883), .B1(new_n857), .B2(new_n884), .ZN(new_n885));
  OR2_X1    g0685(.A1(new_n280), .A2(new_n282), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT16), .B1(new_n886), .B2(new_n272), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n321), .B1(new_n887), .B2(new_n286), .ZN(new_n888));
  INV_X1    g0688(.A(new_n680), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n342), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n303), .A2(new_n287), .ZN(new_n893));
  AND2_X1   g0693(.A1(new_n283), .A2(new_n285), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n318), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n269), .ZN(new_n896));
  NOR3_X1   g0696(.A1(new_n895), .A2(KEYINPUT102), .A3(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT102), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n898), .B1(new_n328), .B2(new_n269), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n328), .A2(new_n889), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT37), .ZN(new_n902));
  AND3_X1   g0702(.A1(new_n901), .A2(new_n902), .A3(new_n340), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n888), .A2(new_n269), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n904), .A2(new_n890), .A3(new_n340), .ZN(new_n905));
  AOI22_X1  g0705(.A1(new_n900), .A2(new_n903), .B1(KEYINPUT37), .B2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(KEYINPUT38), .B1(new_n892), .B2(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n890), .B1(new_n334), .B2(new_n341), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT38), .ZN(new_n910));
  NOR3_X1   g0710(.A1(new_n909), .A2(new_n906), .A3(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n885), .B1(new_n908), .B2(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n333), .A2(new_n319), .A3(new_n680), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(KEYINPUT103), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT39), .ZN(new_n916));
  XNOR2_X1  g0716(.A(KEYINPUT104), .B(KEYINPUT38), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT105), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n340), .B(new_n919), .C1(new_n895), .C2(new_n896), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n901), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n919), .B1(new_n331), .B2(new_n340), .ZN(new_n922));
  OAI21_X1  g0722(.A(KEYINPUT37), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n900), .A2(new_n903), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n901), .B1(new_n655), .B2(new_n341), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n918), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n916), .B1(new_n928), .B2(new_n911), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n877), .A2(new_n419), .A3(new_n689), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n892), .A2(new_n907), .A3(KEYINPUT38), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n910), .B1(new_n909), .B2(new_n906), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n932), .A2(KEYINPUT39), .A3(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n929), .A2(new_n931), .A3(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT103), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n912), .A2(new_n936), .A3(new_n913), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n915), .A2(new_n935), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n660), .A2(new_n376), .ZN(new_n939));
  OAI21_X1  g0739(.A(KEYINPUT106), .B1(new_n725), .B2(new_n449), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT106), .ZN(new_n941));
  AOI22_X1  g0741(.A1(new_n713), .A2(KEYINPUT29), .B1(new_n722), .B2(new_n723), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n450), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n939), .B1(new_n940), .B2(new_n943), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n938), .B(new_n944), .ZN(new_n945));
  NOR3_X1   g0745(.A1(new_n741), .A2(new_n744), .A3(new_n727), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n745), .B1(new_n946), .B2(KEYINPUT107), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT107), .ZN(new_n948));
  OAI211_X1 g0748(.A(new_n948), .B(new_n727), .C1(new_n741), .C2(new_n744), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n947), .A2(new_n726), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n855), .B1(new_n882), .B2(new_n879), .ZN(new_n951));
  OAI211_X1 g0751(.A(new_n950), .B(new_n951), .C1(new_n928), .C2(new_n911), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(KEYINPUT40), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n932), .A2(new_n933), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT40), .ZN(new_n955));
  NAND4_X1  g0755(.A1(new_n954), .A2(new_n955), .A3(new_n950), .A4(new_n951), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n953), .A2(new_n956), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n450), .A2(new_n950), .ZN(new_n958));
  AND2_X1   g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n957), .A2(new_n958), .ZN(new_n960));
  INV_X1    g0760(.A(G330), .ZN(new_n961));
  NOR3_X1   g0761(.A1(new_n959), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  OAI22_X1  g0762(.A1(new_n945), .A2(new_n962), .B1(new_n205), .B2(new_n754), .ZN(new_n963));
  AND2_X1   g0763(.A1(new_n945), .A2(new_n962), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n874), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n965), .B(KEYINPUT108), .Z(G367));
  AOI21_X1  g0766(.A(new_n689), .B1(new_n636), .B2(new_n645), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n967), .B(KEYINPUT109), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n968), .A2(new_n670), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n969), .B1(new_n668), .B2(new_n968), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT43), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(new_n698), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n666), .B1(new_n586), .B2(new_n700), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n665), .A2(new_n747), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n973), .A2(new_n976), .ZN(new_n977));
  OR2_X1    g0777(.A1(new_n977), .A2(KEYINPUT42), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n605), .B1(new_n974), .B2(new_n530), .ZN(new_n979));
  AOI22_X1  g0779(.A1(new_n977), .A2(KEYINPUT42), .B1(new_n700), .B2(new_n979), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n972), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n970), .A2(new_n971), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND4_X1  g0783(.A1(new_n978), .A2(new_n980), .A3(new_n971), .A4(new_n970), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n976), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n696), .A2(new_n986), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n985), .B(new_n987), .Z(new_n988));
  XNOR2_X1  g0788(.A(KEYINPUT110), .B(KEYINPUT41), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n706), .B(new_n989), .Z(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n976), .B1(new_n702), .B2(new_n703), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT45), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  OAI211_X1 g0794(.A(KEYINPUT45), .B(new_n976), .C1(new_n702), .C2(new_n703), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n698), .A2(new_n701), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(KEYINPUT94), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n698), .A2(new_n699), .A3(new_n701), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n998), .A2(new_n999), .A3(new_n986), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT44), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND4_X1  g0802(.A1(new_n998), .A2(KEYINPUT44), .A3(new_n999), .A4(new_n986), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  AND3_X1   g0804(.A1(new_n996), .A2(new_n1004), .A3(new_n696), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n696), .B1(new_n996), .B2(new_n1004), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n690), .A2(new_n697), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n695), .B1(new_n1007), .B2(new_n973), .ZN(new_n1008));
  OAI211_X1 g0808(.A(new_n694), .B(new_n698), .C1(new_n690), .C2(new_n697), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n751), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  NOR3_X1   g0811(.A1(new_n1005), .A2(new_n1006), .A3(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n991), .B1(new_n1012), .B2(new_n751), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n988), .B1(new_n1013), .B2(new_n755), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n970), .A2(new_n812), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n805), .A2(new_n239), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n1016), .B(new_n813), .C1(new_n209), .C2(new_n379), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n801), .A2(new_n1017), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n1018), .B(KEYINPUT111), .Z(new_n1019));
  INV_X1    g0819(.A(G159), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n832), .A2(new_n1020), .B1(new_n779), .B2(new_n220), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1021), .B1(G58), .B2(new_n795), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n776), .A2(new_n833), .B1(new_n766), .B2(new_n834), .ZN(new_n1023));
  AOI211_X1 g0823(.A(new_n289), .B(new_n1023), .C1(G50), .C2(new_n825), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n785), .A2(new_n830), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n784), .A2(G68), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n1022), .A2(new_n1024), .A3(new_n1025), .A4(new_n1026), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(G283), .A2(new_n825), .B1(new_n767), .B2(G317), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n551), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1028), .B1(new_n1029), .B2(new_n776), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n1030), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n783), .A2(new_n391), .B1(new_n779), .B2(new_n536), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1032), .B1(G294), .B2(new_n772), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT46), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(new_n763), .B2(new_n540), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n261), .B1(new_n785), .B2(G311), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1031), .A2(new_n1033), .A3(new_n1035), .A4(new_n1036), .ZN(new_n1037));
  NOR3_X1   g0837(.A1(new_n763), .A2(new_n1034), .A3(new_n540), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT112), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1027), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT47), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n760), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n1015), .B(new_n1019), .C1(new_n1042), .C2(new_n1044), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT113), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n1014), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n1047), .ZN(G387));
  NAND3_X1  g0848(.A1(new_n1011), .A2(KEYINPUT116), .A3(new_n706), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT116), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n706), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1050), .B1(new_n1010), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1049), .B(new_n1052), .C1(new_n752), .C2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1053), .A2(new_n756), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n806), .B1(new_n236), .B2(G45), .ZN(new_n1056));
  AOI211_X1 g0856(.A(G45), .B(new_n708), .C1(G68), .C2(G77), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n1057), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1058), .A2(KEYINPUT114), .ZN(new_n1059));
  OAI21_X1  g0859(.A(KEYINPUT50), .B1(new_n309), .B2(G50), .ZN(new_n1060));
  OR3_X1    g0860(.A1(new_n309), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT114), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n1060), .B(new_n1061), .C1(new_n1057), .C2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1056), .B1(new_n1059), .B2(new_n1063), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n1064), .B1(G107), .B2(new_n209), .C1(new_n707), .C2(new_n802), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n847), .B1(new_n1065), .B2(new_n813), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n821), .A2(new_n1020), .B1(new_n763), .B2(new_n220), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n776), .A2(new_n344), .B1(new_n766), .B2(new_n833), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(G68), .B2(new_n825), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n618), .A2(new_n784), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n598), .B1(G97), .B2(new_n797), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1069), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  AOI211_X1 g0872(.A(new_n1067), .B(new_n1072), .C1(new_n310), .C2(new_n772), .ZN(new_n1073));
  INV_X1    g0873(.A(G283), .ZN(new_n1074));
  INV_X1    g0874(.A(G294), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n783), .A2(new_n1074), .B1(new_n763), .B2(new_n1075), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n777), .A2(G317), .B1(new_n825), .B2(new_n551), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n1077), .B1(new_n832), .B2(new_n790), .C1(new_n788), .C2(new_n821), .ZN(new_n1078));
  INV_X1    g0878(.A(KEYINPUT48), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1076), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1080), .B1(new_n1079), .B2(new_n1078), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1081), .B(KEYINPUT49), .ZN(new_n1082));
  OR2_X1    g0882(.A1(new_n1082), .A2(KEYINPUT115), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n261), .B1(G326), .B2(new_n767), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1084), .B1(new_n540), .B2(new_n779), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1085), .B1(new_n1082), .B2(KEYINPUT115), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1073), .B1(new_n1083), .B2(new_n1086), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n1066), .B1(new_n761), .B2(new_n1087), .C1(new_n690), .C2(new_n817), .ZN(new_n1088));
  AND2_X1   g0888(.A1(new_n1055), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1054), .A2(new_n1089), .ZN(G393));
  OAI21_X1  g0890(.A(new_n1011), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n996), .A2(new_n1004), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n696), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n996), .A2(new_n1004), .A3(new_n696), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1094), .A2(new_n1095), .A3(new_n1010), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1091), .A2(new_n1096), .A3(new_n706), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n986), .A2(new_n812), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n813), .B1(new_n536), .B2(new_n209), .C1(new_n806), .C2(new_n246), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n801), .A2(new_n1100), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n821), .A2(new_n833), .B1(new_n1020), .B2(new_n776), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT51), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n767), .A2(new_n830), .B1(new_n825), .B2(new_n310), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n832), .A2(new_n344), .B1(new_n220), .B2(new_n783), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n214), .A2(new_n763), .B1(new_n779), .B2(new_n216), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n1103), .A2(new_n261), .A3(new_n1104), .A4(new_n1107), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(G317), .A2(new_n785), .B1(new_n777), .B2(G311), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(new_n1109), .B(KEYINPUT117), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1110), .B(KEYINPUT52), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n783), .A2(new_n540), .B1(new_n774), .B2(new_n1075), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1112), .B1(new_n551), .B2(new_n772), .ZN(new_n1113));
  XOR2_X1   g0913(.A(new_n1113), .B(KEYINPUT118), .Z(new_n1114));
  OAI21_X1  g0914(.A(new_n289), .B1(new_n766), .B2(new_n788), .ZN(new_n1115));
  AOI211_X1 g0915(.A(new_n780), .B(new_n1115), .C1(G283), .C2(new_n795), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1108), .B1(new_n1111), .B2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1101), .B1(new_n1118), .B2(new_n760), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n1098), .A2(new_n756), .B1(new_n1099), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1097), .A2(new_n1120), .ZN(G390));
  AOI21_X1  g0921(.A(new_n850), .B1(new_n713), .B2(new_n854), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n930), .B1(new_n1122), .B2(new_n883), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n928), .A2(new_n911), .ZN(new_n1124));
  OR2_X1    g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n929), .A2(new_n934), .ZN(new_n1126));
  OR2_X1    g0926(.A1(new_n885), .A2(new_n931), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n749), .A2(new_n951), .A3(G330), .ZN(new_n1129));
  AND2_X1   g0929(.A1(new_n950), .A2(G330), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1129), .B1(new_n1130), .B2(KEYINPUT119), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1125), .A2(new_n1128), .A3(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n950), .A2(G330), .A3(new_n951), .ZN(new_n1133));
  OR2_X1    g0933(.A1(new_n1133), .A2(KEYINPUT119), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n885), .A2(new_n931), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1135), .B1(new_n929), .B2(new_n934), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1134), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1132), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n811), .B1(new_n929), .B2(new_n934), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n848), .A2(new_n309), .ZN(new_n1142));
  INV_X1    g0942(.A(G125), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n776), .A2(new_n840), .B1(new_n766), .B2(new_n1143), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(KEYINPUT54), .B(G143), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1145), .ZN(new_n1146));
  AOI211_X1 g0946(.A(new_n289), .B(new_n1144), .C1(new_n825), .C2(new_n1146), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n763), .A2(new_n833), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(KEYINPUT121), .B(KEYINPUT53), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n1148), .B(new_n1149), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n785), .A2(G128), .B1(new_n797), .B2(G50), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(G159), .A2(new_n784), .B1(new_n772), .B2(G137), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n1147), .A2(new_n1150), .A3(new_n1151), .A4(new_n1152), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n776), .A2(new_n540), .B1(new_n766), .B2(new_n1075), .ZN(new_n1154));
  AOI211_X1 g0954(.A(new_n357), .B(new_n1154), .C1(G97), .C2(new_n825), .ZN(new_n1155));
  OR2_X1    g0955(.A1(new_n832), .A2(new_n391), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(G77), .A2(new_n784), .B1(new_n785), .B2(G283), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n764), .B1(G68), .B2(new_n797), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1155), .A2(new_n1156), .A3(new_n1157), .A4(new_n1158), .ZN(new_n1159));
  AND2_X1   g0959(.A1(new_n1153), .A2(new_n1159), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n801), .B(new_n1142), .C1(new_n1160), .C2(new_n761), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n1140), .A2(new_n755), .B1(new_n1141), .B2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n883), .B1(new_n750), .B2(new_n855), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n1163), .A2(new_n1133), .B1(new_n857), .B2(new_n884), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n950), .A2(G330), .A3(new_n852), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(new_n883), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT120), .ZN(new_n1168));
  AND2_X1   g0968(.A1(new_n1129), .A2(new_n1122), .ZN(new_n1169));
  AND3_X1   g0969(.A1(new_n1167), .A2(new_n1168), .A3(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1168), .B1(new_n1167), .B2(new_n1169), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1165), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1130), .A2(new_n450), .ZN(new_n1173));
  NOR3_X1   g0973(.A1(new_n725), .A2(KEYINPUT106), .A3(new_n449), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n941), .B1(new_n450), .B2(new_n942), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n661), .B(new_n1173), .C1(new_n1174), .C2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1139), .A2(new_n1172), .A3(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1172), .A2(new_n1177), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1051), .B1(new_n1140), .B2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1162), .B1(new_n1178), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(G378));
  INV_X1    g0982(.A(KEYINPUT123), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n377), .A2(new_n354), .A3(new_n889), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n354), .A2(new_n889), .ZN(new_n1185));
  NAND4_X1  g0985(.A1(new_n371), .A2(new_n376), .A3(new_n373), .A4(new_n1185), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1187));
  AND3_X1   g0987(.A1(new_n1184), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1187), .B1(new_n1184), .B2(new_n1186), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1190), .A2(new_n810), .ZN(new_n1191));
  OAI221_X1 g0991(.A(new_n1026), .B1(new_n1074), .B2(new_n766), .C1(new_n222), .C2(new_n776), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(new_n618), .B2(new_n825), .ZN(new_n1193));
  INV_X1    g0993(.A(G41), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1193), .A2(new_n1194), .A3(new_n598), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n763), .A2(new_n220), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n779), .A2(new_n838), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n832), .A2(new_n536), .B1(new_n821), .B2(new_n540), .ZN(new_n1198));
  NOR4_X1   g0998(.A1(new_n1195), .A2(new_n1196), .A3(new_n1197), .A4(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1199), .A2(KEYINPUT58), .ZN(new_n1200));
  AOI21_X1  g1000(.A(G50), .B1(new_n257), .B2(new_n1194), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1201), .B1(new_n261), .B2(G41), .ZN(new_n1202));
  AND2_X1   g1002(.A1(new_n1200), .A2(new_n1202), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n832), .A2(new_n840), .B1(new_n821), .B2(new_n1143), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n777), .A2(G128), .B1(new_n825), .B2(G137), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1205), .B1(new_n763), .B2(new_n1145), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n1204), .B(new_n1206), .C1(G150), .C2(new_n784), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1208), .A2(KEYINPUT59), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1208), .A2(KEYINPUT59), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n797), .A2(G159), .ZN(new_n1211));
  AOI211_X1 g1011(.A(G33), .B(G41), .C1(new_n767), .C2(G124), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1210), .A2(new_n1211), .A3(new_n1212), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n1203), .B1(KEYINPUT58), .B2(new_n1199), .C1(new_n1209), .C2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1214), .A2(new_n760), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n860), .B1(new_n344), .B2(new_n848), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1191), .A2(new_n1215), .A3(new_n1216), .ZN(new_n1217));
  AND2_X1   g1017(.A1(new_n950), .A2(new_n951), .ZN(new_n1218));
  AOI21_X1  g1018(.A(KEYINPUT40), .B1(new_n932), .B2(new_n933), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(KEYINPUT40), .A2(new_n952), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1190), .B1(new_n1220), .B2(new_n961), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1190), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n957), .A2(G330), .A3(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT122), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n1221), .A2(new_n1223), .B1(new_n938), .B2(new_n1224), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n915), .A2(KEYINPUT122), .A3(new_n935), .A4(new_n937), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1222), .B1(new_n957), .B2(G330), .ZN(new_n1227));
  AOI211_X1 g1027(.A(new_n961), .B(new_n1190), .C1(new_n953), .C2(new_n956), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n937), .A2(new_n935), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n936), .B1(new_n912), .B2(new_n913), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n1225), .A2(new_n1226), .B1(new_n1229), .B2(new_n1232), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1183), .B(new_n1217), .C1(new_n1233), .C2(new_n755), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1224), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n1235), .B(new_n1226), .C1(new_n1227), .C2(new_n1228), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1221), .A2(new_n1232), .A3(new_n1223), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n755), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1217), .ZN(new_n1239));
  OAI21_X1  g1039(.A(KEYINPUT123), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1234), .A2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT57), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1176), .A2(KEYINPUT124), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT124), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n944), .A2(new_n1244), .A3(new_n1173), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1243), .A2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(KEYINPUT120), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1167), .A2(new_n1168), .A3(new_n1169), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1176), .B1(new_n1250), .B2(new_n1165), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1246), .B1(new_n1251), .B2(new_n1139), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1242), .B1(new_n1233), .B2(new_n1252), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n938), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1242), .B1(new_n1254), .B2(new_n1237), .ZN(new_n1255));
  AND2_X1   g1055(.A1(new_n1243), .A2(new_n1245), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1178), .A2(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1051), .B1(new_n1255), .B2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1253), .A2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1241), .A2(new_n1259), .ZN(G375));
  OAI211_X1 g1060(.A(new_n1176), .B(new_n1165), .C1(new_n1170), .C2(new_n1171), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1179), .A2(new_n991), .A3(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n883), .A2(new_n810), .ZN(new_n1263));
  NOR3_X1   g1063(.A1(new_n760), .A2(G68), .A3(new_n810), .ZN(new_n1264));
  OAI22_X1  g1064(.A1(new_n776), .A2(new_n834), .B1(new_n774), .B2(new_n833), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1265), .B1(G128), .B2(new_n767), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(G50), .A2(new_n784), .B1(new_n785), .B2(G132), .ZN(new_n1267));
  AOI22_X1  g1067(.A1(new_n772), .A2(new_n1146), .B1(new_n795), .B2(G159), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1197), .A2(new_n598), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1266), .A2(new_n1267), .A3(new_n1268), .A4(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n772), .A2(G116), .ZN(new_n1271));
  OAI221_X1 g1071(.A(new_n1271), .B1(new_n391), .B2(new_n774), .C1(new_n821), .C2(new_n1075), .ZN(new_n1272));
  XOR2_X1   g1072(.A(new_n1272), .B(KEYINPUT125), .Z(new_n1273));
  OAI21_X1  g1073(.A(new_n289), .B1(new_n766), .B2(new_n547), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1274), .B1(G283), .B2(new_n777), .ZN(new_n1275));
  AOI22_X1  g1075(.A1(new_n795), .A2(G97), .B1(new_n797), .B2(G77), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1070), .A2(new_n1275), .A3(new_n1276), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1270), .B1(new_n1273), .B2(new_n1277), .ZN(new_n1278));
  AOI211_X1 g1078(.A(new_n847), .B(new_n1264), .C1(new_n1278), .C2(new_n760), .ZN(new_n1279));
  AOI22_X1  g1079(.A1(new_n1172), .A2(new_n756), .B1(new_n1263), .B2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1262), .A2(new_n1280), .ZN(G381));
  NOR2_X1   g1081(.A1(G375), .A2(G378), .ZN(new_n1282));
  INV_X1    g1082(.A(G390), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1054), .A2(new_n819), .A3(new_n1089), .ZN(new_n1284));
  NOR3_X1   g1084(.A1(new_n1284), .A2(G384), .A3(G381), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1282), .A2(new_n1047), .A3(new_n1283), .A4(new_n1285), .ZN(G407));
  AOI22_X1  g1086(.A1(new_n1234), .A2(new_n1240), .B1(new_n1253), .B2(new_n1258), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(new_n1181), .ZN(new_n1288));
  OAI211_X1 g1088(.A(G407), .B(G213), .C1(G343), .C2(new_n1288), .ZN(G409));
  NAND3_X1  g1089(.A1(new_n681), .A2(G213), .A3(G2897), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT60), .ZN(new_n1292));
  OAI21_X1  g1092(.A(KEYINPUT127), .B1(new_n1261), .B2(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1164), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT127), .ZN(new_n1295));
  NAND4_X1  g1095(.A1(new_n1294), .A2(new_n1295), .A3(KEYINPUT60), .A4(new_n1176), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1051), .B1(new_n1172), .B2(new_n1177), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1261), .A2(new_n1292), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1293), .A2(new_n1296), .A3(new_n1297), .A4(new_n1298), .ZN(new_n1299));
  AND3_X1   g1099(.A1(new_n1299), .A2(G384), .A3(new_n1280), .ZN(new_n1300));
  AOI21_X1  g1100(.A(G384), .B1(new_n1299), .B2(new_n1280), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1291), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1299), .A2(new_n1280), .ZN(new_n1303));
  INV_X1    g1103(.A(G384), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1299), .A2(G384), .A3(new_n1280), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1305), .A2(new_n1306), .A3(new_n1290), .ZN(new_n1307));
  AND2_X1   g1107(.A1(new_n1302), .A2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n681), .A2(G213), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1257), .A2(new_n1310), .A3(new_n991), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT126), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1257), .A2(new_n1310), .A3(KEYINPUT126), .A4(new_n991), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1254), .A2(new_n1237), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1239), .B1(new_n1315), .B2(new_n756), .ZN(new_n1316));
  NAND4_X1  g1116(.A1(new_n1313), .A2(new_n1181), .A3(new_n1314), .A4(new_n1316), .ZN(new_n1317));
  OAI211_X1 g1117(.A(new_n1309), .B(new_n1317), .C1(new_n1287), .C2(new_n1181), .ZN(new_n1318));
  AOI21_X1  g1118(.A(KEYINPUT61), .B1(new_n1308), .B2(new_n1318), .ZN(new_n1319));
  NOR2_X1   g1119(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1320), .ZN(new_n1321));
  OAI21_X1  g1121(.A(KEYINPUT62), .B1(new_n1318), .B2(new_n1321), .ZN(new_n1322));
  AND2_X1   g1122(.A1(new_n1317), .A2(new_n1309), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(G375), .A2(G378), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT62), .ZN(new_n1325));
  NAND4_X1  g1125(.A1(new_n1323), .A2(new_n1324), .A3(new_n1325), .A4(new_n1320), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1319), .A2(new_n1322), .A3(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(G393), .A2(G396), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1328), .A2(new_n1284), .ZN(new_n1329));
  XNOR2_X1  g1129(.A(new_n985), .B(new_n987), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n990), .B1(new_n1096), .B2(new_n752), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n1330), .B1(new_n1331), .B2(new_n756), .ZN(new_n1332));
  INV_X1    g1132(.A(new_n1046), .ZN(new_n1333));
  AND3_X1   g1133(.A1(new_n1332), .A2(new_n1333), .A3(G390), .ZN(new_n1334));
  AOI21_X1  g1134(.A(G390), .B1(new_n1332), .B2(new_n1333), .ZN(new_n1335));
  OAI21_X1  g1135(.A(new_n1329), .B1(new_n1334), .B2(new_n1335), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1283), .B1(new_n1014), .B2(new_n1046), .ZN(new_n1337));
  INV_X1    g1137(.A(new_n1329), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1332), .A2(new_n1333), .A3(G390), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1337), .A2(new_n1338), .A3(new_n1339), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1336), .A2(new_n1340), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1327), .A2(new_n1341), .ZN(new_n1342));
  NOR3_X1   g1142(.A1(new_n1334), .A2(new_n1335), .A3(new_n1329), .ZN(new_n1343));
  AOI21_X1  g1143(.A(new_n1338), .B1(new_n1337), .B2(new_n1339), .ZN(new_n1344));
  NOR2_X1   g1144(.A1(new_n1343), .A2(new_n1344), .ZN(new_n1345));
  NAND4_X1  g1145(.A1(new_n1323), .A2(new_n1324), .A3(KEYINPUT63), .A4(new_n1320), .ZN(new_n1346));
  INV_X1    g1146(.A(KEYINPUT63), .ZN(new_n1347));
  OAI21_X1  g1147(.A(new_n1347), .B1(new_n1318), .B2(new_n1321), .ZN(new_n1348));
  NAND4_X1  g1148(.A1(new_n1345), .A2(new_n1319), .A3(new_n1346), .A4(new_n1348), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1342), .A2(new_n1349), .ZN(G405));
  NAND2_X1  g1150(.A1(new_n1324), .A2(new_n1288), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1351), .A2(new_n1320), .ZN(new_n1352));
  NAND3_X1  g1152(.A1(new_n1324), .A2(new_n1288), .A3(new_n1321), .ZN(new_n1353));
  AND4_X1   g1153(.A1(new_n1340), .A2(new_n1352), .A3(new_n1336), .A4(new_n1353), .ZN(new_n1354));
  AOI22_X1  g1154(.A1(new_n1352), .A2(new_n1353), .B1(new_n1336), .B2(new_n1340), .ZN(new_n1355));
  NOR2_X1   g1155(.A1(new_n1354), .A2(new_n1355), .ZN(G402));
endmodule


