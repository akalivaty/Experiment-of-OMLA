

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781;

  NOR2_X1 U375 ( .A1(G953), .A2(G237), .ZN(n509) );
  AND2_X2 U376 ( .A1(n666), .A2(n654), .ZN(n359) );
  AND2_X2 U377 ( .A1(n655), .A2(n654), .ZN(n360) );
  AND2_X2 U378 ( .A1(n413), .A2(n412), .ZN(n411) );
  AND2_X1 U379 ( .A1(n771), .A2(n433), .ZN(n432) );
  INV_X1 U380 ( .A(G953), .ZN(n477) );
  BUF_X1 U381 ( .A(n477), .Z(n772) );
  AND2_X2 U382 ( .A1(n672), .A2(n654), .ZN(n353) );
  NOR2_X2 U383 ( .A1(n781), .A2(n780), .ZN(n373) );
  XNOR2_X2 U384 ( .A(n619), .B(n618), .ZN(n781) );
  XNOR2_X2 U385 ( .A(n560), .B(n466), .ZN(n610) );
  OR2_X1 U386 ( .A1(n556), .A2(n555), .ZN(n686) );
  NAND2_X1 U387 ( .A1(n553), .A2(n540), .ZN(n541) );
  AND2_X1 U388 ( .A1(n544), .A2(n605), .ZN(n553) );
  AND2_X1 U389 ( .A1(n611), .A2(n389), .ZN(n709) );
  XNOR2_X1 U390 ( .A(n539), .B(n538), .ZN(n544) );
  NOR2_X1 U391 ( .A1(n713), .A2(n718), .ZN(n540) );
  XNOR2_X1 U392 ( .A(n369), .B(n517), .ZN(n594) );
  OR2_X1 U393 ( .A1(n669), .A2(n426), .ZN(n425) );
  XNOR2_X1 U394 ( .A(n680), .B(n679), .ZN(n681) );
  XNOR2_X1 U395 ( .A(n490), .B(n755), .ZN(n669) );
  XNOR2_X1 U396 ( .A(n484), .B(n458), .ZN(n767) );
  XNOR2_X1 U397 ( .A(n518), .B(KEYINPUT4), .ZN(n484) );
  XNOR2_X1 U398 ( .A(n388), .B(KEYINPUT80), .ZN(n479) );
  XNOR2_X1 U399 ( .A(n423), .B(G104), .ZN(n487) );
  NAND2_X1 U400 ( .A1(n477), .A2(G224), .ZN(n388) );
  XNOR2_X1 U401 ( .A(KEYINPUT3), .B(G119), .ZN(n471) );
  XNOR2_X1 U402 ( .A(G101), .B(KEYINPUT74), .ZN(n469) );
  XNOR2_X1 U403 ( .A(G110), .B(G107), .ZN(n423) );
  XNOR2_X1 U404 ( .A(G146), .B(G125), .ZN(n478) );
  XNOR2_X2 U405 ( .A(n643), .B(KEYINPUT65), .ZN(n354) );
  XNOR2_X1 U406 ( .A(n643), .B(KEYINPUT65), .ZN(n675) );
  NAND2_X2 U407 ( .A1(n642), .A2(n641), .ZN(n643) );
  OR2_X1 U408 ( .A1(n669), .A2(n381), .ZN(n380) );
  NAND2_X1 U409 ( .A1(n600), .A2(n599), .ZN(n397) );
  XNOR2_X1 U410 ( .A(n478), .B(n437), .ZN(n513) );
  INV_X1 U411 ( .A(n709), .ZN(n405) );
  NAND2_X1 U412 ( .A1(n378), .A2(n377), .ZN(n585) );
  INV_X1 U413 ( .A(n705), .ZN(n377) );
  INV_X1 U414 ( .A(n703), .ZN(n378) );
  INV_X1 U415 ( .A(n620), .ZN(n729) );
  OR2_X1 U416 ( .A1(n676), .A2(G902), .ZN(n465) );
  XNOR2_X1 U417 ( .A(n441), .B(n403), .ZN(n522) );
  INV_X1 U418 ( .A(KEYINPUT8), .ZN(n403) );
  XNOR2_X1 U419 ( .A(n438), .B(KEYINPUT70), .ZN(n459) );
  NAND2_X1 U420 ( .A1(n415), .A2(n355), .ZN(n414) );
  NAND2_X1 U421 ( .A1(n424), .A2(n364), .ZN(n606) );
  NAND2_X1 U422 ( .A1(n383), .A2(n382), .ZN(n424) );
  BUF_X1 U423 ( .A(n560), .Z(n581) );
  NAND2_X1 U424 ( .A1(G472), .A2(G902), .ZN(n412) );
  XNOR2_X1 U425 ( .A(n459), .B(n513), .ZN(n769) );
  XNOR2_X1 U426 ( .A(G119), .B(G110), .ZN(n442) );
  XNOR2_X1 U427 ( .A(G143), .B(G104), .ZN(n510) );
  XOR2_X1 U428 ( .A(G140), .B(G122), .Z(n511) );
  XNOR2_X1 U429 ( .A(n385), .B(n506), .ZN(n508) );
  XOR2_X1 U430 ( .A(KEYINPUT95), .B(KEYINPUT11), .Z(n506) );
  XNOR2_X1 U431 ( .A(n505), .B(n386), .ZN(n385) );
  INV_X1 U432 ( .A(KEYINPUT12), .ZN(n386) );
  AND2_X2 U433 ( .A1(n421), .A2(n629), .ZN(n771) );
  XNOR2_X1 U434 ( .A(n371), .B(n623), .ZN(n421) );
  XNOR2_X1 U435 ( .A(n606), .B(n494), .ZN(n583) );
  XNOR2_X1 U436 ( .A(KEYINPUT67), .B(KEYINPUT19), .ZN(n494) );
  XNOR2_X1 U437 ( .A(n447), .B(n357), .ZN(n448) );
  NAND2_X1 U438 ( .A1(n652), .A2(n527), .ZN(n369) );
  AND2_X1 U439 ( .A1(n394), .A2(n407), .ZN(n393) );
  AND2_X1 U440 ( .A1(n398), .A2(n396), .ZN(n395) );
  INV_X1 U441 ( .A(KEYINPUT87), .ZN(n381) );
  OR2_X1 U442 ( .A1(n492), .A2(n381), .ZN(n379) );
  XNOR2_X1 U443 ( .A(G116), .B(G113), .ZN(n470) );
  XNOR2_X1 U444 ( .A(n585), .B(n567), .ZN(n588) );
  XOR2_X1 U445 ( .A(G122), .B(G107), .Z(n520) );
  INV_X1 U446 ( .A(G128), .ZN(n456) );
  XNOR2_X1 U447 ( .A(KEYINPUT18), .B(KEYINPUT90), .ZN(n480) );
  XNOR2_X1 U448 ( .A(KEYINPUT81), .B(KEYINPUT17), .ZN(n481) );
  XNOR2_X1 U449 ( .A(n375), .B(n404), .ZN(n374) );
  XNOR2_X1 U450 ( .A(n373), .B(KEYINPUT46), .ZN(n372) );
  INV_X1 U451 ( .A(KEYINPUT72), .ZN(n404) );
  AND2_X1 U452 ( .A1(n660), .A2(n545), .ZN(n546) );
  AND2_X1 U453 ( .A1(n674), .A2(n549), .ZN(n550) );
  XNOR2_X1 U454 ( .A(n596), .B(n612), .ZN(n620) );
  NAND2_X1 U455 ( .A1(n631), .A2(n492), .ZN(n429) );
  NAND2_X1 U456 ( .A1(n428), .A2(n427), .ZN(n426) );
  INV_X1 U457 ( .A(n631), .ZN(n427) );
  INV_X1 U458 ( .A(n492), .ZN(n428) );
  XNOR2_X1 U459 ( .A(KEYINPUT16), .B(G122), .ZN(n486) );
  XNOR2_X1 U460 ( .A(n390), .B(KEYINPUT41), .ZN(n748) );
  NOR2_X1 U461 ( .A1(n733), .A2(n732), .ZN(n390) );
  NOR2_X1 U462 ( .A1(n605), .A2(n604), .ZN(n624) );
  AND2_X1 U463 ( .A1(n703), .A2(n601), .ZN(n602) );
  BUF_X1 U464 ( .A(n610), .Z(n389) );
  NAND2_X1 U465 ( .A1(n410), .A2(n527), .ZN(n409) );
  XNOR2_X1 U466 ( .A(n401), .B(n358), .ZN(n400) );
  XNOR2_X1 U467 ( .A(n370), .B(n516), .ZN(n652) );
  NOR2_X2 U468 ( .A1(n621), .A2(n584), .ZN(n701) );
  AND2_X1 U469 ( .A1(n566), .A2(n565), .ZN(n705) );
  XNOR2_X1 U470 ( .A(n700), .B(n376), .ZN(G45) );
  INV_X1 U471 ( .A(G143), .ZN(n376) );
  AND2_X1 U472 ( .A1(n610), .A2(n362), .ZN(n355) );
  AND2_X1 U473 ( .A1(n380), .A2(n365), .ZN(n356) );
  XNOR2_X1 U474 ( .A(n528), .B(G478), .ZN(n565) );
  XNOR2_X1 U475 ( .A(KEYINPUT25), .B(KEYINPUT93), .ZN(n357) );
  XOR2_X1 U476 ( .A(n440), .B(n439), .Z(n358) );
  AND2_X1 U477 ( .A1(n429), .A2(n728), .ZN(n361) );
  AND2_X1 U478 ( .A1(n561), .A2(n420), .ZN(n362) );
  AND2_X1 U479 ( .A1(n425), .A2(n429), .ZN(n363) );
  OR2_X1 U480 ( .A1(n430), .A2(KEYINPUT87), .ZN(n364) );
  AND2_X1 U481 ( .A1(n361), .A2(n379), .ZN(n365) );
  XOR2_X1 U482 ( .A(n652), .B(n651), .Z(n366) );
  XOR2_X1 U483 ( .A(n669), .B(n670), .Z(n367) );
  AND2_X1 U484 ( .A1(n631), .A2(n630), .ZN(n368) );
  NOR2_X1 U485 ( .A1(n772), .A2(G952), .ZN(n683) );
  XNOR2_X1 U486 ( .A(n514), .B(n515), .ZN(n370) );
  NAND2_X1 U487 ( .A1(n374), .A2(n372), .ZN(n371) );
  NAND2_X1 U488 ( .A1(n406), .A2(n405), .ZN(n375) );
  INV_X1 U489 ( .A(n585), .ZN(n734) );
  NAND2_X1 U490 ( .A1(n669), .A2(n492), .ZN(n430) );
  NAND2_X1 U491 ( .A1(n425), .A2(n361), .ZN(n384) );
  NAND2_X1 U492 ( .A1(n356), .A2(n425), .ZN(n383) );
  NAND2_X1 U493 ( .A1(n384), .A2(KEYINPUT87), .ZN(n382) );
  NAND2_X1 U494 ( .A1(n586), .A2(KEYINPUT47), .ZN(n394) );
  NAND2_X1 U495 ( .A1(n615), .A2(n614), .ZN(n616) );
  NOR2_X2 U496 ( .A1(n591), .A2(n592), .ZN(n615) );
  NAND2_X1 U497 ( .A1(n578), .A2(n562), .ZN(n580) );
  AND2_X2 U498 ( .A1(n387), .A2(n552), .ZN(n573) );
  NAND2_X1 U499 ( .A1(n546), .A2(n547), .ZN(n387) );
  INV_X1 U500 ( .A(n394), .ZN(n399) );
  NAND2_X1 U501 ( .A1(n395), .A2(n391), .ZN(n406) );
  NAND2_X1 U502 ( .A1(n393), .A2(n392), .ZN(n391) );
  INV_X1 U503 ( .A(n397), .ZN(n392) );
  NAND2_X1 U504 ( .A1(n397), .A2(KEYINPUT77), .ZN(n396) );
  NAND2_X1 U505 ( .A1(n399), .A2(KEYINPUT77), .ZN(n398) );
  NAND2_X1 U506 ( .A1(n522), .A2(G221), .ZN(n401) );
  XNOR2_X1 U507 ( .A(n769), .B(n445), .ZN(n402) );
  XNOR2_X1 U508 ( .A(n402), .B(n400), .ZN(n658) );
  INV_X1 U509 ( .A(KEYINPUT77), .ZN(n407) );
  NAND2_X4 U510 ( .A1(n411), .A2(n408), .ZN(n562) );
  OR2_X1 U511 ( .A1(n662), .A2(n409), .ZN(n408) );
  INV_X1 U512 ( .A(G472), .ZN(n410) );
  NAND2_X1 U513 ( .A1(n662), .A2(G472), .ZN(n413) );
  INV_X1 U514 ( .A(n562), .ZN(n557) );
  NAND2_X2 U515 ( .A1(n573), .A2(n572), .ZN(n422) );
  NOR2_X1 U516 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X2 U517 ( .A(n617), .B(n616), .ZN(n628) );
  OR2_X2 U518 ( .A1(n674), .A2(KEYINPUT68), .ZN(n534) );
  NAND2_X1 U519 ( .A1(n674), .A2(n434), .ZN(n535) );
  XNOR2_X2 U520 ( .A(n532), .B(n531), .ZN(n674) );
  NAND2_X1 U521 ( .A1(n610), .A2(n561), .ZN(n418) );
  NAND2_X1 U522 ( .A1(n416), .A2(n414), .ZN(n737) );
  INV_X1 U523 ( .A(n605), .ZN(n415) );
  AND2_X1 U524 ( .A1(n417), .A2(n419), .ZN(n416) );
  NAND2_X1 U525 ( .A1(n418), .A2(n476), .ZN(n417) );
  NAND2_X1 U526 ( .A1(n605), .A2(n476), .ZN(n419) );
  INV_X1 U527 ( .A(n476), .ZN(n420) );
  XNOR2_X2 U528 ( .A(n562), .B(KEYINPUT6), .ZN(n605) );
  NAND2_X1 U529 ( .A1(n759), .A2(n771), .ZN(n712) );
  XNOR2_X2 U530 ( .A(n422), .B(KEYINPUT45), .ZN(n759) );
  NAND2_X1 U531 ( .A1(n363), .A2(n430), .ZN(n596) );
  NAND2_X1 U532 ( .A1(n431), .A2(n368), .ZN(n637) );
  NAND2_X1 U533 ( .A1(n432), .A2(n759), .ZN(n431) );
  INV_X1 U534 ( .A(KEYINPUT83), .ZN(n433) );
  NOR2_X2 U535 ( .A1(n684), .A2(n683), .ZN(n685) );
  AND2_X1 U536 ( .A1(n533), .A2(KEYINPUT68), .ZN(n434) );
  XOR2_X1 U537 ( .A(n662), .B(n664), .Z(n435) );
  XOR2_X1 U538 ( .A(KEYINPUT100), .B(n625), .Z(n436) );
  INV_X1 U539 ( .A(KEYINPUT82), .ZN(n567) );
  NAND2_X1 U540 ( .A1(n551), .A2(KEYINPUT44), .ZN(n552) );
  XNOR2_X1 U541 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U542 ( .A(KEYINPUT71), .B(KEYINPUT48), .ZN(n623) );
  AND2_X1 U543 ( .A1(n603), .A2(n601), .ZN(n578) );
  INV_X1 U544 ( .A(n683), .ZN(n654) );
  XNOR2_X1 U545 ( .A(KEYINPUT40), .B(KEYINPUT101), .ZN(n618) );
  INV_X1 U546 ( .A(KEYINPUT10), .ZN(n437) );
  XNOR2_X1 U547 ( .A(G137), .B(G140), .ZN(n438) );
  XOR2_X1 U548 ( .A(KEYINPUT78), .B(KEYINPUT75), .Z(n440) );
  XNOR2_X1 U549 ( .A(G128), .B(KEYINPUT24), .ZN(n439) );
  NAND2_X1 U550 ( .A1(n772), .A2(G234), .ZN(n441) );
  XOR2_X1 U551 ( .A(KEYINPUT91), .B(KEYINPUT92), .Z(n443) );
  XNOR2_X1 U552 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U553 ( .A(n444), .B(KEYINPUT23), .ZN(n445) );
  NOR2_X1 U554 ( .A1(G902), .A2(n658), .ZN(n449) );
  XNOR2_X1 U555 ( .A(KEYINPUT15), .B(G902), .ZN(n635) );
  NAND2_X1 U556 ( .A1(n635), .A2(G234), .ZN(n446) );
  XNOR2_X1 U557 ( .A(n446), .B(KEYINPUT20), .ZN(n450) );
  NAND2_X1 U558 ( .A1(n450), .A2(G217), .ZN(n447) );
  XNOR2_X2 U559 ( .A(n449), .B(n448), .ZN(n603) );
  INV_X1 U560 ( .A(n603), .ZN(n455) );
  NAND2_X1 U561 ( .A1(n450), .A2(G221), .ZN(n452) );
  INV_X1 U562 ( .A(KEYINPUT21), .ZN(n451) );
  XNOR2_X1 U563 ( .A(n452), .B(n451), .ZN(n714) );
  INV_X1 U564 ( .A(KEYINPUT94), .ZN(n453) );
  XNOR2_X1 U565 ( .A(n714), .B(n453), .ZN(n536) );
  INV_X1 U566 ( .A(n536), .ZN(n454) );
  AND2_X1 U567 ( .A1(n455), .A2(n454), .ZN(n561) );
  XNOR2_X2 U568 ( .A(KEYINPUT64), .B(G143), .ZN(n457) );
  XNOR2_X2 U569 ( .A(n457), .B(n456), .ZN(n518) );
  XNOR2_X1 U570 ( .A(G134), .B(G131), .ZN(n458) );
  XNOR2_X2 U571 ( .A(n767), .B(G146), .ZN(n475) );
  XNOR2_X1 U572 ( .A(n459), .B(n487), .ZN(n463) );
  XOR2_X1 U573 ( .A(G101), .B(KEYINPUT79), .Z(n461) );
  NAND2_X1 U574 ( .A1(G227), .A2(n772), .ZN(n460) );
  XNOR2_X1 U575 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U576 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U577 ( .A(n475), .B(n464), .ZN(n676) );
  XNOR2_X2 U578 ( .A(n465), .B(G469), .ZN(n560) );
  XNOR2_X1 U579 ( .A(KEYINPUT66), .B(KEYINPUT1), .ZN(n466) );
  XOR2_X1 U580 ( .A(KEYINPUT5), .B(G137), .Z(n468) );
  NAND2_X1 U581 ( .A1(n509), .A2(G210), .ZN(n467) );
  XNOR2_X1 U582 ( .A(n468), .B(n467), .ZN(n473) );
  XNOR2_X1 U583 ( .A(n470), .B(n469), .ZN(n472) );
  XNOR2_X1 U584 ( .A(n472), .B(n471), .ZN(n489) );
  XNOR2_X1 U585 ( .A(n489), .B(n473), .ZN(n474) );
  XNOR2_X1 U586 ( .A(n475), .B(n474), .ZN(n662) );
  XNOR2_X1 U587 ( .A(KEYINPUT88), .B(KEYINPUT33), .ZN(n476) );
  XNOR2_X1 U588 ( .A(n479), .B(n478), .ZN(n483) );
  XNOR2_X1 U589 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U590 ( .A(n483), .B(n482), .ZN(n485) );
  XNOR2_X1 U591 ( .A(n484), .B(n485), .ZN(n490) );
  XNOR2_X1 U592 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U593 ( .A(n489), .B(n488), .ZN(n755) );
  INV_X1 U594 ( .A(n635), .ZN(n631) );
  INV_X1 U595 ( .A(G902), .ZN(n527) );
  INV_X1 U596 ( .A(G237), .ZN(n491) );
  NAND2_X1 U597 ( .A1(n527), .A2(n491), .ZN(n493) );
  NAND2_X1 U598 ( .A1(n493), .A2(G210), .ZN(n492) );
  NAND2_X1 U599 ( .A1(n493), .A2(G214), .ZN(n728) );
  NAND2_X1 U600 ( .A1(G234), .A2(G237), .ZN(n495) );
  XNOR2_X1 U601 ( .A(n495), .B(KEYINPUT14), .ZN(n743) );
  INV_X1 U602 ( .A(G952), .ZN(n496) );
  NAND2_X1 U603 ( .A1(n772), .A2(n496), .ZN(n498) );
  NAND2_X1 U604 ( .A1(G953), .A2(n527), .ZN(n497) );
  AND2_X1 U605 ( .A1(n498), .A2(n497), .ZN(n499) );
  AND2_X1 U606 ( .A1(n743), .A2(n499), .ZN(n575) );
  NAND2_X1 U607 ( .A1(G953), .A2(G898), .ZN(n500) );
  NAND2_X1 U608 ( .A1(n575), .A2(n500), .ZN(n501) );
  NOR2_X2 U609 ( .A1(n583), .A2(n501), .ZN(n502) );
  XNOR2_X2 U610 ( .A(n502), .B(KEYINPUT0), .ZN(n564) );
  NAND2_X1 U611 ( .A1(n737), .A2(n564), .ZN(n504) );
  XOR2_X1 U612 ( .A(KEYINPUT76), .B(KEYINPUT34), .Z(n503) );
  XNOR2_X1 U613 ( .A(n504), .B(n503), .ZN(n530) );
  XNOR2_X1 U614 ( .A(KEYINPUT97), .B(KEYINPUT96), .ZN(n505) );
  XNOR2_X1 U615 ( .A(G113), .B(G131), .ZN(n507) );
  XNOR2_X1 U616 ( .A(n508), .B(n507), .ZN(n516) );
  NAND2_X1 U617 ( .A1(G214), .A2(n509), .ZN(n515) );
  XNOR2_X1 U618 ( .A(n511), .B(n510), .ZN(n512) );
  XOR2_X1 U619 ( .A(KEYINPUT13), .B(G475), .Z(n517) );
  XNOR2_X1 U620 ( .A(G116), .B(G134), .ZN(n519) );
  XNOR2_X1 U621 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U622 ( .A(n518), .B(n521), .ZN(n526) );
  XOR2_X1 U623 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n524) );
  NAND2_X1 U624 ( .A1(G217), .A2(n522), .ZN(n523) );
  XNOR2_X1 U625 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U626 ( .A(n526), .B(n525), .ZN(n644) );
  NAND2_X1 U627 ( .A1(n644), .A2(n527), .ZN(n528) );
  AND2_X1 U628 ( .A1(n594), .A2(n565), .ZN(n529) );
  NAND2_X1 U629 ( .A1(n530), .A2(n529), .ZN(n532) );
  INV_X1 U630 ( .A(KEYINPUT35), .ZN(n531) );
  INV_X1 U631 ( .A(KEYINPUT44), .ZN(n533) );
  NAND2_X1 U632 ( .A1(n535), .A2(n534), .ZN(n547) );
  OR2_X1 U633 ( .A1(n594), .A2(n565), .ZN(n732) );
  NOR2_X1 U634 ( .A1(n732), .A2(n536), .ZN(n537) );
  NAND2_X1 U635 ( .A1(n564), .A2(n537), .ZN(n539) );
  INV_X1 U636 ( .A(KEYINPUT22), .ZN(n538) );
  XNOR2_X1 U637 ( .A(n603), .B(KEYINPUT99), .ZN(n713) );
  INV_X1 U638 ( .A(n389), .ZN(n718) );
  XNOR2_X2 U639 ( .A(n541), .B(KEYINPUT32), .ZN(n660) );
  NAND2_X1 U640 ( .A1(n603), .A2(n557), .ZN(n542) );
  NOR2_X1 U641 ( .A1(n389), .A2(n542), .ZN(n543) );
  AND2_X1 U642 ( .A1(n544), .A2(n543), .ZN(n695) );
  INV_X1 U643 ( .A(n695), .ZN(n545) );
  INV_X1 U644 ( .A(KEYINPUT68), .ZN(n548) );
  NOR2_X1 U645 ( .A1(n695), .A2(n548), .ZN(n549) );
  NAND2_X1 U646 ( .A1(n550), .A2(n660), .ZN(n551) );
  NAND2_X1 U647 ( .A1(n553), .A2(n718), .ZN(n554) );
  XNOR2_X1 U648 ( .A(n554), .B(KEYINPUT86), .ZN(n556) );
  INV_X1 U649 ( .A(n713), .ZN(n555) );
  INV_X1 U650 ( .A(n561), .ZN(n717) );
  NOR2_X1 U651 ( .A1(n717), .A2(n557), .ZN(n558) );
  AND2_X1 U652 ( .A1(n558), .A2(n389), .ZN(n722) );
  NAND2_X1 U653 ( .A1(n564), .A2(n722), .ZN(n559) );
  XNOR2_X1 U654 ( .A(n559), .B(KEYINPUT31), .ZN(n706) );
  NAND2_X1 U655 ( .A1(n561), .A2(n581), .ZN(n592) );
  NOR2_X1 U656 ( .A1(n592), .A2(n562), .ZN(n563) );
  AND2_X1 U657 ( .A1(n564), .A2(n563), .ZN(n692) );
  OR2_X1 U658 ( .A1(n706), .A2(n692), .ZN(n569) );
  INV_X1 U659 ( .A(n565), .ZN(n593) );
  AND2_X1 U660 ( .A1(n594), .A2(n593), .ZN(n703) );
  INV_X1 U661 ( .A(n594), .ZN(n566) );
  INV_X1 U662 ( .A(n588), .ZN(n568) );
  NAND2_X1 U663 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U664 ( .A(n570), .B(KEYINPUT98), .ZN(n571) );
  AND2_X1 U665 ( .A1(n686), .A2(n571), .ZN(n572) );
  INV_X1 U666 ( .A(n714), .ZN(n576) );
  NAND2_X1 U667 ( .A1(G953), .A2(G900), .ZN(n574) );
  NAND2_X1 U668 ( .A1(n575), .A2(n574), .ZN(n613) );
  NOR2_X1 U669 ( .A1(n576), .A2(n613), .ZN(n577) );
  XOR2_X1 U670 ( .A(n577), .B(KEYINPUT73), .Z(n601) );
  INV_X1 U671 ( .A(KEYINPUT28), .ZN(n579) );
  XNOR2_X1 U672 ( .A(n580), .B(n579), .ZN(n582) );
  NAND2_X1 U673 ( .A1(n582), .A2(n581), .ZN(n621) );
  BUF_X1 U674 ( .A(n583), .Z(n584) );
  NAND2_X1 U675 ( .A1(n701), .A2(n585), .ZN(n586) );
  XOR2_X1 U676 ( .A(KEYINPUT47), .B(KEYINPUT69), .Z(n587) );
  NAND2_X1 U677 ( .A1(n701), .A2(n589), .ZN(n600) );
  NAND2_X1 U678 ( .A1(n562), .A2(n728), .ZN(n590) );
  XNOR2_X1 U679 ( .A(n590), .B(KEYINPUT30), .ZN(n591) );
  NOR2_X1 U680 ( .A1(n593), .A2(n613), .ZN(n595) );
  NAND2_X1 U681 ( .A1(n595), .A2(n594), .ZN(n597) );
  NOR2_X1 U682 ( .A1(n597), .A2(n596), .ZN(n598) );
  AND2_X1 U683 ( .A1(n615), .A2(n598), .ZN(n700) );
  INV_X1 U684 ( .A(n700), .ZN(n599) );
  NAND2_X1 U685 ( .A1(n603), .A2(n602), .ZN(n604) );
  INV_X1 U686 ( .A(n606), .ZN(n607) );
  NAND2_X1 U687 ( .A1(n624), .A2(n607), .ZN(n609) );
  INV_X1 U688 ( .A(KEYINPUT36), .ZN(n608) );
  XNOR2_X1 U689 ( .A(n609), .B(n608), .ZN(n611) );
  XOR2_X1 U690 ( .A(KEYINPUT85), .B(KEYINPUT39), .Z(n617) );
  INV_X1 U691 ( .A(KEYINPUT38), .ZN(n612) );
  NOR2_X1 U692 ( .A1(n620), .A2(n613), .ZN(n614) );
  NAND2_X1 U693 ( .A1(n703), .A2(n628), .ZN(n619) );
  NAND2_X1 U694 ( .A1(n729), .A2(n728), .ZN(n733) );
  NOR2_X1 U695 ( .A1(n748), .A2(n621), .ZN(n622) );
  XNOR2_X1 U696 ( .A(n622), .B(KEYINPUT42), .ZN(n780) );
  NAND2_X1 U697 ( .A1(n624), .A2(n728), .ZN(n625) );
  NAND2_X1 U698 ( .A1(n436), .A2(n718), .ZN(n626) );
  XNOR2_X1 U699 ( .A(n626), .B(KEYINPUT43), .ZN(n627) );
  NAND2_X1 U700 ( .A1(n627), .A2(n596), .ZN(n650) );
  NAND2_X1 U701 ( .A1(n628), .A2(n705), .ZN(n711) );
  AND2_X1 U702 ( .A1(n650), .A2(n711), .ZN(n629) );
  NAND2_X1 U703 ( .A1(KEYINPUT2), .A2(KEYINPUT84), .ZN(n630) );
  INV_X1 U704 ( .A(KEYINPUT2), .ZN(n632) );
  NOR2_X1 U705 ( .A1(n632), .A2(KEYINPUT84), .ZN(n633) );
  NOR2_X1 U706 ( .A1(KEYINPUT83), .A2(n633), .ZN(n634) );
  NAND2_X1 U707 ( .A1(n635), .A2(n634), .ZN(n636) );
  NAND2_X1 U708 ( .A1(n637), .A2(n636), .ZN(n639) );
  NAND2_X1 U709 ( .A1(n712), .A2(KEYINPUT83), .ZN(n638) );
  NAND2_X1 U710 ( .A1(n639), .A2(n638), .ZN(n642) );
  INV_X1 U711 ( .A(n712), .ZN(n640) );
  NAND2_X1 U712 ( .A1(n640), .A2(KEYINPUT2), .ZN(n641) );
  NAND2_X1 U713 ( .A1(n675), .A2(G478), .ZN(n646) );
  XOR2_X1 U714 ( .A(KEYINPUT118), .B(n644), .Z(n645) );
  XNOR2_X1 U715 ( .A(n646), .B(n645), .ZN(n647) );
  NOR2_X2 U716 ( .A1(n647), .A2(n683), .ZN(n649) );
  INV_X1 U717 ( .A(KEYINPUT119), .ZN(n648) );
  XNOR2_X1 U718 ( .A(n649), .B(n648), .ZN(G63) );
  XNOR2_X1 U719 ( .A(n650), .B(G140), .ZN(G42) );
  NAND2_X1 U720 ( .A1(n354), .A2(G475), .ZN(n653) );
  XOR2_X1 U721 ( .A(KEYINPUT117), .B(KEYINPUT59), .Z(n651) );
  XNOR2_X1 U722 ( .A(n653), .B(n366), .ZN(n655) );
  XNOR2_X1 U723 ( .A(n360), .B(KEYINPUT60), .ZN(G60) );
  BUF_X1 U724 ( .A(n354), .Z(n656) );
  NAND2_X1 U725 ( .A1(n656), .A2(G217), .ZN(n657) );
  XNOR2_X1 U726 ( .A(n658), .B(n657), .ZN(n659) );
  NOR2_X1 U727 ( .A1(n659), .A2(n683), .ZN(G66) );
  XNOR2_X1 U728 ( .A(G119), .B(KEYINPUT125), .ZN(n661) );
  XOR2_X1 U729 ( .A(n661), .B(n660), .Z(G21) );
  NAND2_X1 U730 ( .A1(n354), .A2(G472), .ZN(n665) );
  XNOR2_X1 U731 ( .A(KEYINPUT102), .B(KEYINPUT103), .ZN(n663) );
  XOR2_X1 U732 ( .A(n663), .B(KEYINPUT62), .Z(n664) );
  XNOR2_X1 U733 ( .A(n665), .B(n435), .ZN(n666) );
  XNOR2_X1 U734 ( .A(KEYINPUT104), .B(KEYINPUT63), .ZN(n667) );
  XNOR2_X1 U735 ( .A(n667), .B(KEYINPUT89), .ZN(n668) );
  XNOR2_X1 U736 ( .A(n359), .B(n668), .ZN(G57) );
  NAND2_X1 U737 ( .A1(n354), .A2(G210), .ZN(n671) );
  XOR2_X1 U738 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n670) );
  XNOR2_X1 U739 ( .A(n671), .B(n367), .ZN(n672) );
  XNOR2_X1 U740 ( .A(n353), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U741 ( .A(G122), .B(KEYINPUT124), .ZN(n673) );
  XNOR2_X1 U742 ( .A(n674), .B(n673), .ZN(G24) );
  NAND2_X1 U743 ( .A1(n675), .A2(G469), .ZN(n682) );
  BUF_X1 U744 ( .A(n676), .Z(n680) );
  XOR2_X1 U745 ( .A(KEYINPUT115), .B(KEYINPUT114), .Z(n678) );
  XNOR2_X1 U746 ( .A(KEYINPUT58), .B(KEYINPUT57), .ZN(n677) );
  XOR2_X1 U747 ( .A(n678), .B(n677), .Z(n679) );
  XNOR2_X1 U748 ( .A(n682), .B(n681), .ZN(n684) );
  XNOR2_X1 U749 ( .A(n685), .B(KEYINPUT116), .ZN(G54) );
  XNOR2_X1 U750 ( .A(n686), .B(G101), .ZN(G3) );
  XOR2_X1 U751 ( .A(G104), .B(KEYINPUT105), .Z(n688) );
  NAND2_X1 U752 ( .A1(n692), .A2(n703), .ZN(n687) );
  XNOR2_X1 U753 ( .A(n688), .B(n687), .ZN(G6) );
  XOR2_X1 U754 ( .A(KEYINPUT107), .B(KEYINPUT27), .Z(n690) );
  XNOR2_X1 U755 ( .A(G107), .B(KEYINPUT26), .ZN(n689) );
  XNOR2_X1 U756 ( .A(n690), .B(n689), .ZN(n691) );
  XOR2_X1 U757 ( .A(KEYINPUT106), .B(n691), .Z(n694) );
  NAND2_X1 U758 ( .A1(n692), .A2(n705), .ZN(n693) );
  XNOR2_X1 U759 ( .A(n694), .B(n693), .ZN(G9) );
  XOR2_X1 U760 ( .A(G110), .B(n695), .Z(n696) );
  XNOR2_X1 U761 ( .A(KEYINPUT108), .B(n696), .ZN(G12) );
  XOR2_X1 U762 ( .A(KEYINPUT109), .B(KEYINPUT29), .Z(n698) );
  NAND2_X1 U763 ( .A1(n701), .A2(n705), .ZN(n697) );
  XNOR2_X1 U764 ( .A(n698), .B(n697), .ZN(n699) );
  XOR2_X1 U765 ( .A(G128), .B(n699), .Z(G30) );
  NAND2_X1 U766 ( .A1(n701), .A2(n703), .ZN(n702) );
  XNOR2_X1 U767 ( .A(n702), .B(G146), .ZN(G48) );
  NAND2_X1 U768 ( .A1(n706), .A2(n703), .ZN(n704) );
  XNOR2_X1 U769 ( .A(n704), .B(G113), .ZN(G15) );
  NAND2_X1 U770 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U771 ( .A(n707), .B(KEYINPUT110), .ZN(n708) );
  XNOR2_X1 U772 ( .A(G116), .B(n708), .ZN(G18) );
  XNOR2_X1 U773 ( .A(n709), .B(G125), .ZN(n710) );
  XNOR2_X1 U774 ( .A(n710), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U775 ( .A(G134), .B(n711), .ZN(G36) );
  XNOR2_X1 U776 ( .A(n712), .B(KEYINPUT2), .ZN(n753) );
  NOR2_X1 U777 ( .A1(n714), .A2(n713), .ZN(n715) );
  XOR2_X1 U778 ( .A(KEYINPUT49), .B(n715), .Z(n716) );
  NOR2_X1 U779 ( .A1(n716), .A2(n562), .ZN(n721) );
  NAND2_X1 U780 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U781 ( .A(n719), .B(KEYINPUT50), .ZN(n720) );
  NAND2_X1 U782 ( .A1(n721), .A2(n720), .ZN(n724) );
  INV_X1 U783 ( .A(n722), .ZN(n723) );
  NAND2_X1 U784 ( .A1(n724), .A2(n723), .ZN(n726) );
  XOR2_X1 U785 ( .A(KEYINPUT111), .B(KEYINPUT51), .Z(n725) );
  XNOR2_X1 U786 ( .A(n726), .B(n725), .ZN(n727) );
  NOR2_X1 U787 ( .A1(n727), .A2(n748), .ZN(n741) );
  NOR2_X1 U788 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U789 ( .A(n730), .B(KEYINPUT112), .ZN(n731) );
  NOR2_X1 U790 ( .A1(n732), .A2(n731), .ZN(n736) );
  NOR2_X1 U791 ( .A1(n734), .A2(n733), .ZN(n735) );
  NOR2_X1 U792 ( .A1(n736), .A2(n735), .ZN(n739) );
  BUF_X1 U793 ( .A(n737), .Z(n738) );
  INV_X1 U794 ( .A(n738), .ZN(n747) );
  NOR2_X1 U795 ( .A1(n739), .A2(n747), .ZN(n740) );
  NOR2_X1 U796 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U797 ( .A(KEYINPUT52), .B(n742), .ZN(n745) );
  NAND2_X1 U798 ( .A1(G952), .A2(n743), .ZN(n744) );
  NOR2_X1 U799 ( .A1(n745), .A2(n744), .ZN(n746) );
  NOR2_X1 U800 ( .A1(G953), .A2(n746), .ZN(n751) );
  NOR2_X1 U801 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U802 ( .A(n749), .B(KEYINPUT113), .ZN(n750) );
  NAND2_X1 U803 ( .A1(n751), .A2(n750), .ZN(n752) );
  NOR2_X1 U804 ( .A1(n753), .A2(n752), .ZN(n754) );
  XNOR2_X1 U805 ( .A(KEYINPUT53), .B(n754), .ZN(G75) );
  XOR2_X1 U806 ( .A(KEYINPUT121), .B(n755), .Z(n757) );
  NOR2_X1 U807 ( .A1(G898), .A2(n772), .ZN(n756) );
  NOR2_X1 U808 ( .A1(n757), .A2(n756), .ZN(n758) );
  XOR2_X1 U809 ( .A(KEYINPUT122), .B(n758), .Z(n766) );
  NAND2_X1 U810 ( .A1(n759), .A2(n772), .ZN(n760) );
  XNOR2_X1 U811 ( .A(n760), .B(KEYINPUT120), .ZN(n764) );
  NAND2_X1 U812 ( .A1(G953), .A2(G224), .ZN(n761) );
  XNOR2_X1 U813 ( .A(KEYINPUT61), .B(n761), .ZN(n762) );
  NAND2_X1 U814 ( .A1(n762), .A2(G898), .ZN(n763) );
  NAND2_X1 U815 ( .A1(n764), .A2(n763), .ZN(n765) );
  XOR2_X1 U816 ( .A(n766), .B(n765), .Z(G69) );
  BUF_X1 U817 ( .A(n767), .Z(n768) );
  XNOR2_X1 U818 ( .A(n769), .B(KEYINPUT123), .ZN(n770) );
  XNOR2_X1 U819 ( .A(n768), .B(n770), .ZN(n774) );
  XOR2_X1 U820 ( .A(n774), .B(n771), .Z(n773) );
  NAND2_X1 U821 ( .A1(n773), .A2(n772), .ZN(n778) );
  XNOR2_X1 U822 ( .A(G227), .B(n774), .ZN(n775) );
  NAND2_X1 U823 ( .A1(n775), .A2(G900), .ZN(n776) );
  NAND2_X1 U824 ( .A1(n776), .A2(G953), .ZN(n777) );
  NAND2_X1 U825 ( .A1(n778), .A2(n777), .ZN(G72) );
  XOR2_X1 U826 ( .A(G137), .B(KEYINPUT126), .Z(n779) );
  XNOR2_X1 U827 ( .A(n780), .B(n779), .ZN(G39) );
  XOR2_X1 U828 ( .A(G131), .B(n781), .Z(G33) );
endmodule

