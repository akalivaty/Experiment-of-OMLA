//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 0 1 1 1 1 0 0 0 1 0 0 0 1 0 0 1 0 1 1 0 0 1 1 0 0 0 0 0 1 1 1 1 0 0 1 1 1 1 1 1 1 0 0 1 0 0 0 1 0 1 0 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n632, new_n633, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n704, new_n706, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n800, new_n802, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n862, new_n863, new_n864, new_n866, new_n867, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n879, new_n880, new_n882, new_n883, new_n884, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT0), .ZN(new_n203));
  XOR2_X1   g002(.A(G57gat), .B(G85gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G162gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT74), .ZN(new_n208));
  INV_X1    g007(.A(G155gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(KEYINPUT74), .A2(G155gat), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n207), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT2), .ZN(new_n213));
  OAI21_X1  g012(.A(KEYINPUT75), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(new_n211), .ZN(new_n215));
  NOR2_X1   g014(.A1(KEYINPUT74), .A2(G155gat), .ZN(new_n216));
  OAI21_X1  g015(.A(G162gat), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT75), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n217), .A2(new_n218), .A3(KEYINPUT2), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n207), .A2(G155gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n209), .A2(G162gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OR2_X1    g021(.A1(KEYINPUT73), .A2(G148gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(KEYINPUT73), .A2(G148gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n223), .A2(G141gat), .A3(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(G141gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(G148gat), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n222), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  AND3_X1   g027(.A1(new_n214), .A2(new_n219), .A3(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(G141gat), .B(G148gat), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n222), .B1(new_n230), .B2(KEYINPUT2), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT72), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  OAI211_X1 g032(.A(new_n222), .B(KEYINPUT72), .C1(new_n230), .C2(KEYINPUT2), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  OAI21_X1  g034(.A(KEYINPUT3), .B1(new_n229), .B2(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n214), .A2(new_n228), .A3(new_n219), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n238));
  NAND4_X1  g037(.A1(new_n237), .A2(new_n238), .A3(new_n233), .A4(new_n234), .ZN(new_n239));
  INV_X1    g038(.A(G134gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(G127gat), .ZN(new_n241));
  INV_X1    g040(.A(G127gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(G134gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(G113gat), .B(G120gat), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n244), .B1(new_n245), .B2(KEYINPUT1), .ZN(new_n246));
  INV_X1    g045(.A(G120gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(G113gat), .ZN(new_n248));
  INV_X1    g047(.A(G113gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(G120gat), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(G127gat), .B(G134gat), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT1), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n251), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  AND2_X1   g053(.A1(new_n246), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n236), .A2(new_n239), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(G225gat), .A2(G233gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n258), .B(KEYINPUT76), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n237), .A2(new_n255), .A3(new_n233), .A4(new_n234), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT4), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n235), .ZN(new_n264));
  NAND4_X1  g063(.A1(new_n264), .A2(KEYINPUT4), .A3(new_n237), .A4(new_n255), .ZN(new_n265));
  NAND4_X1  g064(.A1(new_n257), .A2(new_n260), .A3(new_n263), .A4(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT5), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n206), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT78), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT77), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n266), .A2(new_n271), .ZN(new_n272));
  AND2_X1   g071(.A1(new_n263), .A2(new_n265), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n273), .A2(KEYINPUT77), .A3(new_n260), .A4(new_n257), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n255), .B1(new_n264), .B2(new_n237), .ZN(new_n276));
  INV_X1    g075(.A(new_n261), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n259), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(KEYINPUT5), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n270), .B1(new_n275), .B2(new_n280), .ZN(new_n281));
  AOI211_X1 g080(.A(KEYINPUT78), .B(new_n279), .C1(new_n272), .C2(new_n274), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n269), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT79), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  OAI211_X1 g084(.A(KEYINPUT79), .B(new_n269), .C1(new_n281), .C2(new_n282), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n267), .A2(new_n268), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n288), .B1(new_n281), .B2(new_n282), .ZN(new_n289));
  AOI21_X1  g088(.A(KEYINPUT6), .B1(new_n289), .B2(new_n206), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n287), .A2(new_n290), .ZN(new_n291));
  AND3_X1   g090(.A1(new_n289), .A2(KEYINPUT6), .A3(new_n206), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  XOR2_X1   g093(.A(G197gat), .B(G204gat), .Z(new_n295));
  AOI21_X1  g094(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(G211gat), .B(G218gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n297), .B(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(G226gat), .A2(G233gat), .ZN(new_n300));
  AND2_X1   g099(.A1(G183gat), .A2(G190gat), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT68), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n302), .B1(G169gat), .B2(G176gat), .ZN(new_n303));
  NOR3_X1   g102(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n304));
  MUX2_X1   g103(.A(new_n303), .B(new_n302), .S(new_n304), .Z(new_n305));
  OAI21_X1  g104(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n306));
  XOR2_X1   g105(.A(new_n306), .B(KEYINPUT67), .Z(new_n307));
  AOI21_X1  g106(.A(new_n301), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(KEYINPUT27), .B(G183gat), .ZN(new_n309));
  INV_X1    g108(.A(G190gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT28), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  XNOR2_X1  g112(.A(new_n309), .B(KEYINPUT66), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n310), .A2(KEYINPUT28), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n313), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n308), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT24), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n318), .A2(G183gat), .A3(G190gat), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n319), .B1(new_n301), .B2(new_n318), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n320), .B1(G183gat), .B2(G190gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(G169gat), .A2(G176gat), .ZN(new_n322));
  INV_X1    g121(.A(G169gat), .ZN(new_n323));
  INV_X1    g122(.A(G176gat), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n323), .A2(new_n324), .A3(KEYINPUT23), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT23), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n326), .B1(G169gat), .B2(G176gat), .ZN(new_n327));
  NAND4_X1  g126(.A1(new_n321), .A2(new_n322), .A3(new_n325), .A4(new_n327), .ZN(new_n328));
  OAI21_X1  g127(.A(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n329));
  OR3_X1    g128(.A1(KEYINPUT65), .A2(G183gat), .A3(G190gat), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n320), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n325), .A2(new_n327), .A3(new_n322), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n332), .A2(KEYINPUT25), .ZN(new_n333));
  AOI22_X1  g132(.A1(new_n328), .A2(KEYINPUT25), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n317), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(KEYINPUT69), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT69), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n317), .A2(new_n334), .A3(new_n337), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n300), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n300), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n340), .A2(KEYINPUT29), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n335), .A2(KEYINPUT71), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT71), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n317), .A2(new_n334), .A3(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n342), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n299), .B1(new_n339), .B2(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(KEYINPUT70), .B(KEYINPUT29), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n336), .A2(new_n300), .A3(new_n338), .A4(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n299), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n343), .A2(new_n340), .A3(new_n345), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n347), .A2(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(G8gat), .B(G36gat), .ZN(new_n354));
  XNOR2_X1  g153(.A(G64gat), .B(G92gat), .ZN(new_n355));
  XOR2_X1   g154(.A(new_n354), .B(new_n355), .Z(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  OR3_X1    g156(.A1(new_n353), .A2(KEYINPUT30), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n336), .A2(new_n338), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(new_n340), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n343), .A2(new_n345), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(new_n341), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n350), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  AND3_X1   g162(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n357), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n347), .A2(new_n352), .A3(new_n356), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n365), .A2(KEYINPUT30), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n358), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n294), .A2(KEYINPUT80), .A3(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT80), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n292), .B1(new_n287), .B2(new_n290), .ZN(new_n371));
  INV_X1    g170(.A(new_n368), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n370), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(new_n335), .B(new_n256), .ZN(new_n374));
  NAND2_X1  g173(.A1(G227gat), .A2(G233gat), .ZN(new_n375));
  XNOR2_X1  g174(.A(new_n375), .B(KEYINPUT64), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(KEYINPUT32), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n374), .A2(new_n376), .ZN(new_n379));
  XOR2_X1   g178(.A(new_n379), .B(KEYINPUT34), .Z(new_n380));
  XNOR2_X1  g179(.A(G15gat), .B(G43gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(G71gat), .B(G99gat), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n381), .B(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT33), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n383), .B1(new_n377), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n380), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n380), .A2(new_n385), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n378), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  OR2_X1    g188(.A1(new_n380), .A2(new_n385), .ZN(new_n390));
  INV_X1    g189(.A(new_n378), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n390), .A2(new_n386), .A3(new_n391), .ZN(new_n392));
  OR2_X1    g191(.A1(new_n350), .A2(KEYINPUT29), .ZN(new_n393));
  AOI22_X1  g192(.A1(new_n393), .A2(new_n238), .B1(new_n237), .B2(new_n264), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n299), .B1(new_n239), .B2(new_n348), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(G228gat), .A2(G233gat), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n299), .A2(KEYINPUT81), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n297), .A2(KEYINPUT81), .A3(new_n298), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(new_n348), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n238), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n401), .B1(new_n229), .B2(new_n235), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(new_n397), .ZN(new_n403));
  OAI22_X1  g202(.A1(new_n396), .A2(new_n397), .B1(new_n403), .B2(new_n395), .ZN(new_n404));
  INV_X1    g203(.A(G22gat), .ZN(new_n405));
  AND2_X1   g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n404), .A2(new_n405), .ZN(new_n407));
  XNOR2_X1  g206(.A(G78gat), .B(G106gat), .ZN(new_n408));
  XNOR2_X1  g207(.A(KEYINPUT31), .B(G50gat), .ZN(new_n409));
  XOR2_X1   g208(.A(new_n408), .B(new_n409), .Z(new_n410));
  XNOR2_X1  g209(.A(new_n410), .B(KEYINPUT82), .ZN(new_n411));
  OR3_X1    g210(.A1(new_n406), .A2(new_n407), .A3(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT82), .ZN(new_n413));
  OAI22_X1  g212(.A1(new_n406), .A2(new_n407), .B1(new_n413), .B2(new_n410), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  AND3_X1   g214(.A1(new_n389), .A2(new_n392), .A3(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n369), .A2(new_n373), .A3(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT35), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n415), .A2(new_n418), .ZN(new_n419));
  NOR3_X1   g218(.A1(new_n387), .A2(new_n388), .A3(new_n378), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n391), .B1(new_n390), .B2(new_n386), .ZN(new_n421));
  NOR4_X1   g220(.A1(new_n419), .A2(new_n420), .A3(new_n421), .A4(new_n372), .ZN(new_n422));
  AOI21_X1  g221(.A(KEYINPUT6), .B1(new_n285), .B2(new_n286), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT85), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n289), .A2(new_n424), .ZN(new_n425));
  OAI211_X1 g224(.A(KEYINPUT85), .B(new_n288), .C1(new_n281), .C2(new_n282), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n425), .A2(new_n206), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n423), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(KEYINPUT86), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT86), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n423), .A2(new_n430), .A3(new_n427), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n429), .A2(new_n293), .A3(new_n431), .ZN(new_n432));
  AOI22_X1  g231(.A1(new_n417), .A2(KEYINPUT35), .B1(new_n422), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT88), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n357), .A2(KEYINPUT37), .ZN(new_n435));
  AOI22_X1  g234(.A1(new_n365), .A2(new_n435), .B1(KEYINPUT37), .B2(new_n353), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT38), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n434), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n366), .ZN(new_n439));
  AOI21_X1  g238(.A(KEYINPUT38), .B1(new_n365), .B2(new_n435), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n350), .B1(new_n339), .B2(new_n346), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n349), .A2(new_n299), .A3(new_n351), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n441), .A2(KEYINPUT37), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(KEYINPUT87), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT87), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n441), .A2(new_n445), .A3(KEYINPUT37), .A4(new_n442), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n439), .B1(new_n440), .B2(new_n447), .ZN(new_n448));
  AND2_X1   g247(.A1(new_n353), .A2(KEYINPUT37), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n357), .B1(new_n353), .B2(KEYINPUT37), .ZN(new_n450));
  OAI211_X1 g249(.A(KEYINPUT88), .B(KEYINPUT38), .C1(new_n449), .C2(new_n450), .ZN(new_n451));
  AND3_X1   g250(.A1(new_n438), .A2(new_n448), .A3(new_n451), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n429), .A2(new_n293), .A3(new_n431), .A4(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n415), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n260), .B1(new_n273), .B2(new_n257), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT39), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n206), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  OR2_X1    g256(.A1(new_n276), .A2(new_n277), .ZN(new_n458));
  OAI21_X1  g257(.A(KEYINPUT39), .B1(new_n458), .B2(new_n259), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n457), .B1(new_n455), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT84), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  XNOR2_X1  g261(.A(new_n462), .B(KEYINPUT40), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n463), .A2(new_n368), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n454), .B1(new_n464), .B2(new_n427), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n453), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(KEYINPUT80), .B1(new_n294), .B2(new_n368), .ZN(new_n468));
  NOR3_X1   g267(.A1(new_n371), .A2(new_n370), .A3(new_n372), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n454), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT36), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n471), .B1(new_n420), .B2(new_n421), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n389), .A2(new_n392), .A3(KEYINPUT36), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n470), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT83), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n467), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n470), .A2(KEYINPUT83), .A3(new_n474), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n433), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(G29gat), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n480), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n481));
  XOR2_X1   g280(.A(KEYINPUT14), .B(G29gat), .Z(new_n482));
  OAI21_X1  g281(.A(new_n481), .B1(new_n482), .B2(G36gat), .ZN(new_n483));
  XNOR2_X1  g282(.A(G43gat), .B(G50gat), .ZN(new_n484));
  AOI22_X1  g283(.A1(new_n483), .A2(KEYINPUT89), .B1(KEYINPUT15), .B2(new_n484), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n483), .B1(KEYINPUT15), .B2(new_n484), .ZN(new_n486));
  OR2_X1    g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n485), .A2(new_n486), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  OR2_X1    g288(.A1(new_n489), .A2(KEYINPUT17), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT90), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n490), .B(new_n491), .ZN(new_n492));
  AND2_X1   g291(.A1(new_n489), .A2(KEYINPUT17), .ZN(new_n493));
  XNOR2_X1  g292(.A(G15gat), .B(G22gat), .ZN(new_n494));
  OR2_X1    g293(.A1(new_n494), .A2(G1gat), .ZN(new_n495));
  INV_X1    g294(.A(G8gat), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT16), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n494), .B1(new_n497), .B2(G1gat), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n495), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  XNOR2_X1  g298(.A(new_n499), .B(KEYINPUT92), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n495), .A2(KEYINPUT91), .A3(new_n498), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n501), .B(G8gat), .C1(KEYINPUT91), .C2(new_n498), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n493), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n492), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(G229gat), .A2(G233gat), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n506), .B(KEYINPUT93), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n489), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(new_n503), .ZN(new_n510));
  AND3_X1   g309(.A1(new_n505), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(KEYINPUT18), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT94), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n511), .A2(KEYINPUT94), .A3(KEYINPUT18), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n511), .A2(KEYINPUT18), .ZN(new_n517));
  XOR2_X1   g316(.A(KEYINPUT95), .B(KEYINPUT13), .Z(new_n518));
  XNOR2_X1  g317(.A(new_n507), .B(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(KEYINPUT96), .B1(new_n509), .B2(new_n503), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n509), .A2(new_n503), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n520), .B(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n517), .B1(new_n519), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n516), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(G113gat), .B(G141gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n525), .B(G197gat), .ZN(new_n526));
  XOR2_X1   g325(.A(KEYINPUT11), .B(G169gat), .Z(new_n527));
  XNOR2_X1  g326(.A(new_n526), .B(new_n527), .ZN(new_n528));
  XOR2_X1   g327(.A(new_n528), .B(KEYINPUT12), .Z(new_n529));
  NAND2_X1  g328(.A1(new_n524), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n529), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n516), .A2(new_n523), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n479), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(G85gat), .A2(G92gat), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n536), .B(KEYINPUT7), .ZN(new_n537));
  NAND2_X1  g336(.A1(G99gat), .A2(G106gat), .ZN(new_n538));
  INV_X1    g337(.A(G85gat), .ZN(new_n539));
  INV_X1    g338(.A(G92gat), .ZN(new_n540));
  AOI22_X1  g339(.A1(KEYINPUT8), .A2(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT101), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n542), .B(new_n543), .ZN(new_n544));
  XOR2_X1   g343(.A(G99gat), .B(G106gat), .Z(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n542), .B(KEYINPUT101), .ZN(new_n547));
  INV_X1    g346(.A(new_n545), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  AND2_X1   g349(.A1(G232gat), .A2(G233gat), .ZN(new_n551));
  AOI22_X1  g350(.A1(new_n509), .A2(new_n550), .B1(KEYINPUT41), .B2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n550), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n493), .B1(KEYINPUT102), .B2(new_n553), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n554), .B1(KEYINPUT102), .B2(new_n553), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n490), .B(KEYINPUT90), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n552), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  XOR2_X1   g356(.A(G190gat), .B(G218gat), .Z(new_n558));
  XNOR2_X1  g357(.A(new_n557), .B(new_n558), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n551), .A2(KEYINPUT41), .ZN(new_n560));
  XNOR2_X1  g359(.A(G134gat), .B(G162gat), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n560), .B(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n559), .B(new_n562), .ZN(new_n563));
  XOR2_X1   g362(.A(G57gat), .B(G64gat), .Z(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  OR2_X1    g364(.A1(new_n565), .A2(KEYINPUT99), .ZN(new_n566));
  AOI21_X1  g365(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n567));
  XOR2_X1   g366(.A(new_n567), .B(KEYINPUT98), .Z(new_n568));
  XNOR2_X1  g367(.A(G71gat), .B(G78gat), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n565), .A2(KEYINPUT99), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n566), .A2(new_n568), .A3(new_n569), .A4(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n568), .A2(new_n564), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT97), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n573), .B1(G71gat), .B2(G78gat), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n574), .B1(new_n569), .B2(new_n573), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n571), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT21), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(G231gat), .A2(G233gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(G127gat), .ZN(new_n582));
  XOR2_X1   g381(.A(G183gat), .B(G211gat), .Z(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  OAI211_X1 g383(.A(new_n500), .B(new_n502), .C1(new_n577), .C2(new_n578), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(KEYINPUT100), .ZN(new_n586));
  XNOR2_X1  g385(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n587), .B(new_n209), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n586), .B(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n584), .B(new_n589), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n563), .A2(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n550), .B(new_n577), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT10), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND4_X1  g393(.A1(new_n550), .A2(KEYINPUT10), .A3(new_n576), .A4(new_n571), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(G230gat), .A2(G233gat), .ZN(new_n597));
  XOR2_X1   g396(.A(new_n597), .B(KEYINPUT103), .Z(new_n598));
  AND2_X1   g397(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n592), .A2(new_n598), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  XOR2_X1   g400(.A(G120gat), .B(G148gat), .Z(new_n602));
  XNOR2_X1  g401(.A(G176gat), .B(G204gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  OR2_X1    g403(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n601), .A2(new_n604), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n606), .A2(KEYINPUT104), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT104), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n608), .B1(new_n601), .B2(new_n604), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n605), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n591), .A2(new_n611), .ZN(new_n612));
  XOR2_X1   g411(.A(new_n612), .B(KEYINPUT105), .Z(new_n613));
  NAND2_X1  g412(.A1(new_n535), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(new_n371), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g416(.A(KEYINPUT16), .B(G8gat), .Z(new_n618));
  NAND3_X1  g417(.A1(new_n615), .A2(new_n372), .A3(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(KEYINPUT42), .ZN(new_n620));
  OAI21_X1  g419(.A(G8gat), .B1(new_n614), .B2(new_n368), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(KEYINPUT106), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n620), .A2(new_n622), .ZN(G1325gat));
  AND2_X1   g422(.A1(new_n472), .A2(new_n473), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(KEYINPUT107), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  OAI21_X1  g425(.A(G15gat), .B1(new_n614), .B2(new_n626), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n420), .A2(new_n421), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  OR2_X1    g428(.A1(new_n629), .A2(G15gat), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n627), .B1(new_n614), .B2(new_n630), .ZN(G1326gat));
  NOR2_X1   g430(.A1(new_n614), .A2(new_n415), .ZN(new_n632));
  XOR2_X1   g431(.A(KEYINPUT43), .B(G22gat), .Z(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(G1327gat));
  INV_X1    g433(.A(new_n563), .ZN(new_n635));
  INV_X1    g434(.A(new_n590), .ZN(new_n636));
  NOR3_X1   g435(.A1(new_n635), .A2(new_n636), .A3(new_n610), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(KEYINPUT108), .ZN(new_n638));
  AND2_X1   g437(.A1(new_n535), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n639), .A2(new_n480), .A3(new_n371), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(KEYINPUT45), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n533), .A2(new_n590), .A3(new_n611), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT44), .ZN(new_n643));
  AND3_X1   g442(.A1(new_n470), .A2(new_n466), .A3(new_n474), .ZN(new_n644));
  OAI211_X1 g443(.A(new_n643), .B(new_n563), .C1(new_n644), .C2(new_n433), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(KEYINPUT109), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n417), .A2(KEYINPUT35), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n422), .A2(new_n432), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n470), .A2(new_n466), .A3(new_n474), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n635), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT109), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n651), .A2(new_n652), .A3(new_n643), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n646), .A2(new_n653), .ZN(new_n654));
  OAI21_X1  g453(.A(KEYINPUT44), .B1(new_n479), .B2(new_n635), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n642), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  AND2_X1   g455(.A1(new_n656), .A2(new_n371), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n641), .B1(new_n480), .B2(new_n657), .ZN(G1328gat));
  INV_X1    g457(.A(G36gat), .ZN(new_n659));
  NAND4_X1  g458(.A1(new_n535), .A2(new_n659), .A3(new_n372), .A4(new_n638), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(KEYINPUT46), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n659), .B1(new_n656), .B2(new_n372), .ZN(new_n662));
  OR3_X1    g461(.A1(new_n661), .A2(KEYINPUT110), .A3(new_n662), .ZN(new_n663));
  OAI21_X1  g462(.A(KEYINPUT110), .B1(new_n661), .B2(new_n662), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(G1329gat));
  NAND2_X1  g464(.A1(new_n656), .A2(new_n625), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(G43gat), .ZN(new_n667));
  INV_X1    g466(.A(G43gat), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n639), .A2(new_n668), .A3(new_n628), .ZN(new_n669));
  AND2_X1   g468(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n668), .B1(new_n656), .B2(new_n624), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n669), .A2(KEYINPUT47), .ZN(new_n672));
  OAI22_X1  g471(.A1(new_n670), .A2(KEYINPUT47), .B1(new_n671), .B2(new_n672), .ZN(G1330gat));
  INV_X1    g472(.A(KEYINPUT48), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n415), .A2(G50gat), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n639), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(G50gat), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n677), .B1(new_n656), .B2(new_n454), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT111), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n676), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  AOI211_X1 g479(.A(KEYINPUT111), .B(new_n677), .C1(new_n656), .C2(new_n454), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n674), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT112), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n674), .B1(new_n639), .B2(new_n675), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n683), .B1(new_n685), .B2(new_n678), .ZN(new_n686));
  AND2_X1   g485(.A1(new_n656), .A2(new_n454), .ZN(new_n687));
  OAI211_X1 g486(.A(KEYINPUT112), .B(new_n684), .C1(new_n687), .C2(new_n677), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n682), .A2(new_n689), .ZN(G1331gat));
  NAND2_X1  g489(.A1(new_n649), .A2(new_n650), .ZN(new_n691));
  NOR4_X1   g490(.A1(new_n533), .A2(new_n590), .A3(new_n563), .A4(new_n611), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(new_n371), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g495(.A1(new_n693), .A2(new_n368), .ZN(new_n697));
  NOR2_X1   g496(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n698));
  AND2_X1   g497(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n697), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n700), .B1(new_n697), .B2(new_n698), .ZN(G1333gat));
  NOR3_X1   g500(.A1(new_n693), .A2(G71gat), .A3(new_n629), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n694), .A2(new_n625), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n702), .B1(G71gat), .B2(new_n703), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g504(.A1(new_n694), .A2(new_n454), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g506(.A1(new_n533), .A2(new_n636), .ZN(new_n708));
  INV_X1    g507(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n709), .A2(new_n611), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n711), .B1(new_n654), .B2(new_n655), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(new_n371), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT113), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n539), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n715), .B1(new_n714), .B2(new_n713), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n691), .A2(new_n563), .A3(new_n708), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT51), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n651), .A2(KEYINPUT51), .A3(new_n708), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n721), .A2(new_n539), .A3(new_n371), .A4(new_n610), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n716), .A2(new_n722), .ZN(G1336gat));
  INV_X1    g522(.A(new_n721), .ZN(new_n724));
  NOR4_X1   g523(.A1(new_n724), .A2(G92gat), .A3(new_n368), .A4(new_n611), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n540), .B1(new_n712), .B2(new_n372), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT52), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n727), .B(new_n728), .ZN(G1337gat));
  AND2_X1   g528(.A1(new_n712), .A2(new_n625), .ZN(new_n730));
  INV_X1    g529(.A(G99gat), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n628), .A2(new_n610), .A3(new_n731), .ZN(new_n732));
  XOR2_X1   g531(.A(new_n732), .B(KEYINPUT114), .Z(new_n733));
  OAI22_X1  g532(.A1(new_n730), .A2(new_n731), .B1(new_n724), .B2(new_n733), .ZN(G1338gat));
  NOR2_X1   g533(.A1(new_n415), .A2(G106gat), .ZN(new_n735));
  AND3_X1   g534(.A1(new_n651), .A2(KEYINPUT51), .A3(new_n708), .ZN(new_n736));
  AOI21_X1  g535(.A(KEYINPUT51), .B1(new_n651), .B2(new_n708), .ZN(new_n737));
  OAI211_X1 g536(.A(new_n610), .B(new_n735), .C1(new_n736), .C2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  AND4_X1   g538(.A1(new_n652), .A2(new_n691), .A3(new_n643), .A4(new_n563), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n652), .B1(new_n651), .B2(new_n643), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n415), .B1(new_n369), .B2(new_n373), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n476), .B1(new_n742), .B2(new_n624), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n478), .A2(new_n743), .A3(new_n466), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n635), .B1(new_n744), .B2(new_n649), .ZN(new_n745));
  OAI22_X1  g544(.A1(new_n740), .A2(new_n741), .B1(new_n643), .B2(new_n745), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n746), .A2(new_n454), .A3(new_n710), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n739), .B1(new_n747), .B2(G106gat), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT53), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n738), .A2(KEYINPUT115), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT115), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n721), .A2(new_n751), .A3(new_n610), .A4(new_n735), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n750), .A2(new_n749), .A3(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(G106gat), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n754), .B1(new_n712), .B2(new_n454), .ZN(new_n755));
  OAI22_X1  g554(.A1(new_n748), .A2(new_n749), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT116), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(KEYINPUT53), .B1(new_n755), .B2(new_n739), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n747), .A2(G106gat), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n760), .A2(new_n749), .A3(new_n750), .A4(new_n752), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n759), .A2(new_n761), .A3(KEYINPUT116), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n758), .A2(new_n762), .ZN(G1339gat));
  NOR2_X1   g562(.A1(new_n612), .A2(new_n533), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n508), .B1(new_n505), .B2(new_n510), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n522), .A2(new_n519), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n528), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n532), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n606), .B(KEYINPUT104), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT117), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT54), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n604), .B1(new_n599), .B2(new_n772), .ZN(new_n773));
  OR2_X1    g572(.A1(new_n596), .A2(new_n598), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n596), .A2(new_n598), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n774), .A2(KEYINPUT54), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n773), .A2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT55), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n771), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(new_n777), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n780), .A2(KEYINPUT117), .A3(KEYINPUT55), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n770), .A2(new_n779), .A3(new_n781), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n780), .A2(KEYINPUT55), .ZN(new_n783));
  NOR4_X1   g582(.A1(new_n769), .A2(new_n782), .A3(new_n635), .A4(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n532), .A2(new_n610), .A3(new_n768), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(KEYINPUT118), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT118), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n532), .A2(new_n610), .A3(new_n787), .A4(new_n768), .ZN(new_n788));
  INV_X1    g587(.A(new_n783), .ZN(new_n789));
  AND3_X1   g588(.A1(new_n516), .A2(new_n523), .A3(new_n531), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n531), .B1(new_n516), .B2(new_n523), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n789), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  OAI211_X1 g591(.A(new_n786), .B(new_n788), .C1(new_n792), .C2(new_n782), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n784), .B1(new_n793), .B2(new_n635), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n765), .B1(new_n794), .B2(new_n636), .ZN(new_n795));
  AND3_X1   g594(.A1(new_n795), .A2(new_n371), .A3(new_n415), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n796), .A2(new_n368), .A3(new_n628), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n797), .A2(new_n534), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n798), .B(new_n249), .ZN(G1340gat));
  NOR2_X1   g598(.A1(new_n797), .A2(new_n611), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n800), .B(new_n247), .ZN(G1341gat));
  NOR2_X1   g600(.A1(new_n797), .A2(new_n590), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n802), .B(new_n242), .ZN(G1342gat));
  NOR2_X1   g602(.A1(new_n635), .A2(new_n372), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n796), .A2(new_n240), .A3(new_n628), .A4(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT120), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n805), .B1(new_n806), .B2(KEYINPUT56), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT56), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n807), .B1(KEYINPUT120), .B2(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n805), .A2(new_n806), .A3(KEYINPUT56), .ZN(new_n810));
  OAI21_X1  g609(.A(G134gat), .B1(new_n797), .B2(new_n635), .ZN(new_n811));
  AND2_X1   g610(.A1(new_n811), .A2(KEYINPUT119), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT119), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n813), .B(G134gat), .C1(new_n797), .C2(new_n635), .ZN(new_n814));
  INV_X1    g613(.A(new_n814), .ZN(new_n815));
  OAI211_X1 g614(.A(new_n809), .B(new_n810), .C1(new_n812), .C2(new_n815), .ZN(G1343gat));
  INV_X1    g615(.A(new_n785), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n783), .B1(new_n530), .B2(new_n532), .ZN(new_n818));
  INV_X1    g617(.A(new_n782), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n817), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n819), .A2(new_n563), .A3(new_n789), .ZN(new_n821));
  OAI22_X1  g620(.A1(new_n820), .A2(new_n563), .B1(new_n769), .B2(new_n821), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n764), .B1(new_n822), .B2(new_n590), .ZN(new_n823));
  OAI21_X1  g622(.A(KEYINPUT57), .B1(new_n823), .B2(new_n415), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT57), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n795), .A2(new_n825), .A3(new_n454), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n624), .A2(new_n294), .A3(new_n372), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n824), .A2(new_n826), .A3(new_n533), .A4(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT121), .ZN(new_n829));
  AND3_X1   g628(.A1(new_n828), .A2(new_n829), .A3(G141gat), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n829), .B1(new_n828), .B2(G141gat), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n625), .A2(new_n294), .ZN(new_n832));
  AND3_X1   g631(.A1(new_n795), .A2(new_n454), .A3(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT122), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n534), .A2(G141gat), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n833), .A2(new_n834), .A3(new_n368), .A4(new_n835), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n795), .A2(new_n368), .A3(new_n454), .A4(new_n832), .ZN(new_n837));
  INV_X1    g636(.A(new_n835), .ZN(new_n838));
  OAI21_X1  g637(.A(KEYINPUT122), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n830), .A2(new_n831), .A3(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT58), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n828), .A2(G141gat), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n837), .A2(new_n838), .ZN(new_n844));
  XOR2_X1   g643(.A(KEYINPUT123), .B(KEYINPUT58), .Z(new_n845));
  NOR2_X1   g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(KEYINPUT124), .B1(new_n843), .B2(new_n846), .ZN(new_n847));
  AND3_X1   g646(.A1(new_n843), .A2(new_n846), .A3(KEYINPUT124), .ZN(new_n848));
  OAI22_X1  g647(.A1(new_n841), .A2(new_n842), .B1(new_n847), .B2(new_n848), .ZN(G1344gat));
  NAND2_X1  g648(.A1(new_n822), .A2(new_n590), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n613), .A2(new_n534), .ZN(new_n851));
  AOI211_X1 g650(.A(KEYINPUT57), .B(new_n415), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n825), .B1(new_n795), .B2(new_n454), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n854), .A2(new_n610), .A3(new_n827), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n855), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n856));
  OAI21_X1  g655(.A(KEYINPUT59), .B1(new_n837), .B2(new_n611), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n857), .A2(new_n223), .A3(new_n224), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n824), .A2(new_n826), .A3(new_n827), .ZN(new_n859));
  OR3_X1    g658(.A1(new_n859), .A2(KEYINPUT59), .A3(new_n611), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n856), .A2(new_n858), .A3(new_n860), .ZN(G1345gat));
  NAND2_X1  g660(.A1(new_n210), .A2(new_n211), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n862), .B1(new_n859), .B2(new_n590), .ZN(new_n863));
  OR2_X1    g662(.A1(new_n590), .A2(new_n862), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n863), .B1(new_n837), .B2(new_n864), .ZN(G1346gat));
  OAI21_X1  g664(.A(G162gat), .B1(new_n859), .B2(new_n635), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n833), .A2(new_n207), .A3(new_n804), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(G1347gat));
  AND2_X1   g667(.A1(new_n795), .A2(new_n415), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n371), .A2(new_n368), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n870), .A2(new_n628), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n872), .A2(new_n323), .A3(new_n534), .ZN(new_n873));
  AND2_X1   g672(.A1(new_n795), .A2(new_n294), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n874), .A2(new_n372), .A3(new_n416), .ZN(new_n875));
  XNOR2_X1  g674(.A(new_n875), .B(KEYINPUT125), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(new_n533), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n873), .B1(new_n877), .B2(new_n323), .ZN(G1348gat));
  NAND3_X1  g677(.A1(new_n876), .A2(new_n324), .A3(new_n610), .ZN(new_n879));
  OAI21_X1  g678(.A(G176gat), .B1(new_n872), .B2(new_n611), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(G1349gat));
  OAI21_X1  g680(.A(G183gat), .B1(new_n872), .B2(new_n590), .ZN(new_n882));
  OR2_X1    g681(.A1(new_n590), .A2(new_n314), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n882), .B1(new_n875), .B2(new_n883), .ZN(new_n884));
  XNOR2_X1  g683(.A(new_n884), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g684(.A1(new_n876), .A2(new_n310), .A3(new_n563), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT126), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n869), .A2(new_n563), .A3(new_n871), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT61), .ZN(new_n889));
  AND4_X1   g688(.A1(new_n887), .A2(new_n888), .A3(new_n889), .A4(G190gat), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n310), .B1(KEYINPUT126), .B2(KEYINPUT61), .ZN(new_n891));
  AOI22_X1  g690(.A1(new_n888), .A2(new_n891), .B1(new_n887), .B2(new_n889), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n886), .B1(new_n890), .B2(new_n892), .ZN(G1351gat));
  NOR3_X1   g692(.A1(new_n625), .A2(new_n368), .A3(new_n415), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n874), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g694(.A(G197gat), .B1(new_n895), .B2(new_n533), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n626), .A2(new_n870), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n852), .A2(new_n853), .A3(new_n897), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n533), .A2(G197gat), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n896), .B1(new_n898), .B2(new_n899), .ZN(G1352gat));
  INV_X1    g699(.A(G204gat), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n895), .A2(new_n901), .A3(new_n610), .ZN(new_n902));
  OR2_X1    g701(.A1(new_n902), .A2(KEYINPUT62), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(KEYINPUT62), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n898), .A2(new_n610), .ZN(new_n905));
  OAI211_X1 g704(.A(new_n903), .B(new_n904), .C1(new_n901), .C2(new_n905), .ZN(G1353gat));
  INV_X1    g705(.A(G211gat), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n895), .A2(new_n907), .A3(new_n636), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n898), .A2(new_n636), .ZN(new_n909));
  AND3_X1   g708(.A1(new_n909), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n910));
  AOI21_X1  g709(.A(KEYINPUT63), .B1(new_n909), .B2(G211gat), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n908), .B1(new_n910), .B2(new_n911), .ZN(G1354gat));
  INV_X1    g711(.A(G218gat), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n895), .A2(new_n913), .A3(new_n563), .ZN(new_n914));
  NOR4_X1   g713(.A1(new_n852), .A2(new_n853), .A3(new_n635), .A4(new_n897), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n914), .B1(new_n915), .B2(new_n913), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT127), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI211_X1 g717(.A(new_n914), .B(KEYINPUT127), .C1(new_n915), .C2(new_n913), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(G1355gat));
endmodule


