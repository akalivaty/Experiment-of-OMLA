//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 1 1 1 0 0 1 1 0 0 1 0 1 1 1 0 1 0 0 0 1 1 1 1 0 0 1 1 1 0 0 0 0 1 0 1 1 0 0 1 0 0 0 0 0 1 1 0 1 1 0 1 0 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:19 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n726, new_n727, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993;
  INV_X1    g000(.A(KEYINPUT98), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT12), .ZN(new_n188));
  INV_X1    g002(.A(G104), .ZN(new_n189));
  OAI21_X1  g003(.A(KEYINPUT3), .B1(new_n189), .B2(G107), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT3), .ZN(new_n191));
  INV_X1    g005(.A(G107), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n191), .A2(new_n192), .A3(G104), .ZN(new_n193));
  INV_X1    g007(.A(G101), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n189), .A2(G107), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n190), .A2(new_n193), .A3(new_n194), .A4(new_n195), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n189), .A2(G107), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n192), .A2(G104), .ZN(new_n198));
  OAI21_X1  g012(.A(G101), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  AND2_X1   g013(.A1(new_n196), .A2(new_n199), .ZN(new_n200));
  XNOR2_X1  g014(.A(G143), .B(G146), .ZN(new_n201));
  INV_X1    g015(.A(G128), .ZN(new_n202));
  INV_X1    g016(.A(G143), .ZN(new_n203));
  OAI21_X1  g017(.A(KEYINPUT1), .B1(new_n203), .B2(G146), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT81), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n202), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G146), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G143), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n208), .A2(KEYINPUT81), .A3(KEYINPUT1), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n201), .B1(new_n206), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT1), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n203), .A2(G146), .ZN(new_n212));
  AND4_X1   g026(.A1(new_n211), .A2(new_n208), .A3(new_n212), .A4(G128), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n200), .B1(new_n210), .B2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(new_n213), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n196), .A2(new_n199), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n202), .B1(new_n208), .B2(KEYINPUT1), .ZN(new_n217));
  NOR3_X1   g031(.A1(new_n217), .A2(new_n201), .A3(KEYINPUT66), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT66), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n204), .A2(G128), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n208), .A2(new_n212), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n219), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n215), .B(new_n216), .C1(new_n218), .C2(new_n222), .ZN(new_n223));
  AND2_X1   g037(.A1(new_n214), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT11), .ZN(new_n225));
  INV_X1    g039(.A(G134), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n225), .B1(new_n226), .B2(G137), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(G137), .ZN(new_n228));
  INV_X1    g042(.A(G137), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n229), .A2(KEYINPUT11), .A3(G134), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n227), .A2(new_n228), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G131), .ZN(new_n232));
  XNOR2_X1  g046(.A(KEYINPUT65), .B(G131), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n233), .A2(new_n227), .A3(new_n228), .A4(new_n230), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n188), .B1(new_n224), .B2(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n236), .B1(new_n214), .B2(new_n223), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(KEYINPUT12), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n237), .A2(KEYINPUT83), .A3(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT83), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n238), .A2(KEYINPUT12), .ZN(new_n242));
  AOI211_X1 g056(.A(new_n188), .B(new_n236), .C1(new_n214), .C2(new_n223), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n241), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n240), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n190), .A2(new_n193), .A3(new_n195), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(KEYINPUT79), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT79), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n190), .A2(new_n193), .A3(new_n249), .A4(new_n195), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n247), .A2(new_n248), .A3(G101), .A4(new_n250), .ZN(new_n251));
  AND4_X1   g065(.A1(KEYINPUT0), .A2(new_n208), .A3(new_n212), .A4(G128), .ZN(new_n252));
  XNOR2_X1  g066(.A(KEYINPUT0), .B(G128), .ZN(new_n253));
  OAI21_X1  g067(.A(KEYINPUT64), .B1(new_n201), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n202), .A2(KEYINPUT0), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT0), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G128), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT64), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n221), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n252), .B1(new_n254), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n251), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n196), .A2(KEYINPUT4), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n247), .A2(G101), .A3(new_n250), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT80), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n263), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND4_X1  g080(.A1(new_n247), .A2(KEYINPUT80), .A3(G101), .A4(new_n250), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n262), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  XOR2_X1   g082(.A(KEYINPUT82), .B(KEYINPUT10), .Z(new_n269));
  NAND2_X1  g083(.A1(new_n204), .A2(new_n205), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n270), .A2(G128), .A3(new_n209), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n213), .B1(new_n271), .B2(new_n221), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n269), .B1(new_n272), .B2(new_n216), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n215), .B1(new_n218), .B2(new_n222), .ZN(new_n274));
  AND3_X1   g088(.A1(new_n196), .A2(new_n199), .A3(KEYINPUT10), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  NOR3_X1   g091(.A1(new_n268), .A2(new_n277), .A3(new_n235), .ZN(new_n278));
  XNOR2_X1  g092(.A(G110), .B(G140), .ZN(new_n279));
  INV_X1    g093(.A(G953), .ZN(new_n280));
  AND2_X1   g094(.A1(new_n280), .A2(G227), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n279), .B(new_n281), .ZN(new_n282));
  OAI21_X1  g096(.A(KEYINPUT84), .B1(new_n278), .B2(new_n282), .ZN(new_n283));
  AOI22_X1  g097(.A1(new_n214), .A2(new_n269), .B1(new_n274), .B2(new_n275), .ZN(new_n284));
  AND2_X1   g098(.A1(new_n266), .A2(new_n267), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n236), .B(new_n284), .C1(new_n285), .C2(new_n262), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT84), .ZN(new_n287));
  INV_X1    g101(.A(new_n282), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n245), .A2(new_n283), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(KEYINPUT85), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT85), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n245), .A2(new_n283), .A3(new_n292), .A4(new_n289), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n235), .B1(new_n268), .B2(new_n277), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n288), .B1(new_n286), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n291), .A2(new_n293), .A3(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G469), .ZN(new_n298));
  INV_X1    g112(.A(G902), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n286), .A2(new_n288), .A3(new_n294), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n242), .A2(new_n243), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n302), .A2(new_n278), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n301), .B1(new_n303), .B2(new_n288), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n304), .A2(new_n298), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n298), .A2(new_n299), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n300), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g122(.A(KEYINPUT9), .B(G234), .ZN(new_n309));
  OAI21_X1  g123(.A(G221), .B1(new_n309), .B2(G902), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(G214), .B1(G237), .B2(G902), .ZN(new_n312));
  XNOR2_X1  g126(.A(new_n312), .B(KEYINPUT86), .ZN(new_n313));
  XOR2_X1   g127(.A(G116), .B(G119), .Z(new_n314));
  XNOR2_X1  g128(.A(KEYINPUT2), .B(G113), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT87), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT5), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n314), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G119), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n318), .A2(new_n320), .A3(G116), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G113), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n317), .B1(new_n319), .B2(new_n322), .ZN(new_n323));
  XNOR2_X1  g137(.A(G116), .B(G119), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n322), .B1(KEYINPUT5), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(KEYINPUT87), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n316), .B1(new_n323), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(new_n200), .ZN(new_n328));
  XNOR2_X1  g142(.A(G110), .B(G122), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n314), .B(new_n315), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n251), .A2(new_n330), .ZN(new_n331));
  OAI211_X1 g145(.A(new_n328), .B(new_n329), .C1(new_n285), .C2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n329), .ZN(new_n333));
  AND2_X1   g147(.A1(new_n333), .A2(KEYINPUT88), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n331), .B1(new_n266), .B2(new_n267), .ZN(new_n335));
  AOI211_X1 g149(.A(new_n316), .B(new_n216), .C1(new_n323), .C2(new_n326), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n334), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n332), .A2(new_n337), .A3(KEYINPUT6), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT6), .ZN(new_n339));
  OAI211_X1 g153(.A(new_n339), .B(new_n334), .C1(new_n335), .C2(new_n336), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n274), .A2(G125), .ZN(new_n341));
  INV_X1    g155(.A(G125), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n261), .A2(new_n342), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n280), .A2(G224), .ZN(new_n345));
  XNOR2_X1  g159(.A(new_n345), .B(KEYINPUT89), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n344), .B(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n338), .A2(new_n340), .A3(new_n347), .ZN(new_n348));
  XNOR2_X1  g162(.A(new_n329), .B(KEYINPUT8), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n325), .A2(new_n316), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n349), .B1(new_n350), .B2(new_n216), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n351), .B1(new_n216), .B2(new_n327), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n345), .A2(KEYINPUT7), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n344), .A2(new_n353), .ZN(new_n354));
  OAI211_X1 g168(.A(KEYINPUT7), .B(new_n345), .C1(new_n341), .C2(new_n343), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n352), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(G902), .B1(new_n356), .B2(new_n332), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n348), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g172(.A(G210), .B1(G237), .B2(G902), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(KEYINPUT90), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n358), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n348), .A2(new_n357), .A3(new_n361), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n313), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT97), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT20), .ZN(new_n367));
  XNOR2_X1  g181(.A(G113), .B(G122), .ZN(new_n368));
  XNOR2_X1  g182(.A(new_n368), .B(new_n189), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT16), .ZN(new_n371));
  INV_X1    g185(.A(G140), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n371), .A2(new_n372), .A3(G125), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(G125), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n342), .A2(G140), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  OAI211_X1 g190(.A(G146), .B(new_n373), .C1(new_n376), .C2(new_n371), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT77), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n374), .A2(new_n375), .A3(KEYINPUT77), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT19), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n376), .A2(KEYINPUT19), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n377), .B1(new_n384), .B2(G146), .ZN(new_n385));
  INV_X1    g199(.A(new_n233), .ZN(new_n386));
  INV_X1    g200(.A(G237), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(KEYINPUT70), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT70), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(G237), .ZN(new_n390));
  AOI21_X1  g204(.A(G953), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  XNOR2_X1  g205(.A(KEYINPUT91), .B(G143), .ZN(new_n392));
  AND3_X1   g206(.A1(new_n391), .A2(G214), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(KEYINPUT91), .A2(G143), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n395), .B1(new_n391), .B2(G214), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n386), .B1(new_n393), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n391), .A2(G214), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(new_n394), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n391), .A2(G214), .A3(new_n392), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n399), .A2(new_n233), .A3(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n385), .B1(new_n397), .B2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT18), .ZN(new_n403));
  INV_X1    g217(.A(G131), .ZN(new_n404));
  NOR3_X1   g218(.A1(new_n403), .A2(new_n404), .A3(KEYINPUT92), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n406), .B1(new_n393), .B2(new_n396), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n399), .A2(new_n405), .A3(new_n400), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n379), .A2(new_n380), .A3(new_n207), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n376), .A2(G146), .ZN(new_n410));
  AOI22_X1  g224(.A1(new_n407), .A2(new_n408), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n370), .B1(new_n402), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n373), .B1(new_n376), .B2(new_n371), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(new_n207), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(new_n377), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n233), .B1(new_n399), .B2(new_n400), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n415), .B1(new_n416), .B2(KEYINPUT17), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT17), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n397), .A2(new_n401), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n407), .A2(new_n408), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n409), .A2(new_n410), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n420), .A2(new_n369), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n412), .A2(new_n424), .ZN(new_n425));
  NOR2_X1   g239(.A1(G475), .A2(G902), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n367), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n426), .ZN(new_n428));
  AOI211_X1 g242(.A(KEYINPUT20), .B(new_n428), .C1(new_n412), .C2(new_n424), .ZN(new_n429));
  INV_X1    g243(.A(G475), .ZN(new_n430));
  AND3_X1   g244(.A1(new_n397), .A2(new_n401), .A3(new_n418), .ZN(new_n431));
  OAI211_X1 g245(.A(new_n414), .B(new_n377), .C1(new_n397), .C2(new_n418), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n423), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n370), .ZN(new_n434));
  AOI21_X1  g248(.A(G902), .B1(new_n434), .B2(new_n424), .ZN(new_n435));
  OAI22_X1  g249(.A1(new_n427), .A2(new_n429), .B1(new_n430), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(G234), .A2(G237), .ZN(new_n438));
  AND3_X1   g252(.A1(new_n438), .A2(G952), .A3(new_n280), .ZN(new_n439));
  XOR2_X1   g253(.A(KEYINPUT21), .B(G898), .Z(new_n440));
  XNOR2_X1  g254(.A(new_n440), .B(KEYINPUT96), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n438), .A2(G902), .A3(G953), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n443), .B(KEYINPUT95), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n439), .B1(new_n442), .B2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n203), .A2(G128), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n202), .A2(G143), .ZN(new_n449));
  AND3_X1   g263(.A1(new_n448), .A2(new_n449), .A3(new_n226), .ZN(new_n450));
  XOR2_X1   g264(.A(G116), .B(G122), .Z(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(G107), .ZN(new_n452));
  XNOR2_X1  g266(.A(G116), .B(G122), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(new_n192), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n450), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT13), .ZN(new_n456));
  OAI21_X1  g270(.A(KEYINPUT93), .B1(new_n448), .B2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT93), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n458), .A2(new_n203), .A3(KEYINPUT13), .A4(G128), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n448), .A2(new_n456), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n457), .A2(new_n459), .A3(new_n449), .A4(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(G134), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n455), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(G116), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n464), .A2(KEYINPUT14), .A3(G122), .ZN(new_n465));
  OAI211_X1 g279(.A(G107), .B(new_n465), .C1(new_n451), .C2(KEYINPUT14), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n226), .B1(new_n448), .B2(new_n449), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n466), .B(new_n454), .C1(new_n450), .C2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(G217), .ZN(new_n469));
  NOR3_X1   g283(.A1(new_n309), .A2(new_n469), .A3(G953), .ZN(new_n470));
  AND3_X1   g284(.A1(new_n463), .A2(new_n468), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n470), .B1(new_n463), .B2(new_n468), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n299), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(G478), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n474), .A2(KEYINPUT15), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  OAI221_X1 g290(.A(new_n299), .B1(KEYINPUT15), .B2(new_n474), .C1(new_n471), .C2(new_n472), .ZN(new_n477));
  AND3_X1   g291(.A1(new_n476), .A2(KEYINPUT94), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(KEYINPUT94), .B1(new_n476), .B2(new_n477), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n447), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n366), .B1(new_n437), .B2(new_n481), .ZN(new_n482));
  NOR3_X1   g296(.A1(new_n436), .A2(new_n480), .A3(KEYINPUT97), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n365), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n187), .B1(new_n311), .B2(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n469), .B1(G234), .B2(new_n299), .ZN(new_n486));
  OAI21_X1  g300(.A(KEYINPUT23), .B1(new_n202), .B2(G119), .ZN(new_n487));
  OAI21_X1  g301(.A(KEYINPUT74), .B1(new_n320), .B2(G128), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n487), .B(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(G110), .ZN(new_n490));
  OR3_X1    g304(.A1(new_n489), .A2(KEYINPUT75), .A3(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(KEYINPUT75), .B1(new_n489), .B2(new_n490), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  XOR2_X1   g307(.A(G119), .B(G128), .Z(new_n494));
  XNOR2_X1  g308(.A(KEYINPUT24), .B(G110), .ZN(new_n495));
  OR2_X1    g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n493), .A2(new_n496), .A3(new_n415), .ZN(new_n497));
  XNOR2_X1  g311(.A(KEYINPUT76), .B(G110), .ZN(new_n498));
  AOI22_X1  g312(.A1(new_n489), .A2(new_n498), .B1(new_n494), .B2(new_n495), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n409), .A2(new_n377), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n497), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n280), .A2(G221), .A3(G234), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n504), .B(KEYINPUT22), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n505), .B(G137), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n503), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n497), .A2(new_n502), .A3(new_n506), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n508), .A2(new_n299), .A3(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT78), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT25), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  AND2_X1   g327(.A1(new_n510), .A2(new_n512), .ZN(new_n514));
  OAI21_X1  g328(.A(KEYINPUT78), .B1(new_n510), .B2(new_n512), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n486), .B(new_n513), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n486), .A2(G902), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n508), .A2(new_n509), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n228), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n226), .A2(G137), .ZN(new_n521));
  OAI21_X1  g335(.A(G131), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n234), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(KEYINPUT68), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT68), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n234), .A2(new_n525), .A3(new_n522), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n274), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n261), .A2(new_n235), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n527), .A2(KEYINPUT30), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(KEYINPUT69), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT69), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n527), .A2(new_n531), .A3(KEYINPUT30), .A4(new_n528), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n523), .ZN(new_n534));
  AOI22_X1  g348(.A1(new_n274), .A2(new_n534), .B1(new_n261), .B2(new_n235), .ZN(new_n535));
  OAI21_X1  g349(.A(KEYINPUT67), .B1(new_n535), .B2(KEYINPUT30), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT67), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT30), .ZN(new_n538));
  AND2_X1   g352(.A1(new_n261), .A2(new_n235), .ZN(new_n539));
  OAI21_X1  g353(.A(KEYINPUT66), .B1(new_n217), .B2(new_n201), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n220), .A2(new_n219), .A3(new_n221), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n523), .B1(new_n542), .B2(new_n215), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n537), .B(new_n538), .C1(new_n539), .C2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n536), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n533), .A2(new_n330), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n391), .A2(G210), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(KEYINPUT27), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT26), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT27), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n391), .A2(new_n550), .A3(G210), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n548), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n549), .B1(new_n548), .B2(new_n551), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n194), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n554), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n556), .A2(G101), .A3(new_n552), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n330), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n527), .A2(new_n560), .A3(new_n528), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n546), .A2(new_n559), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(KEYINPUT31), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT28), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n330), .B1(new_n539), .B2(new_n543), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n527), .A2(KEYINPUT28), .A3(new_n560), .A4(new_n528), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(new_n558), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT31), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n546), .A2(new_n570), .A3(new_n559), .A4(new_n561), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n563), .A2(new_n569), .A3(new_n571), .ZN(new_n572));
  NOR2_X1   g386(.A1(G472), .A2(G902), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n573), .B(KEYINPUT71), .ZN(new_n574));
  AND3_X1   g388(.A1(new_n572), .A2(KEYINPUT32), .A3(new_n574), .ZN(new_n575));
  XOR2_X1   g389(.A(KEYINPUT72), .B(KEYINPUT32), .Z(new_n576));
  AOI21_X1  g390(.A(new_n576), .B1(new_n572), .B2(new_n574), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT29), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n579), .B1(new_n568), .B2(new_n558), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n546), .A2(new_n561), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n580), .B1(new_n581), .B2(new_n558), .ZN(new_n582));
  AND2_X1   g396(.A1(new_n565), .A2(new_n567), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n527), .A2(new_n528), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n330), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n583), .A2(KEYINPUT29), .A3(new_n559), .A4(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(new_n299), .ZN(new_n587));
  OAI21_X1  g401(.A(G472), .B1(new_n582), .B2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT73), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n583), .A2(new_n559), .A3(new_n566), .ZN(new_n591));
  INV_X1    g405(.A(new_n561), .ZN(new_n592));
  AOI22_X1  g406(.A1(new_n530), .A2(new_n532), .B1(new_n536), .B2(new_n544), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n592), .B1(new_n593), .B2(new_n330), .ZN(new_n594));
  OAI211_X1 g408(.A(new_n579), .B(new_n591), .C1(new_n594), .C2(new_n559), .ZN(new_n595));
  AND2_X1   g409(.A1(new_n586), .A2(new_n299), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n597), .A2(KEYINPUT73), .A3(G472), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n590), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n519), .B1(new_n578), .B2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n310), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n601), .B1(new_n300), .B2(new_n307), .ZN(new_n602));
  INV_X1    g416(.A(new_n483), .ZN(new_n603));
  OAI21_X1  g417(.A(KEYINPUT97), .B1(new_n436), .B2(new_n480), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n602), .A2(new_n605), .A3(KEYINPUT98), .A4(new_n365), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n485), .A2(new_n600), .A3(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(G101), .ZN(G3));
  NAND2_X1  g422(.A1(new_n572), .A2(new_n299), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(G472), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n572), .A2(new_n574), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NOR3_X1   g426(.A1(new_n311), .A2(new_n612), .A3(new_n519), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n313), .B1(new_n358), .B2(new_n359), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n348), .A2(new_n357), .A3(new_n360), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n614), .A2(new_n447), .A3(new_n615), .ZN(new_n616));
  OR2_X1    g430(.A1(new_n471), .A2(new_n472), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT33), .ZN(new_n618));
  OR2_X1    g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n617), .A2(new_n618), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n619), .A2(G478), .A3(new_n299), .A4(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n473), .A2(new_n474), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n436), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n616), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n613), .A2(new_n625), .ZN(new_n626));
  XOR2_X1   g440(.A(KEYINPUT34), .B(G104), .Z(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G6));
  INV_X1    g442(.A(KEYINPUT99), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n629), .B1(new_n435), .B2(new_n430), .ZN(new_n630));
  AND3_X1   g444(.A1(new_n420), .A2(new_n369), .A3(new_n423), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n369), .B1(new_n420), .B2(new_n423), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n299), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n633), .A2(KEYINPUT99), .A3(G475), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n630), .A2(new_n634), .ZN(new_n635));
  AND2_X1   g449(.A1(new_n412), .A2(new_n424), .ZN(new_n636));
  OAI21_X1  g450(.A(KEYINPUT20), .B1(new_n636), .B2(new_n428), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n425), .A2(new_n367), .A3(new_n426), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n478), .A2(new_n479), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n635), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n616), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n613), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT35), .B(G107), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G9));
  INV_X1    g459(.A(KEYINPUT100), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n507), .A2(KEYINPUT36), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n503), .B(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n517), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n516), .A2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n646), .B1(new_n612), .B2(new_n651), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n610), .A2(KEYINPUT100), .A3(new_n611), .A4(new_n650), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n485), .A2(new_n606), .A3(new_n652), .A4(new_n653), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT37), .B(G110), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G12));
  INV_X1    g470(.A(G900), .ZN(new_n657));
  AOI21_X1  g471(.A(KEYINPUT101), .B1(new_n445), .B2(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n658), .A2(new_n439), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n445), .A2(KEYINPUT101), .A3(new_n657), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n635), .A2(new_n639), .A3(new_n640), .A4(new_n661), .ZN(new_n662));
  AOI211_X1 g476(.A(new_n601), .B(new_n662), .C1(new_n300), .C2(new_n307), .ZN(new_n663));
  INV_X1    g477(.A(new_n576), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n611), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n572), .A2(KEYINPUT32), .A3(new_n574), .ZN(new_n666));
  AOI21_X1  g480(.A(KEYINPUT73), .B1(new_n597), .B2(G472), .ZN(new_n667));
  INV_X1    g481(.A(G472), .ZN(new_n668));
  AOI211_X1 g482(.A(new_n589), .B(new_n668), .C1(new_n595), .C2(new_n596), .ZN(new_n669));
  OAI211_X1 g483(.A(new_n665), .B(new_n666), .C1(new_n667), .C2(new_n669), .ZN(new_n670));
  AND2_X1   g484(.A1(new_n614), .A2(new_n615), .ZN(new_n671));
  AND2_X1   g485(.A1(new_n650), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n663), .A2(new_n670), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G128), .ZN(G30));
  XOR2_X1   g488(.A(new_n661), .B(KEYINPUT106), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(KEYINPUT39), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n602), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(KEYINPUT40), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n363), .A2(new_n364), .ZN(new_n679));
  XOR2_X1   g493(.A(new_n679), .B(KEYINPUT102), .Z(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(KEYINPUT38), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n585), .A2(new_n561), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n558), .ZN(new_n683));
  XOR2_X1   g497(.A(new_n683), .B(KEYINPUT103), .Z(new_n684));
  INV_X1    g498(.A(new_n562), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n299), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(G472), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n665), .A2(new_n687), .A3(new_n666), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n436), .A2(new_n640), .ZN(new_n689));
  NOR3_X1   g503(.A1(new_n650), .A2(new_n689), .A3(new_n313), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(KEYINPUT104), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n681), .A2(new_n688), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(KEYINPUT105), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT105), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n681), .A2(new_n694), .A3(new_n688), .A4(new_n691), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n678), .B1(new_n693), .B2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(new_n203), .ZN(G45));
  NAND3_X1  g511(.A1(new_n436), .A2(new_n623), .A3(new_n661), .ZN(new_n698));
  AOI211_X1 g512(.A(new_n601), .B(new_n698), .C1(new_n300), .C2(new_n307), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n670), .A2(new_n699), .A3(new_n672), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(KEYINPUT107), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G146), .ZN(G48));
  AOI21_X1  g516(.A(new_n295), .B1(new_n290), .B2(KEYINPUT85), .ZN(new_n703));
  AOI211_X1 g517(.A(G469), .B(G902), .C1(new_n703), .C2(new_n293), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n298), .B1(new_n297), .B2(new_n299), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n704), .A2(new_n705), .A3(new_n601), .ZN(new_n706));
  INV_X1    g520(.A(new_n519), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n670), .A2(new_n706), .A3(new_n707), .A4(new_n625), .ZN(new_n708));
  XNOR2_X1  g522(.A(KEYINPUT41), .B(G113), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n708), .B(new_n709), .ZN(G15));
  NAND4_X1  g524(.A1(new_n670), .A2(new_n706), .A3(new_n707), .A4(new_n642), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G116), .ZN(G18));
  NAND2_X1  g526(.A1(new_n297), .A2(new_n299), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(G469), .ZN(new_n714));
  AND4_X1   g528(.A1(new_n310), .A2(new_n714), .A3(new_n300), .A4(new_n671), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n715), .A2(new_n670), .A3(new_n605), .A4(new_n650), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G119), .ZN(G21));
  AND2_X1   g531(.A1(new_n583), .A2(new_n585), .ZN(new_n718));
  OAI211_X1 g532(.A(new_n563), .B(new_n571), .C1(new_n559), .C2(new_n718), .ZN(new_n719));
  AND2_X1   g533(.A1(new_n719), .A2(new_n574), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n668), .B1(new_n572), .B2(new_n299), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n720), .A2(new_n519), .A3(new_n721), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n616), .A2(new_n689), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n722), .A2(new_n706), .A3(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G122), .ZN(G24));
  NOR3_X1   g539(.A1(new_n720), .A2(new_n721), .A3(new_n698), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n726), .A2(new_n706), .A3(new_n671), .A4(new_n650), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G125), .ZN(G27));
  OAI21_X1  g542(.A(KEYINPUT108), .B1(new_n303), .B2(new_n288), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT108), .ZN(new_n730));
  OAI211_X1 g544(.A(new_n730), .B(new_n282), .C1(new_n302), .C2(new_n278), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n729), .A2(new_n301), .A3(new_n731), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n298), .B1(new_n732), .B2(new_n299), .ZN(new_n733));
  AOI21_X1  g547(.A(G902), .B1(new_n703), .B2(new_n293), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n733), .B1(new_n734), .B2(new_n298), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n601), .A2(new_n313), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n363), .A2(new_n364), .A3(new_n736), .ZN(new_n737));
  OAI21_X1  g551(.A(KEYINPUT109), .B1(new_n735), .B2(new_n737), .ZN(new_n738));
  AND3_X1   g552(.A1(new_n729), .A2(new_n301), .A3(new_n731), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n306), .B1(new_n739), .B2(G469), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n300), .A2(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(new_n737), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT109), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n741), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n738), .A2(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(new_n698), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n745), .A2(new_n600), .A3(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT42), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  AOI21_X1  g563(.A(KEYINPUT32), .B1(new_n572), .B2(new_n574), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  AND3_X1   g565(.A1(new_n599), .A2(new_n666), .A3(new_n751), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n752), .A2(new_n519), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n698), .A2(new_n748), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n753), .A2(new_n745), .A3(new_n754), .ZN(new_n755));
  AND2_X1   g569(.A1(new_n749), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(new_n404), .ZN(G33));
  INV_X1    g571(.A(new_n662), .ZN(new_n758));
  AND3_X1   g572(.A1(new_n745), .A2(new_n600), .A3(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(new_n226), .ZN(G36));
  NAND2_X1  g574(.A1(new_n739), .A2(KEYINPUT45), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT45), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n298), .B1(new_n304), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n764), .B1(new_n298), .B2(new_n299), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT46), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n704), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n767), .B1(new_n766), .B2(new_n765), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n768), .A2(new_n310), .A3(new_n676), .ZN(new_n769));
  INV_X1    g583(.A(new_n679), .ZN(new_n770));
  INV_X1    g584(.A(new_n313), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n437), .A2(KEYINPUT43), .A3(new_n623), .ZN(new_n774));
  XOR2_X1   g588(.A(new_n774), .B(KEYINPUT111), .Z(new_n775));
  INV_X1    g589(.A(KEYINPUT43), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n623), .B(KEYINPUT110), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n776), .B1(new_n777), .B2(new_n436), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n651), .B1(new_n775), .B2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT44), .ZN(new_n780));
  AND3_X1   g594(.A1(new_n779), .A2(new_n780), .A3(new_n612), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n780), .B1(new_n779), .B2(new_n612), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n769), .B(new_n773), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G137), .ZN(G39));
  NAND2_X1  g598(.A1(new_n768), .A2(new_n310), .ZN(new_n785));
  OR2_X1    g599(.A1(new_n785), .A2(KEYINPUT47), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(KEYINPUT47), .ZN(new_n787));
  NOR4_X1   g601(.A1(new_n670), .A2(new_n707), .A3(new_n698), .A4(new_n772), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n786), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G140), .ZN(G42));
  INV_X1    g604(.A(new_n681), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n707), .A2(new_n736), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT112), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n437), .B(new_n623), .C1(new_n792), .C2(new_n793), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n794), .B1(new_n793), .B2(new_n792), .ZN(new_n795));
  INV_X1    g609(.A(new_n688), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n704), .A2(new_n705), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(KEYINPUT49), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n791), .A2(new_n795), .A3(new_n796), .A4(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(KEYINPUT113), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT51), .ZN(new_n801));
  AOI22_X1  g615(.A1(new_n787), .A2(new_n786), .B1(new_n601), .B2(new_n797), .ZN(new_n802));
  INV_X1    g616(.A(new_n439), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n803), .B1(new_n775), .B2(new_n778), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n804), .A2(new_n722), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(new_n773), .ZN(new_n806));
  OR2_X1    g620(.A1(new_n802), .A2(new_n806), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n704), .A2(new_n705), .A3(new_n737), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n804), .A2(new_n808), .ZN(new_n809));
  NOR4_X1   g623(.A1(new_n809), .A2(new_n721), .A3(new_n651), .A4(new_n720), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n796), .A2(new_n707), .A3(new_n439), .A4(new_n808), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n811), .A2(new_n436), .A3(new_n623), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n807), .A2(new_n813), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n805), .A2(new_n313), .A3(new_n791), .A4(new_n706), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(KEYINPUT50), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n801), .B1(new_n814), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n280), .A2(G952), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n818), .B1(new_n805), .B2(new_n715), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT48), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(KEYINPUT119), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n753), .B1(KEYINPUT119), .B2(new_n820), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n809), .A2(new_n822), .ZN(new_n823));
  OAI221_X1 g637(.A(new_n819), .B1(new_n624), .B2(new_n811), .C1(new_n821), .C2(new_n823), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n824), .B1(new_n821), .B2(new_n823), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n813), .B(KEYINPUT118), .ZN(new_n826));
  INV_X1    g640(.A(new_n816), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n827), .A2(KEYINPUT51), .A3(new_n807), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n817), .B(new_n825), .C1(new_n826), .C2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT114), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n612), .A2(new_n519), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n679), .A2(new_n771), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n832), .A2(new_n624), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n831), .A2(new_n602), .A3(new_n447), .A4(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n830), .B1(new_n607), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n476), .A2(new_n477), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n437), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n832), .A2(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n831), .A2(new_n602), .A3(new_n447), .A4(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n654), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n835), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n759), .B1(new_n749), .B2(new_n755), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n716), .A2(new_n708), .A3(new_n711), .A4(new_n724), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n743), .B1(new_n741), .B2(new_n742), .ZN(new_n844));
  AOI211_X1 g658(.A(KEYINPUT109), .B(new_n737), .C1(new_n300), .C2(new_n740), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n726), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n635), .A2(new_n639), .ZN(new_n847));
  INV_X1    g661(.A(new_n661), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n847), .A2(new_n836), .A3(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n670), .A2(new_n602), .A3(new_n773), .A4(new_n849), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n651), .B1(new_n846), .B2(new_n850), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n843), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n607), .A2(new_n830), .A3(new_n834), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n841), .A2(new_n842), .A3(new_n852), .A4(new_n853), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n671), .A2(new_n436), .A3(new_n640), .ZN(new_n855));
  AND4_X1   g669(.A1(new_n516), .A2(new_n310), .A3(new_n649), .A4(new_n661), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n855), .A2(new_n688), .A3(new_n741), .A4(new_n856), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n727), .A2(new_n673), .A3(new_n700), .A4(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT52), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT115), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n670), .B(new_n672), .C1(new_n663), .C2(new_n699), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n862), .A2(KEYINPUT52), .A3(new_n727), .A4(new_n857), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n860), .A2(new_n861), .A3(new_n863), .ZN(new_n864));
  OR2_X1    g678(.A1(new_n863), .A2(new_n861), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n854), .A2(new_n866), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n607), .A2(new_n830), .A3(new_n834), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n868), .A2(new_n835), .A3(new_n840), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n860), .A2(new_n863), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n869), .A2(new_n842), .A3(new_n852), .A4(new_n870), .ZN(new_n871));
  XOR2_X1   g685(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n872));
  OAI22_X1  g686(.A1(new_n867), .A2(KEYINPUT53), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(KEYINPUT54), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n842), .A2(new_n852), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n607), .A2(new_n834), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(KEYINPUT114), .ZN(new_n877));
  AND2_X1   g691(.A1(new_n654), .A2(new_n839), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n877), .A2(new_n878), .A3(new_n853), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n875), .A2(new_n879), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n864), .A2(new_n865), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n880), .A2(new_n881), .A3(KEYINPUT53), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n871), .A2(new_n872), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  XOR2_X1   g698(.A(KEYINPUT117), .B(KEYINPUT54), .Z(new_n885));
  INV_X1    g699(.A(new_n885), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n874), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n829), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(G952), .A2(G953), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n800), .B1(new_n888), .B2(new_n889), .ZN(G75));
  AOI22_X1  g704(.A1(new_n867), .A2(KEYINPUT53), .B1(new_n871), .B2(new_n872), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n891), .A2(new_n299), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(G210), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n338), .A2(new_n340), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n894), .B(new_n347), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(KEYINPUT55), .ZN(new_n896));
  XNOR2_X1  g710(.A(KEYINPUT120), .B(KEYINPUT56), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n893), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT56), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n896), .B1(new_n893), .B2(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n280), .A2(G952), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n898), .A2(new_n900), .A3(new_n901), .ZN(G51));
  XNOR2_X1  g716(.A(new_n891), .B(new_n886), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n306), .B(KEYINPUT57), .Z(new_n904));
  OAI21_X1  g718(.A(new_n297), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n892), .A2(new_n761), .A3(new_n763), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n901), .B1(new_n905), .B2(new_n906), .ZN(G54));
  NAND3_X1  g721(.A1(new_n892), .A2(KEYINPUT58), .A3(G475), .ZN(new_n908));
  AND3_X1   g722(.A1(new_n908), .A2(KEYINPUT121), .A3(new_n636), .ZN(new_n909));
  INV_X1    g723(.A(new_n901), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n910), .B1(new_n908), .B2(new_n636), .ZN(new_n911));
  AOI21_X1  g725(.A(KEYINPUT121), .B1(new_n908), .B2(new_n636), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n909), .A2(new_n911), .A3(new_n912), .ZN(G60));
  AND2_X1   g727(.A1(new_n619), .A2(new_n620), .ZN(new_n914));
  NAND2_X1  g728(.A1(G478), .A2(G902), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(KEYINPUT59), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n910), .B1(new_n903), .B2(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n914), .B1(new_n887), .B2(new_n916), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n918), .A2(new_n919), .ZN(G63));
  NAND2_X1  g734(.A1(new_n508), .A2(new_n509), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT122), .ZN(new_n922));
  NAND2_X1  g736(.A1(G217), .A2(G902), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT60), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n922), .B1(new_n891), .B2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(new_n924), .ZN(new_n926));
  INV_X1    g740(.A(new_n872), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n927), .B1(new_n880), .B2(new_n870), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT53), .ZN(new_n929));
  NOR3_X1   g743(.A1(new_n854), .A2(new_n866), .A3(new_n929), .ZN(new_n930));
  OAI211_X1 g744(.A(new_n648), .B(new_n926), .C1(new_n928), .C2(new_n930), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n925), .A2(KEYINPUT61), .A3(new_n910), .A4(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(KEYINPUT124), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n926), .B1(new_n928), .B2(new_n930), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n901), .B1(new_n934), .B2(new_n922), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT124), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n935), .A2(new_n936), .A3(KEYINPUT61), .A4(new_n931), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n933), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n935), .A2(new_n931), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT61), .ZN(new_n940));
  AOI21_X1  g754(.A(KEYINPUT123), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n924), .B1(new_n882), .B2(new_n883), .ZN(new_n942));
  INV_X1    g756(.A(new_n922), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n910), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(new_n931), .ZN(new_n945));
  OAI211_X1 g759(.A(KEYINPUT123), .B(new_n940), .C1(new_n944), .C2(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(new_n946), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n938), .B1(new_n941), .B2(new_n947), .ZN(G66));
  INV_X1    g762(.A(G224), .ZN(new_n949));
  OAI21_X1  g763(.A(G953), .B1(new_n442), .B2(new_n949), .ZN(new_n950));
  OR2_X1    g764(.A1(new_n879), .A2(new_n843), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT125), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n950), .B1(new_n952), .B2(G953), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n894), .B1(G898), .B2(new_n280), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n953), .B(new_n954), .ZN(G69));
  NAND2_X1  g769(.A1(new_n862), .A2(new_n727), .ZN(new_n956));
  INV_X1    g770(.A(new_n956), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n769), .A2(new_n753), .A3(new_n855), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n789), .A2(new_n783), .A3(new_n957), .A4(new_n958), .ZN(new_n959));
  NOR3_X1   g773(.A1(new_n959), .A2(new_n756), .A3(new_n759), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(new_n280), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n593), .B(new_n384), .Z(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n963), .B1(G900), .B2(G953), .ZN(new_n964));
  AOI21_X1  g778(.A(KEYINPUT127), .B1(new_n961), .B2(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT126), .ZN(new_n966));
  INV_X1    g780(.A(new_n696), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT62), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n967), .A2(new_n968), .A3(new_n957), .ZN(new_n969));
  OAI21_X1  g783(.A(KEYINPUT62), .B1(new_n696), .B2(new_n956), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n772), .B1(new_n624), .B2(new_n837), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n600), .A2(new_n602), .A3(new_n676), .A4(new_n971), .ZN(new_n972));
  AND3_X1   g786(.A1(new_n789), .A2(new_n783), .A3(new_n972), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n969), .A2(new_n970), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n974), .A2(new_n280), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n966), .B1(new_n975), .B2(new_n963), .ZN(new_n976));
  AOI211_X1 g790(.A(KEYINPUT126), .B(new_n962), .C1(new_n974), .C2(new_n280), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n965), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n280), .B1(G227), .B2(G900), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(new_n979), .ZN(new_n981));
  OAI211_X1 g795(.A(new_n981), .B(new_n965), .C1(new_n976), .C2(new_n977), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n980), .A2(new_n982), .ZN(G72));
  NAND2_X1  g797(.A1(G472), .A2(G902), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n984), .B(KEYINPUT63), .Z(new_n985));
  XOR2_X1   g799(.A(new_n951), .B(KEYINPUT125), .Z(new_n986));
  OAI21_X1  g800(.A(new_n985), .B1(new_n986), .B2(new_n974), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n987), .A2(new_n559), .A3(new_n581), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n594), .A2(new_n559), .ZN(new_n989));
  OAI211_X1 g803(.A(new_n873), .B(new_n985), .C1(new_n989), .C2(new_n685), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n988), .A2(new_n910), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n952), .A2(new_n960), .ZN(new_n992));
  AOI211_X1 g806(.A(new_n559), .B(new_n581), .C1(new_n992), .C2(new_n985), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n991), .A2(new_n993), .ZN(G57));
endmodule


