//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 1 0 0 1 1 1 0 1 1 1 0 0 1 0 0 0 1 1 1 1 0 0 0 1 1 1 1 0 1 0 0 0 0 1 0 0 1 0 0 0 0 1 1 1 0 0 0 0 1 0 0 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:30 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n559, new_n560, new_n561,
    new_n562, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n572, new_n574, new_n575, new_n576, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n590,
    new_n591, new_n592, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n621, new_n622, new_n625,
    new_n627, new_n628, new_n629, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1124,
    new_n1125;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT64), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT65), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n447), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT66), .Z(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT67), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT2), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n454), .A2(new_n456), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(new_n456), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n453), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT68), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT68), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g043(.A(KEYINPUT3), .B(G2104), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n468), .A2(new_n469), .A3(G137), .ZN(new_n470));
  AND3_X1   g045(.A1(new_n464), .A2(KEYINPUT70), .A3(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(KEYINPUT70), .B1(new_n464), .B2(G2104), .ZN(new_n472));
  OAI21_X1  g047(.A(G101), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(KEYINPUT71), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT71), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n470), .A2(new_n473), .A3(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n468), .ZN(new_n478));
  INV_X1    g053(.A(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(KEYINPUT3), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT3), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G2104), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n480), .A2(new_n482), .A3(G125), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(KEYINPUT69), .ZN(new_n484));
  NAND2_X1  g059(.A1(G113), .A2(G2104), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT69), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n480), .A2(new_n482), .A3(new_n486), .A4(G125), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n484), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  AOI22_X1  g063(.A1(new_n475), .A2(new_n477), .B1(new_n478), .B2(new_n488), .ZN(new_n489));
  XNOR2_X1  g064(.A(new_n489), .B(KEYINPUT72), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G160));
  AND3_X1   g066(.A1(new_n469), .A2(new_n465), .A3(new_n467), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n469), .A2(new_n464), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  AOI22_X1  g069(.A1(G124), .A2(new_n492), .B1(new_n494), .B2(G136), .ZN(new_n495));
  OAI221_X1 g070(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n468), .C2(G112), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  XNOR2_X1  g072(.A(new_n497), .B(KEYINPUT73), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G162));
  NAND3_X1  g074(.A1(new_n468), .A2(new_n469), .A3(G138), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n501), .A2(KEYINPUT76), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n502), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n468), .A2(new_n469), .A3(new_n504), .A4(G138), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  OR2_X1    g081(.A1(KEYINPUT74), .A2(G114), .ZN(new_n507));
  NAND2_X1  g082(.A1(KEYINPUT74), .A2(G114), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n507), .A2(G2105), .A3(new_n508), .ZN(new_n509));
  OAI21_X1  g084(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND4_X1  g087(.A1(new_n480), .A2(new_n482), .A3(G126), .A4(G2105), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(KEYINPUT75), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT75), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n512), .A2(new_n516), .A3(new_n513), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n506), .A2(new_n515), .A3(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(G164));
  INV_X1    g094(.A(KEYINPUT78), .ZN(new_n520));
  INV_X1    g095(.A(G651), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n520), .B1(new_n521), .B2(KEYINPUT6), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT6), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n523), .A2(KEYINPUT78), .A3(G651), .ZN(new_n524));
  AND2_X1   g099(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(G543), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(KEYINPUT5), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT5), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G543), .ZN(new_n529));
  AND2_X1   g104(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  OAI21_X1  g105(.A(KEYINPUT77), .B1(new_n523), .B2(G651), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT77), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n532), .A2(new_n521), .A3(KEYINPUT6), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND4_X1  g109(.A1(new_n525), .A2(G88), .A3(new_n530), .A4(new_n534), .ZN(new_n535));
  NAND4_X1  g110(.A1(new_n525), .A2(G50), .A3(G543), .A4(new_n534), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT79), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n535), .A2(new_n536), .A3(KEYINPUT79), .ZN(new_n540));
  NAND2_X1  g115(.A1(G75), .A2(G543), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n527), .A2(new_n529), .ZN(new_n542));
  INV_X1    g117(.A(G62), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n539), .A2(new_n540), .B1(G651), .B2(new_n544), .ZN(G166));
  NAND3_X1  g120(.A1(new_n525), .A2(new_n530), .A3(new_n534), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(KEYINPUT80), .A2(G89), .ZN(new_n548));
  OR2_X1    g123(.A1(KEYINPUT80), .A2(G89), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n525), .A2(G543), .A3(new_n534), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G51), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n530), .A2(G63), .A3(G651), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n550), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NAND3_X1  g130(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n556));
  XOR2_X1   g131(.A(new_n556), .B(KEYINPUT7), .Z(new_n557));
  NOR2_X1   g132(.A1(new_n555), .A2(new_n557), .ZN(G168));
  NAND2_X1  g133(.A1(new_n547), .A2(G90), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n552), .A2(G52), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n530), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n561));
  OR2_X1    g136(.A1(new_n561), .A2(new_n521), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n559), .A2(new_n560), .A3(new_n562), .ZN(G301));
  INV_X1    g138(.A(G301), .ZN(G171));
  NAND2_X1  g139(.A1(new_n547), .A2(G81), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n552), .A2(G43), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n530), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n567));
  OR2_X1    g142(.A1(new_n567), .A2(new_n521), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n565), .A2(new_n566), .A3(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G860), .ZN(G153));
  AND3_X1   g146(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(G36), .ZN(G176));
  NAND2_X1  g148(.A1(G1), .A2(G3), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n574), .B(KEYINPUT8), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  XOR2_X1   g151(.A(new_n576), .B(KEYINPUT81), .Z(G188));
  NAND4_X1  g152(.A1(new_n525), .A2(G53), .A3(G543), .A4(new_n534), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT9), .ZN(new_n579));
  NAND2_X1  g154(.A1(G78), .A2(G543), .ZN(new_n580));
  INV_X1    g155(.A(G65), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n542), .B2(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n578), .A2(new_n579), .B1(G651), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n547), .A2(G91), .ZN(new_n584));
  AND3_X1   g159(.A1(new_n534), .A2(new_n522), .A3(new_n524), .ZN(new_n585));
  NAND4_X1  g160(.A1(new_n585), .A2(KEYINPUT9), .A3(G53), .A4(G543), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n583), .A2(new_n584), .A3(new_n586), .ZN(G299));
  INV_X1    g162(.A(G168), .ZN(G286));
  INV_X1    g163(.A(G166), .ZN(G303));
  NAND4_X1  g164(.A1(new_n525), .A2(G49), .A3(G543), .A4(new_n534), .ZN(new_n590));
  OAI21_X1  g165(.A(G651), .B1(new_n530), .B2(G74), .ZN(new_n591));
  INV_X1    g166(.A(G87), .ZN(new_n592));
  OAI211_X1 g167(.A(new_n590), .B(new_n591), .C1(new_n546), .C2(new_n592), .ZN(G288));
  NAND2_X1  g168(.A1(G73), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G61), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n542), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n596), .A2(G651), .ZN(new_n597));
  NAND4_X1  g172(.A1(new_n525), .A2(G48), .A3(G543), .A4(new_n534), .ZN(new_n598));
  NAND4_X1  g173(.A1(new_n525), .A2(G86), .A3(new_n530), .A4(new_n534), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(G305));
  NAND2_X1  g175(.A1(new_n547), .A2(G85), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n552), .A2(G47), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n530), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n603));
  OAI211_X1 g178(.A(new_n601), .B(new_n602), .C1(new_n521), .C2(new_n603), .ZN(G290));
  NAND2_X1  g179(.A1(G301), .A2(G868), .ZN(new_n605));
  INV_X1    g180(.A(G54), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n551), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n547), .A2(KEYINPUT10), .A3(G92), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT10), .ZN(new_n609));
  INV_X1    g184(.A(G92), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n546), .B2(new_n610), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n607), .B1(new_n608), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n530), .A2(G66), .ZN(new_n613));
  NAND2_X1  g188(.A1(G79), .A2(G543), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT82), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n521), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(new_n617));
  AND2_X1   g192(.A1(new_n612), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n605), .B1(new_n618), .B2(G868), .ZN(G284));
  OAI21_X1  g194(.A(new_n605), .B1(new_n618), .B2(G868), .ZN(G321));
  INV_X1    g195(.A(G868), .ZN(new_n621));
  NAND2_X1  g196(.A1(G299), .A2(new_n621), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(G168), .B2(new_n621), .ZN(G297));
  OAI21_X1  g198(.A(new_n622), .B1(G168), .B2(new_n621), .ZN(G280));
  INV_X1    g199(.A(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n618), .B1(new_n625), .B2(G860), .ZN(G148));
  NAND2_X1  g201(.A1(new_n569), .A2(new_n621), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n612), .A2(new_n617), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n628), .A2(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n627), .B1(new_n629), .B2(new_n621), .ZN(G323));
  XNOR2_X1  g205(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g206(.A1(new_n471), .A2(new_n472), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(new_n469), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(KEYINPUT12), .Z(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(KEYINPUT13), .Z(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT83), .B(G2100), .ZN(new_n636));
  INV_X1    g211(.A(KEYINPUT84), .ZN(new_n637));
  AND2_X1   g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g213(.A1(new_n636), .A2(new_n637), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n635), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  AOI22_X1  g215(.A1(G123), .A2(new_n492), .B1(new_n494), .B2(G135), .ZN(new_n641));
  OAI221_X1 g216(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n468), .C2(G111), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(G2096), .Z(new_n644));
  OAI211_X1 g219(.A(new_n640), .B(new_n644), .C1(new_n635), .C2(new_n638), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(KEYINPUT85), .Z(G156));
  XNOR2_X1  g221(.A(KEYINPUT15), .B(G2430), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2435), .ZN(new_n648));
  XOR2_X1   g223(.A(G2427), .B(G2438), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n650), .A2(KEYINPUT14), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2443), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2451), .B(G2454), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT86), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n652), .B(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(KEYINPUT16), .B(G2446), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G1341), .B(G1348), .Z(new_n658));
  AND2_X1   g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n657), .A2(new_n658), .ZN(new_n660));
  OAI21_X1  g235(.A(G14), .B1(new_n660), .B2(KEYINPUT87), .ZN(new_n661));
  AOI211_X1 g236(.A(new_n659), .B(new_n661), .C1(KEYINPUT87), .C2(new_n660), .ZN(G401));
  XOR2_X1   g237(.A(G2072), .B(G2078), .Z(new_n663));
  XOR2_X1   g238(.A(G2084), .B(G2090), .Z(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G2067), .B(G2678), .Z(new_n666));
  OR2_X1    g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g242(.A(new_n663), .B1(new_n667), .B2(KEYINPUT18), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(G2100), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n665), .A2(new_n666), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n667), .A2(new_n670), .A3(KEYINPUT17), .ZN(new_n671));
  INV_X1    g246(.A(KEYINPUT18), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n669), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT88), .B(G2096), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(G227));
  XNOR2_X1  g251(.A(G1971), .B(G1976), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT89), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n678), .B(KEYINPUT19), .Z(new_n679));
  XOR2_X1   g254(.A(G1956), .B(G2474), .Z(new_n680));
  XOR2_X1   g255(.A(G1961), .B(G1966), .Z(new_n681));
  AND2_X1   g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT20), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n680), .A2(new_n681), .ZN(new_n685));
  OR3_X1    g260(.A1(new_n679), .A2(new_n682), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n679), .A2(new_n685), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n684), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1991), .B(G1996), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1981), .B(G1986), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(G229));
  MUX2_X1   g269(.A(G24), .B(G290), .S(G16), .Z(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT91), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(G1986), .ZN(new_n697));
  MUX2_X1   g272(.A(G6), .B(G305), .S(G16), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT92), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT32), .B(G1981), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  MUX2_X1   g276(.A(G23), .B(G288), .S(G16), .Z(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT93), .B(KEYINPUT33), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(G1976), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n702), .B(new_n704), .ZN(new_n705));
  MUX2_X1   g280(.A(G22), .B(G303), .S(G16), .Z(new_n706));
  OR2_X1    g281(.A1(new_n706), .A2(G1971), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n706), .A2(G1971), .ZN(new_n708));
  NAND4_X1  g283(.A1(new_n701), .A2(new_n705), .A3(new_n707), .A4(new_n708), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n697), .B1(new_n709), .B2(KEYINPUT34), .ZN(new_n710));
  AOI22_X1  g285(.A1(G119), .A2(new_n492), .B1(new_n494), .B2(G131), .ZN(new_n711));
  OAI221_X1 g286(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n468), .C2(G107), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  MUX2_X1   g288(.A(G25), .B(new_n713), .S(G29), .Z(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT35), .B(G1991), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT90), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n714), .B(new_n716), .ZN(new_n717));
  OAI211_X1 g292(.A(new_n710), .B(new_n717), .C1(KEYINPUT34), .C2(new_n709), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT36), .ZN(new_n719));
  INV_X1    g294(.A(G29), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(G27), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G164), .B2(new_n720), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT100), .B(G2078), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  OR2_X1    g299(.A1(G29), .A2(G33), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(KEYINPUT25), .Z(new_n727));
  AOI22_X1  g302(.A1(new_n469), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n728), .A2(new_n468), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n494), .A2(G139), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n727), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n725), .B1(new_n731), .B2(new_n720), .ZN(new_n732));
  INV_X1    g307(.A(G2072), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT95), .ZN(new_n735));
  NOR2_X1   g310(.A1(G29), .A2(G32), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n632), .A2(G105), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT96), .ZN(new_n738));
  NAND3_X1  g313(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT26), .Z(new_n740));
  AOI22_X1  g315(.A1(G129), .A2(new_n492), .B1(new_n494), .B2(G141), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n738), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(new_n742), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n736), .B1(new_n743), .B2(G29), .ZN(new_n744));
  XOR2_X1   g319(.A(KEYINPUT27), .B(G1996), .Z(new_n745));
  NAND2_X1  g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n641), .A2(G29), .A3(new_n642), .ZN(new_n747));
  XNOR2_X1  g322(.A(KEYINPUT97), .B(KEYINPUT30), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(G28), .ZN(new_n749));
  OAI211_X1 g324(.A(new_n746), .B(new_n747), .C1(G29), .C2(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n744), .A2(new_n745), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n732), .A2(new_n733), .ZN(new_n752));
  XOR2_X1   g327(.A(KEYINPUT31), .B(G11), .Z(new_n753));
  NOR4_X1   g328(.A1(new_n750), .A2(new_n751), .A3(new_n752), .A4(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT28), .ZN(new_n755));
  INV_X1    g330(.A(G26), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n755), .B1(new_n756), .B2(G29), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n756), .A2(G29), .ZN(new_n758));
  AOI22_X1  g333(.A1(G128), .A2(new_n492), .B1(new_n494), .B2(G140), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n468), .A2(G116), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT94), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G104), .B2(G2105), .ZN(new_n762));
  OR3_X1    g337(.A1(new_n761), .A2(G104), .A3(G2105), .ZN(new_n763));
  NAND4_X1  g338(.A1(new_n760), .A2(G2104), .A3(new_n762), .A4(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n759), .A2(new_n764), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n758), .B1(new_n765), .B2(G29), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n757), .B1(new_n766), .B2(new_n755), .ZN(new_n767));
  OR2_X1    g342(.A1(new_n767), .A2(G2067), .ZN(new_n768));
  NOR2_X1   g343(.A1(G5), .A2(G16), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(G171), .B2(G16), .ZN(new_n770));
  AOI22_X1  g345(.A1(G2067), .A2(new_n767), .B1(new_n770), .B2(G1961), .ZN(new_n771));
  AND4_X1   g346(.A1(new_n735), .A2(new_n754), .A3(new_n768), .A4(new_n771), .ZN(new_n772));
  MUX2_X1   g347(.A(G19), .B(new_n569), .S(G16), .Z(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(G1341), .Z(new_n774));
  OR2_X1    g349(.A1(KEYINPUT24), .A2(G34), .ZN(new_n775));
  NAND2_X1  g350(.A1(KEYINPUT24), .A2(G34), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n775), .A2(new_n720), .A3(new_n776), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G160), .B2(new_n720), .ZN(new_n778));
  OR2_X1    g353(.A1(new_n778), .A2(G2084), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n779), .A2(KEYINPUT99), .ZN(new_n780));
  OR2_X1    g355(.A1(new_n779), .A2(KEYINPUT99), .ZN(new_n781));
  NAND4_X1  g356(.A1(new_n772), .A2(new_n774), .A3(new_n780), .A4(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(G168), .A2(G16), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G16), .B2(G21), .ZN(new_n784));
  INV_X1    g359(.A(G1966), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT98), .Z(new_n787));
  NOR2_X1   g362(.A1(G29), .A2(G35), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(G162), .B2(G29), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT29), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(G2090), .ZN(new_n791));
  NAND2_X1  g366(.A1(G299), .A2(G16), .ZN(new_n792));
  XNOR2_X1  g367(.A(KEYINPUT101), .B(KEYINPUT23), .ZN(new_n793));
  INV_X1    g368(.A(G20), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n794), .A2(G16), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n793), .B(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n792), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(G1956), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(G2084), .B2(new_n778), .ZN(new_n799));
  OR2_X1    g374(.A1(new_n770), .A2(G1961), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n784), .A2(new_n785), .ZN(new_n801));
  INV_X1    g376(.A(G4), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n802), .A2(G16), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(new_n628), .B2(G16), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(G1348), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n799), .A2(new_n800), .A3(new_n801), .A4(new_n805), .ZN(new_n806));
  NOR4_X1   g381(.A1(new_n782), .A2(new_n787), .A3(new_n791), .A4(new_n806), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n719), .A2(new_n724), .A3(new_n807), .ZN(G150));
  INV_X1    g383(.A(G150), .ZN(G311));
  NAND2_X1  g384(.A1(new_n547), .A2(G93), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n552), .A2(G55), .ZN(new_n811));
  AOI22_X1  g386(.A1(new_n530), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n812), .A2(new_n521), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n810), .A2(new_n811), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n814), .A2(G860), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(KEYINPUT37), .Z(new_n816));
  NOR2_X1   g391(.A1(new_n628), .A2(new_n625), .ZN(new_n817));
  XNOR2_X1  g392(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT102), .ZN(new_n820));
  OR2_X1    g395(.A1(new_n814), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n814), .A2(new_n820), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n821), .A2(new_n570), .A3(new_n822), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n569), .A2(new_n814), .A3(new_n820), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n819), .B(new_n825), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n816), .B1(new_n826), .B2(G860), .ZN(G145));
  OR2_X1    g402(.A1(new_n468), .A2(G118), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n479), .B1(new_n828), .B2(KEYINPUT105), .ZN(new_n829));
  OAI221_X1 g404(.A(new_n829), .B1(KEYINPUT105), .B2(new_n828), .C1(G106), .C2(G2105), .ZN(new_n830));
  AOI22_X1  g405(.A1(G130), .A2(new_n492), .B1(new_n494), .B2(G142), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n832), .B(KEYINPUT106), .Z(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(new_n634), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n713), .B(KEYINPUT107), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(new_n514), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n506), .A2(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n765), .B(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(new_n742), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n841), .A2(new_n731), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(KEYINPUT103), .Z(new_n843));
  NAND2_X1  g418(.A1(new_n841), .A2(new_n731), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(KEYINPUT104), .Z(new_n845));
  NAND2_X1  g420(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n837), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n836), .A2(new_n843), .A3(new_n845), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n490), .B(new_n643), .Z(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(G162), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n847), .A2(new_n848), .A3(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(G37), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n847), .A2(new_n848), .ZN(new_n854));
  AOI21_X1  g429(.A(KEYINPUT108), .B1(new_n854), .B2(new_n850), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT108), .ZN(new_n856));
  AOI211_X1 g431(.A(new_n856), .B(new_n851), .C1(new_n847), .C2(new_n848), .ZN(new_n857));
  OAI211_X1 g432(.A(new_n852), .B(new_n853), .C1(new_n855), .C2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g434(.A1(new_n814), .A2(new_n621), .ZN(new_n860));
  INV_X1    g435(.A(G288), .ZN(new_n861));
  XNOR2_X1  g436(.A(G166), .B(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(G305), .ZN(new_n863));
  OR2_X1    g438(.A1(new_n863), .A2(G290), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(G290), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT42), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n825), .B(new_n629), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n628), .B(G299), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n869), .B(KEYINPUT41), .Z(new_n872));
  AOI21_X1  g447(.A(new_n871), .B1(new_n868), .B2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n867), .B(new_n873), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n860), .B1(new_n874), .B2(new_n621), .ZN(G295));
  OAI21_X1  g450(.A(new_n860), .B1(new_n874), .B2(new_n621), .ZN(G331));
  OR2_X1    g451(.A1(new_n866), .A2(KEYINPUT109), .ZN(new_n877));
  XNOR2_X1  g452(.A(G168), .B(G171), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n825), .B(new_n878), .ZN(new_n879));
  OR2_X1    g454(.A1(new_n879), .A2(new_n870), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n872), .A2(new_n879), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(G37), .B1(new_n877), .B2(new_n882), .ZN(new_n883));
  NAND4_X1  g458(.A1(new_n880), .A2(new_n864), .A3(new_n865), .A4(new_n881), .ZN(new_n884));
  OR2_X1    g459(.A1(new_n884), .A2(KEYINPUT109), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(KEYINPUT43), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n882), .A2(new_n866), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n888), .A2(new_n853), .A3(new_n884), .ZN(new_n889));
  OR2_X1    g464(.A1(new_n889), .A2(KEYINPUT43), .ZN(new_n890));
  AND2_X1   g465(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT43), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n883), .A2(new_n892), .A3(new_n885), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT44), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n894), .B1(new_n889), .B2(KEYINPUT43), .ZN(new_n895));
  AND3_X1   g470(.A1(new_n893), .A2(new_n895), .A3(KEYINPUT110), .ZN(new_n896));
  AOI21_X1  g471(.A(KEYINPUT110), .B1(new_n893), .B2(new_n895), .ZN(new_n897));
  OAI22_X1  g472(.A1(new_n891), .A2(KEYINPUT44), .B1(new_n896), .B2(new_n897), .ZN(G397));
  INV_X1    g473(.A(G1384), .ZN(new_n899));
  AOI21_X1  g474(.A(KEYINPUT45), .B1(new_n518), .B2(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n514), .B1(new_n505), .B2(new_n503), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT45), .ZN(new_n902));
  NOR3_X1   g477(.A1(new_n901), .A2(new_n902), .A3(G1384), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n488), .A2(new_n478), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n476), .B1(new_n470), .B2(new_n473), .ZN(new_n905));
  AND3_X1   g480(.A1(new_n470), .A2(new_n473), .A3(new_n476), .ZN(new_n906));
  OAI211_X1 g481(.A(new_n904), .B(G40), .C1(new_n905), .C2(new_n906), .ZN(new_n907));
  NOR3_X1   g482(.A1(new_n900), .A2(new_n903), .A3(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(KEYINPUT56), .B(G2072), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT50), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n518), .A2(new_n910), .A3(new_n899), .ZN(new_n911));
  INV_X1    g486(.A(G40), .ZN(new_n912));
  AOI221_X4 g487(.A(new_n912), .B1(new_n488), .B2(new_n478), .C1(new_n475), .C2(new_n477), .ZN(new_n913));
  OAI21_X1  g488(.A(KEYINPUT50), .B1(new_n901), .B2(G1384), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n911), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(G1956), .ZN(new_n916));
  AOI22_X1  g491(.A1(new_n908), .A2(new_n909), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT57), .ZN(new_n918));
  NAND2_X1  g493(.A1(G299), .A2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT119), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n583), .A2(new_n584), .A3(KEYINPUT57), .A4(new_n586), .ZN(new_n921));
  AND3_X1   g496(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n920), .B1(new_n919), .B2(new_n921), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n917), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(G1384), .B1(new_n506), .B2(new_n838), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(new_n910), .ZN(new_n927));
  AND3_X1   g502(.A1(new_n512), .A2(new_n516), .A3(new_n513), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n516), .B1(new_n512), .B2(new_n513), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(G1384), .B1(new_n930), .B2(new_n506), .ZN(new_n931));
  OAI211_X1 g506(.A(new_n913), .B(new_n927), .C1(new_n931), .C2(new_n910), .ZN(new_n932));
  INV_X1    g507(.A(G1348), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n839), .A2(new_n899), .ZN(new_n935));
  NOR3_X1   g510(.A1(new_n935), .A2(new_n907), .A3(G2067), .ZN(new_n936));
  INV_X1    g511(.A(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n628), .B1(new_n934), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n915), .A2(new_n916), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n903), .A2(new_n907), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n518), .A2(new_n899), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(new_n902), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n940), .A2(new_n942), .A3(new_n909), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n919), .A2(new_n921), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n939), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n925), .B1(new_n938), .B2(new_n945), .ZN(new_n946));
  AOI211_X1 g521(.A(new_n936), .B(new_n618), .C1(new_n933), .C2(new_n932), .ZN(new_n947));
  OAI21_X1  g522(.A(KEYINPUT60), .B1(new_n947), .B2(new_n938), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT59), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n926), .A2(KEYINPUT45), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n913), .A2(new_n950), .ZN(new_n951));
  NOR3_X1   g526(.A1(new_n951), .A2(G1996), .A3(new_n900), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n935), .A2(new_n907), .ZN(new_n953));
  XOR2_X1   g528(.A(KEYINPUT120), .B(G1341), .Z(new_n954));
  XNOR2_X1  g529(.A(new_n954), .B(KEYINPUT58), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n570), .B1(new_n952), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT122), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n949), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  OR2_X1    g534(.A1(new_n953), .A2(new_n955), .ZN(new_n960));
  INV_X1    g535(.A(G1996), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n940), .A2(new_n961), .A3(new_n942), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n569), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT121), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n963), .A2(new_n964), .A3(KEYINPUT122), .A4(KEYINPUT59), .ZN(new_n965));
  OAI211_X1 g540(.A(KEYINPUT61), .B(new_n945), .C1(new_n917), .C2(new_n924), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n948), .A2(new_n959), .A3(new_n965), .A4(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT61), .ZN(new_n968));
  AND3_X1   g543(.A1(new_n939), .A2(new_n943), .A3(new_n944), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n944), .B1(new_n939), .B2(new_n943), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n968), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n957), .A2(KEYINPUT121), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n628), .A2(KEYINPUT60), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n934), .A2(new_n937), .A3(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n971), .A2(new_n972), .A3(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n946), .B1(new_n967), .B2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT55), .ZN(new_n977));
  INV_X1    g552(.A(G8), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n977), .B1(G166), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(KEYINPUT115), .ZN(new_n980));
  NAND3_X1  g555(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT115), .ZN(new_n982));
  OAI211_X1 g557(.A(new_n982), .B(new_n977), .C1(G166), .C2(new_n978), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n980), .A2(new_n981), .A3(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT114), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n985), .B1(new_n951), .B2(new_n900), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n940), .A2(KEYINPUT114), .A3(new_n942), .ZN(new_n987));
  AOI21_X1  g562(.A(G1971), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n932), .A2(G2090), .ZN(new_n989));
  OAI211_X1 g564(.A(G8), .B(new_n984), .C1(new_n988), .C2(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n489), .A2(new_n926), .A3(G40), .ZN(new_n991));
  XNOR2_X1  g566(.A(KEYINPUT116), .B(G1976), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n991), .A2(G8), .A3(G288), .A4(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT117), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n861), .A2(G1976), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n991), .A2(new_n994), .A3(G8), .A4(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT52), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n993), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n993), .A2(new_n997), .ZN(new_n999));
  INV_X1    g574(.A(new_n996), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  AND2_X1   g576(.A1(new_n597), .A2(new_n599), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT118), .ZN(new_n1003));
  INV_X1    g578(.A(G1981), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n1002), .A2(new_n1003), .A3(new_n1004), .A4(new_n598), .ZN(new_n1005));
  OAI21_X1  g580(.A(KEYINPUT118), .B1(G305), .B2(G1981), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(G305), .A2(G1981), .ZN(new_n1008));
  AND3_X1   g583(.A1(new_n1007), .A2(KEYINPUT49), .A3(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(KEYINPUT49), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n953), .A2(new_n978), .ZN(new_n1012));
  AOI22_X1  g587(.A1(new_n998), .A2(new_n1001), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(G1971), .ZN(new_n1014));
  AOI21_X1  g589(.A(KEYINPUT114), .B1(new_n940), .B2(new_n942), .ZN(new_n1015));
  NOR4_X1   g590(.A1(new_n900), .A2(new_n903), .A3(new_n985), .A4(new_n907), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1014), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  OR2_X1    g592(.A1(new_n915), .A2(G2090), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n978), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  OAI211_X1 g594(.A(new_n990), .B(new_n1013), .C1(new_n1019), .C2(new_n984), .ZN(new_n1020));
  INV_X1    g595(.A(G2078), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n986), .A2(new_n1021), .A3(new_n987), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT53), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G1961), .ZN(new_n1025));
  AND3_X1   g600(.A1(new_n932), .A2(KEYINPUT124), .A3(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(KEYINPUT124), .B1(new_n932), .B2(new_n1025), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  XOR2_X1   g603(.A(G301), .B(KEYINPUT54), .Z(new_n1029));
  NAND2_X1  g604(.A1(new_n935), .A2(new_n902), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1030), .A2(KEYINPUT53), .A3(new_n1021), .A4(new_n913), .ZN(new_n1031));
  OR2_X1    g606(.A1(new_n1031), .A2(new_n903), .ZN(new_n1032));
  AND4_X1   g607(.A1(new_n1024), .A2(new_n1028), .A3(new_n1029), .A4(new_n1032), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1020), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT51), .ZN(new_n1035));
  NAND2_X1  g610(.A1(G286), .A2(G8), .ZN(new_n1036));
  INV_X1    g611(.A(new_n932), .ZN(new_n1037));
  INV_X1    g612(.A(G2084), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n1030), .B(new_n913), .C1(new_n902), .C2(new_n941), .ZN(new_n1039));
  AOI22_X1  g614(.A1(new_n1037), .A2(new_n1038), .B1(new_n1039), .B2(new_n785), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n1035), .B(new_n1036), .C1(new_n1040), .C2(new_n978), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1039), .A2(new_n785), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n907), .B1(new_n941), .B2(KEYINPUT50), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1043), .A2(new_n1038), .A3(new_n927), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1045));
  OAI211_X1 g620(.A(KEYINPUT51), .B(G8), .C1(new_n1045), .C2(G286), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1041), .A2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1045), .A2(G8), .A3(G286), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n932), .A2(new_n1025), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n941), .A2(new_n902), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1049), .B1(new_n1050), .B2(new_n1031), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(KEYINPUT123), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT123), .ZN(new_n1053));
  OAI211_X1 g628(.A(new_n1049), .B(new_n1053), .C1(new_n1031), .C2(new_n1050), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1052), .A2(new_n1024), .A3(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1029), .ZN(new_n1056));
  AOI22_X1  g631(.A1(new_n1047), .A2(new_n1048), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n976), .A2(new_n1034), .A3(new_n1057), .ZN(new_n1058));
  AOI21_X1  g633(.A(G1976), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(new_n861), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(new_n1007), .ZN(new_n1061));
  INV_X1    g636(.A(new_n990), .ZN(new_n1062));
  AOI22_X1  g637(.A1(new_n1061), .A2(new_n1012), .B1(new_n1062), .B2(new_n1013), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT63), .ZN(new_n1064));
  NOR3_X1   g639(.A1(new_n1040), .A2(new_n978), .A3(G286), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1064), .B1(new_n1020), .B2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(G8), .B1(new_n988), .B2(new_n989), .ZN(new_n1068));
  INV_X1    g643(.A(new_n984), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1064), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1070), .A2(new_n990), .A3(new_n1013), .A4(new_n1065), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1067), .A2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1058), .A2(new_n1063), .A3(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT125), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1076), .A2(KEYINPUT62), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1077), .A2(new_n1020), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1076), .A2(KEYINPUT62), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1078), .A2(G171), .A3(new_n1055), .A4(new_n1079), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1058), .A2(new_n1072), .A3(KEYINPUT125), .A4(new_n1063), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1075), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n926), .A2(KEYINPUT45), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(new_n913), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1084), .A2(G1996), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(new_n743), .ZN(new_n1086));
  XNOR2_X1  g661(.A(new_n1086), .B(KEYINPUT111), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1084), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n765), .A2(G2067), .ZN(new_n1089));
  INV_X1    g664(.A(G2067), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n759), .A2(new_n1090), .A3(new_n764), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1088), .A2(new_n1092), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1084), .A2(new_n743), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1094), .ZN(new_n1095));
  OAI211_X1 g670(.A(new_n1087), .B(new_n1093), .C1(new_n961), .C2(new_n1095), .ZN(new_n1096));
  OR2_X1    g671(.A1(new_n1096), .A2(KEYINPUT112), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(KEYINPUT112), .ZN(new_n1098));
  XNOR2_X1  g673(.A(new_n713), .B(new_n715), .ZN(new_n1099));
  XOR2_X1   g674(.A(new_n1099), .B(KEYINPUT113), .Z(new_n1100));
  OAI211_X1 g675(.A(new_n1097), .B(new_n1098), .C1(new_n1084), .C2(new_n1100), .ZN(new_n1101));
  XNOR2_X1  g676(.A(G290), .B(G1986), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1101), .B1(new_n1088), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1082), .A2(new_n1103), .ZN(new_n1104));
  NOR3_X1   g679(.A1(new_n1084), .A2(G1986), .A3(G290), .ZN(new_n1105));
  XNOR2_X1  g680(.A(new_n1105), .B(KEYINPUT48), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1101), .A2(new_n1106), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n713), .A2(new_n715), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1097), .A2(new_n1098), .A3(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1084), .B1(new_n1109), .B2(new_n1091), .ZN(new_n1110));
  AND3_X1   g685(.A1(new_n1095), .A2(KEYINPUT126), .A3(new_n1093), .ZN(new_n1111));
  AOI21_X1  g686(.A(KEYINPUT126), .B1(new_n1095), .B2(new_n1093), .ZN(new_n1112));
  AND2_X1   g687(.A1(new_n1085), .A2(KEYINPUT46), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1085), .A2(KEYINPUT46), .ZN(new_n1114));
  NOR4_X1   g689(.A1(new_n1111), .A2(new_n1112), .A3(new_n1113), .A4(new_n1114), .ZN(new_n1115));
  XNOR2_X1  g690(.A(new_n1115), .B(KEYINPUT47), .ZN(new_n1116));
  NOR3_X1   g691(.A1(new_n1107), .A2(new_n1110), .A3(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1104), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(KEYINPUT127), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT127), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1104), .A2(new_n1120), .A3(new_n1117), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1119), .A2(new_n1121), .ZN(G329));
  assign    G231 = 1'b0;
  AOI211_X1 g697(.A(new_n462), .B(G229), .C1(new_n887), .C2(new_n890), .ZN(new_n1124));
  NOR2_X1   g698(.A1(G401), .A2(G227), .ZN(new_n1125));
  AND3_X1   g699(.A1(new_n1124), .A2(new_n858), .A3(new_n1125), .ZN(G308));
  NAND3_X1  g700(.A1(new_n1124), .A2(new_n858), .A3(new_n1125), .ZN(G225));
endmodule


