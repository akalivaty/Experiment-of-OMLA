//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 0 0 0 1 0 0 0 1 0 0 1 1 0 1 0 1 1 1 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 1 1 1 1 0 0 0 0 1 1 1 0 1 0 1 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:30 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1065, new_n1066,
    new_n1067, new_n1068, new_n1069, new_n1070, new_n1071, new_n1072,
    new_n1073, new_n1075, new_n1076, new_n1077, new_n1078, new_n1079,
    new_n1080, new_n1081, new_n1082, new_n1083, new_n1084, new_n1085,
    new_n1086;
  INV_X1    g000(.A(KEYINPUT94), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT20), .ZN(new_n188));
  XNOR2_X1  g002(.A(G113), .B(G122), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT92), .B(G104), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G140), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G125), .ZN(new_n193));
  INV_X1    g007(.A(G125), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G140), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n193), .A2(new_n195), .A3(KEYINPUT76), .ZN(new_n196));
  OR3_X1    g010(.A1(new_n192), .A2(KEYINPUT76), .A3(G125), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(KEYINPUT90), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT90), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n196), .A2(new_n197), .A3(new_n200), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n199), .A2(KEYINPUT19), .A3(new_n201), .ZN(new_n202));
  AND2_X1   g016(.A1(KEYINPUT64), .A2(G146), .ZN(new_n203));
  NOR2_X1   g017(.A1(KEYINPUT64), .A2(G146), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n193), .A2(new_n195), .ZN(new_n206));
  OR2_X1    g020(.A1(new_n206), .A2(KEYINPUT19), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n202), .A2(new_n205), .A3(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G146), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n196), .A2(new_n197), .A3(KEYINPUT16), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT16), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n193), .A2(new_n211), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n209), .B1(new_n210), .B2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G131), .ZN(new_n215));
  INV_X1    g029(.A(G143), .ZN(new_n216));
  INV_X1    g030(.A(G237), .ZN(new_n217));
  INV_X1    g031(.A(G953), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G214), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n216), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(G143), .A2(G214), .ZN(new_n222));
  NOR4_X1   g036(.A1(new_n222), .A2(KEYINPUT88), .A3(G237), .A4(G953), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT88), .ZN(new_n224));
  AND2_X1   g038(.A1(G143), .A2(G214), .ZN(new_n225));
  NOR2_X1   g039(.A1(G237), .A2(G953), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n224), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  OAI211_X1 g041(.A(new_n215), .B(new_n221), .C1(new_n223), .C2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(KEYINPUT91), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n221), .B1(new_n223), .B2(new_n227), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G131), .ZN(new_n231));
  AOI21_X1  g045(.A(G143), .B1(new_n226), .B2(G214), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n232), .A2(G131), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT91), .ZN(new_n234));
  OAI211_X1 g048(.A(new_n233), .B(new_n234), .C1(new_n223), .C2(new_n227), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n229), .A2(new_n231), .A3(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n208), .A2(new_n214), .A3(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n199), .A2(G146), .A3(new_n201), .ZN(new_n238));
  XNOR2_X1  g052(.A(KEYINPUT64), .B(G146), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n206), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n238), .A2(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(KEYINPUT88), .B1(new_n219), .B2(new_n222), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n225), .A2(new_n226), .A3(new_n224), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n232), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(KEYINPUT18), .A2(G131), .ZN(new_n246));
  OAI21_X1  g060(.A(KEYINPUT89), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT89), .ZN(new_n248));
  INV_X1    g062(.A(new_n246), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n230), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n247), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n245), .A2(new_n246), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n242), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n191), .B1(new_n237), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT17), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n229), .A2(new_n231), .A3(new_n235), .A4(new_n255), .ZN(new_n256));
  AND3_X1   g070(.A1(new_n210), .A2(new_n209), .A3(new_n212), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n257), .A2(new_n213), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n230), .A2(KEYINPUT17), .A3(G131), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n256), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n260), .A2(new_n253), .A3(new_n191), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT93), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n260), .A2(new_n253), .A3(KEYINPUT93), .A4(new_n191), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n254), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NOR2_X1   g079(.A1(G475), .A2(G902), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n187), .B(new_n188), .C1(new_n265), .C2(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n191), .B1(new_n260), .B2(new_n253), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n269), .B1(new_n263), .B2(new_n264), .ZN(new_n270));
  OAI21_X1  g084(.A(G475), .B1(new_n270), .B2(G902), .ZN(new_n271));
  AND2_X1   g085(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n263), .A2(new_n264), .ZN(new_n273));
  INV_X1    g087(.A(new_n254), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n275), .A2(KEYINPUT94), .A3(new_n266), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n187), .B1(new_n265), .B2(new_n267), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n276), .A2(KEYINPUT20), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n272), .A2(new_n278), .ZN(new_n279));
  AND2_X1   g093(.A1(new_n218), .A2(G952), .ZN(new_n280));
  INV_X1    g094(.A(G234), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n280), .B1(new_n281), .B2(new_n217), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  XNOR2_X1  g097(.A(KEYINPUT21), .B(G898), .ZN(new_n284));
  XNOR2_X1  g098(.A(new_n284), .B(KEYINPUT97), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(G902), .ZN(new_n287));
  AOI211_X1 g101(.A(new_n287), .B(new_n218), .C1(G234), .C2(G237), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n283), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(G116), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n290), .A2(KEYINPUT14), .A3(G122), .ZN(new_n291));
  XOR2_X1   g105(.A(G116), .B(G122), .Z(new_n292));
  OAI211_X1 g106(.A(G107), .B(new_n291), .C1(new_n292), .C2(KEYINPUT14), .ZN(new_n293));
  XNOR2_X1  g107(.A(G116), .B(G122), .ZN(new_n294));
  INV_X1    g108(.A(G107), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  XNOR2_X1  g110(.A(KEYINPUT65), .B(G134), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n216), .A2(G128), .ZN(new_n298));
  INV_X1    g112(.A(G128), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G143), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n297), .A2(new_n298), .A3(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n297), .B1(new_n298), .B2(new_n300), .ZN(new_n303));
  OAI211_X1 g117(.A(new_n293), .B(new_n296), .C1(new_n302), .C2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n292), .A2(G107), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(new_n296), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT13), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n298), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(new_n300), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n298), .A2(new_n307), .ZN(new_n310));
  OAI21_X1  g124(.A(G134), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n306), .A2(new_n311), .A3(new_n301), .ZN(new_n312));
  XNOR2_X1  g126(.A(KEYINPUT9), .B(G234), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT79), .ZN(new_n314));
  XNOR2_X1  g128(.A(new_n313), .B(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n218), .A2(G217), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  AND3_X1   g131(.A1(new_n304), .A2(new_n312), .A3(new_n317), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n317), .B1(new_n304), .B2(new_n312), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n287), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(KEYINPUT95), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT95), .ZN(new_n322));
  OAI211_X1 g136(.A(new_n322), .B(new_n287), .C1(new_n318), .C2(new_n319), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(G478), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n325), .A2(KEYINPUT15), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n324), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT96), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n323), .A2(new_n326), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n326), .B1(new_n321), .B2(new_n323), .ZN(new_n332));
  INV_X1    g146(.A(new_n330), .ZN(new_n333));
  OAI21_X1  g147(.A(KEYINPUT96), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n331), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NOR3_X1   g150(.A1(new_n279), .A2(new_n289), .A3(new_n336), .ZN(new_n337));
  OAI21_X1  g151(.A(G221), .B1(new_n315), .B2(G902), .ZN(new_n338));
  XOR2_X1   g152(.A(new_n338), .B(KEYINPUT80), .Z(new_n339));
  INV_X1    g153(.A(G469), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n340), .A2(new_n287), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT64), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(new_n209), .ZN(new_n343));
  NAND2_X1  g157(.A1(KEYINPUT64), .A2(G146), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n343), .A2(G143), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n216), .A2(G146), .ZN(new_n346));
  AND2_X1   g160(.A1(KEYINPUT0), .A2(G128), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n209), .A2(G143), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n350), .B1(new_n239), .B2(new_n216), .ZN(new_n351));
  NOR2_X1   g165(.A1(KEYINPUT0), .A2(G128), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n347), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n348), .B1(new_n351), .B2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT4), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n295), .A2(G104), .ZN(new_n358));
  OR2_X1    g172(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n359));
  NAND2_X1  g173(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n358), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(G104), .ZN(new_n362));
  OAI22_X1  g176(.A1(new_n362), .A2(G107), .B1(KEYINPUT81), .B2(KEYINPUT3), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(G107), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n357), .B(G101), .C1(new_n361), .C2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n356), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n359), .A2(new_n360), .ZN(new_n368));
  INV_X1    g182(.A(new_n358), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(G101), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n370), .A2(new_n371), .A3(new_n364), .A4(new_n363), .ZN(new_n372));
  OAI21_X1  g186(.A(G101), .B1(new_n361), .B2(new_n365), .ZN(new_n373));
  AND3_X1   g187(.A1(new_n372), .A2(KEYINPUT4), .A3(new_n373), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n367), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n358), .A2(new_n364), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(G101), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT1), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n345), .A2(new_n378), .A3(G128), .A4(new_n346), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n299), .B1(new_n349), .B2(KEYINPUT1), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n381), .B1(new_n345), .B2(new_n346), .ZN(new_n382));
  OAI211_X1 g196(.A(new_n372), .B(new_n377), .C1(new_n380), .C2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT10), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT82), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n383), .A2(KEYINPUT82), .A3(new_n384), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n375), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NOR3_X1   g203(.A1(new_n203), .A2(new_n204), .A3(new_n216), .ZN(new_n390));
  OAI21_X1  g204(.A(G128), .B1(new_n390), .B2(new_n378), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n349), .B1(new_n205), .B2(G143), .ZN(new_n392));
  AOI21_X1  g206(.A(KEYINPUT67), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n299), .B1(new_n345), .B2(KEYINPUT1), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT67), .ZN(new_n395));
  NOR3_X1   g209(.A1(new_n394), .A2(new_n351), .A3(new_n395), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n379), .B1(new_n393), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(KEYINPUT70), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n395), .B1(new_n394), .B2(new_n351), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n378), .B1(new_n205), .B2(G143), .ZN(new_n400));
  OAI211_X1 g214(.A(KEYINPUT67), .B(new_n392), .C1(new_n400), .C2(new_n299), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT70), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n402), .A2(new_n403), .A3(new_n379), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n372), .A2(new_n377), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n405), .A2(new_n384), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n398), .A2(new_n404), .A3(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT11), .ZN(new_n408));
  INV_X1    g222(.A(G134), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(KEYINPUT65), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT65), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(G134), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n410), .A2(new_n412), .A3(G137), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n409), .A2(G137), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n408), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n410), .A2(new_n412), .ZN(new_n417));
  INV_X1    g231(.A(G137), .ZN(new_n418));
  AOI21_X1  g232(.A(KEYINPUT11), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(G131), .B1(new_n416), .B2(new_n419), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n408), .B1(new_n297), .B2(G137), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n414), .B1(new_n297), .B2(G137), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n215), .B(new_n421), .C1(new_n422), .C2(new_n408), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n420), .A2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n389), .A2(new_n407), .A3(new_n425), .ZN(new_n426));
  XNOR2_X1  g240(.A(G110), .B(G140), .ZN(new_n427));
  AND2_X1   g241(.A1(new_n218), .A2(G227), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n427), .B(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n380), .B1(new_n372), .B2(new_n377), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n402), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT83), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n402), .A2(new_n431), .A3(KEYINPUT83), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n434), .A2(new_n383), .A3(new_n435), .ZN(new_n436));
  AND3_X1   g250(.A1(new_n436), .A2(KEYINPUT12), .A3(new_n424), .ZN(new_n437));
  AOI21_X1  g251(.A(KEYINPUT12), .B1(new_n436), .B2(new_n424), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n426), .B(new_n430), .C1(new_n437), .C2(new_n438), .ZN(new_n439));
  AND3_X1   g253(.A1(new_n389), .A2(new_n407), .A3(new_n425), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n425), .B1(new_n389), .B2(new_n407), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n429), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(G902), .B1(new_n439), .B2(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n341), .B1(new_n443), .B2(new_n340), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n426), .B1(new_n437), .B2(new_n438), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n429), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n440), .A2(new_n429), .ZN(new_n447));
  AND3_X1   g261(.A1(new_n398), .A2(new_n404), .A3(new_n406), .ZN(new_n448));
  AND3_X1   g262(.A1(new_n383), .A2(KEYINPUT82), .A3(new_n384), .ZN(new_n449));
  AOI21_X1  g263(.A(KEYINPUT82), .B1(new_n383), .B2(new_n384), .ZN(new_n450));
  OAI22_X1  g264(.A1(new_n449), .A2(new_n450), .B1(new_n374), .B2(new_n367), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n424), .B1(new_n448), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n447), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n446), .A2(new_n453), .A3(G469), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n339), .B1(new_n444), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(G214), .B1(G237), .B2(G902), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(G210), .B1(G237), .B2(G902), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  XNOR2_X1  g273(.A(G110), .B(G122), .ZN(new_n460));
  XOR2_X1   g274(.A(new_n460), .B(KEYINPUT8), .Z(new_n461));
  XNOR2_X1  g275(.A(G116), .B(G119), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(KEYINPUT5), .ZN(new_n463));
  OR3_X1    g277(.A1(new_n290), .A2(KEYINPUT5), .A3(G119), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n463), .A2(G113), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(KEYINPUT2), .A2(G113), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT69), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n466), .B(new_n467), .ZN(new_n468));
  NOR2_X1   g282(.A1(KEYINPUT2), .A2(G113), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(KEYINPUT68), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT68), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n471), .B1(KEYINPUT2), .B2(G113), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n468), .A2(new_n462), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n465), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n405), .A2(new_n475), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n372), .A2(new_n474), .A3(new_n465), .A4(new_n377), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n461), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n379), .A2(new_n194), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n402), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n355), .A2(G125), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(G224), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n484), .A2(G953), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(KEYINPUT7), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n478), .B1(new_n483), .B2(new_n487), .ZN(new_n488));
  OR2_X1    g302(.A1(new_n486), .A2(KEYINPUT85), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n486), .A2(KEYINPUT85), .ZN(new_n490));
  AND2_X1   g304(.A1(new_n490), .A2(KEYINPUT7), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n482), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n479), .B1(new_n399), .B2(new_n401), .ZN(new_n493));
  OAI21_X1  g307(.A(KEYINPUT86), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n491), .A2(new_n489), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n495), .B1(new_n355), .B2(G125), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT86), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n481), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n494), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n488), .A2(new_n499), .A3(KEYINPUT87), .ZN(new_n500));
  INV_X1    g314(.A(new_n474), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n462), .B1(new_n468), .B2(new_n473), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n366), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n477), .B(new_n460), .C1(new_n503), .C2(new_n374), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n500), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(KEYINPUT87), .B1(new_n488), .B2(new_n499), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT84), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n481), .A2(new_n508), .A3(new_n482), .ZN(new_n509));
  INV_X1    g323(.A(new_n482), .ZN(new_n510));
  OAI21_X1  g324(.A(KEYINPUT84), .B1(new_n493), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(new_n486), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n477), .B1(new_n503), .B2(new_n374), .ZN(new_n514));
  INV_X1    g328(.A(new_n460), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n516), .A2(KEYINPUT6), .A3(new_n504), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n509), .A2(new_n511), .A3(new_n485), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT6), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n514), .A2(new_n519), .A3(new_n515), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n513), .A2(new_n517), .A3(new_n518), .A4(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n287), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n459), .B1(new_n507), .B2(new_n522), .ZN(new_n523));
  AND2_X1   g337(.A1(new_n517), .A2(new_n520), .ZN(new_n524));
  INV_X1    g338(.A(new_n518), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n485), .B1(new_n509), .B2(new_n511), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(G902), .B1(new_n524), .B2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n506), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n529), .A2(new_n504), .A3(new_n500), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n528), .A2(new_n530), .A3(new_n458), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n457), .B1(new_n523), .B2(new_n531), .ZN(new_n532));
  AND3_X1   g346(.A1(new_n337), .A2(new_n455), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n417), .A2(new_n418), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n409), .A2(G137), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(G131), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n423), .A2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n398), .A2(new_n404), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n355), .B1(new_n420), .B2(new_n423), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n501), .A2(new_n502), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(KEYINPUT71), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT71), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n544), .B1(new_n501), .B2(new_n502), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n541), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(KEYINPUT28), .B1(new_n540), .B2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT72), .ZN(new_n549));
  AND3_X1   g363(.A1(new_n540), .A2(new_n549), .A3(new_n546), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n549), .B1(new_n540), .B2(new_n546), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT66), .ZN(new_n552));
  AOI22_X1  g366(.A1(new_n402), .A2(new_n379), .B1(new_n538), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n423), .A2(new_n537), .A3(KEYINPUT66), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n541), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n555), .A2(new_n542), .ZN(new_n556));
  NOR3_X1   g370(.A1(new_n550), .A2(new_n551), .A3(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT28), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n548), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n226), .A2(G210), .ZN(new_n560));
  XOR2_X1   g374(.A(new_n560), .B(KEYINPUT27), .Z(new_n561));
  XNOR2_X1  g375(.A(KEYINPUT26), .B(G101), .ZN(new_n562));
  XOR2_X1   g376(.A(new_n561), .B(new_n562), .Z(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  NOR3_X1   g378(.A1(new_n416), .A2(new_n419), .A3(G131), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n215), .B1(new_n534), .B2(new_n535), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n552), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n397), .A2(new_n567), .A3(new_n554), .ZN(new_n568));
  INV_X1    g382(.A(new_n541), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT30), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n542), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n540), .A2(KEYINPUT30), .A3(new_n569), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n540), .A2(new_n546), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(KEYINPUT72), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n540), .A2(new_n549), .A3(new_n546), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n574), .A2(new_n576), .A3(new_n577), .A4(new_n563), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT31), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n550), .A2(new_n551), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n581), .A2(KEYINPUT31), .A3(new_n563), .A4(new_n574), .ZN(new_n582));
  AOI22_X1  g396(.A1(new_n559), .A2(new_n564), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(KEYINPUT73), .B1(G472), .B2(G902), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NOR3_X1   g399(.A1(KEYINPUT73), .A2(G472), .A3(G902), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  OAI21_X1  g401(.A(KEYINPUT32), .B1(new_n583), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n559), .A2(new_n564), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n580), .A2(new_n582), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT32), .ZN(new_n592));
  INV_X1    g406(.A(new_n587), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n574), .A2(new_n576), .A3(new_n577), .ZN(new_n595));
  AOI21_X1  g409(.A(KEYINPUT29), .B1(new_n595), .B2(new_n564), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n596), .B1(new_n559), .B2(new_n564), .ZN(new_n597));
  AND2_X1   g411(.A1(new_n563), .A2(KEYINPUT29), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n576), .A2(new_n577), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n540), .A2(new_n569), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n543), .A2(new_n545), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(KEYINPUT74), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT74), .ZN(new_n605));
  AOI211_X1 g419(.A(new_n605), .B(new_n601), .C1(new_n540), .C2(new_n569), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n599), .B1(new_n604), .B2(new_n607), .ZN(new_n608));
  OAI211_X1 g422(.A(new_n548), .B(new_n598), .C1(new_n608), .C2(new_n558), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n597), .A2(new_n609), .A3(new_n287), .ZN(new_n610));
  AOI22_X1  g424(.A1(new_n588), .A2(new_n594), .B1(G472), .B2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(G217), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n612), .B1(G234), .B2(new_n287), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT25), .ZN(new_n615));
  OAI21_X1  g429(.A(KEYINPUT23), .B1(new_n299), .B2(G119), .ZN(new_n616));
  AOI21_X1  g430(.A(KEYINPUT75), .B1(new_n299), .B2(G119), .ZN(new_n617));
  OR2_X1    g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n616), .A2(new_n617), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(G110), .ZN(new_n621));
  XOR2_X1   g435(.A(G119), .B(G128), .Z(new_n622));
  XNOR2_X1  g436(.A(KEYINPUT24), .B(G110), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  OR2_X1    g438(.A1(new_n624), .A2(new_n258), .ZN(new_n625));
  XNOR2_X1  g439(.A(KEYINPUT77), .B(G110), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n618), .A2(new_n619), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n622), .A2(new_n623), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n240), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(new_n214), .ZN(new_n630));
  XNOR2_X1  g444(.A(KEYINPUT22), .B(G137), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n218), .A2(G221), .A3(G234), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n625), .A2(new_n630), .A3(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n633), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n624), .A2(new_n258), .ZN(new_n636));
  INV_X1    g450(.A(new_n630), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n635), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n615), .B1(new_n639), .B2(G902), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n634), .A2(new_n638), .A3(KEYINPUT25), .A4(new_n287), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n614), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n613), .A2(G902), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n634), .A2(new_n638), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  NOR3_X1   g460(.A1(new_n611), .A2(KEYINPUT78), .A3(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT78), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n610), .A2(G472), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n592), .B1(new_n591), .B2(new_n593), .ZN(new_n650));
  AOI211_X1 g464(.A(KEYINPUT32), .B(new_n587), .C1(new_n589), .C2(new_n590), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n649), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n646), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n648), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n533), .B1(new_n647), .B2(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT98), .B(G101), .Z(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G3));
  OAI21_X1  g471(.A(G472), .B1(new_n583), .B2(G902), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n591), .A2(new_n593), .ZN(new_n659));
  AND2_X1   g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n439), .A2(new_n442), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n661), .A2(new_n340), .A3(new_n287), .ZN(new_n662));
  INV_X1    g476(.A(new_n341), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n662), .A2(new_n454), .A3(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n339), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n666), .A2(new_n646), .ZN(new_n667));
  AND2_X1   g481(.A1(new_n660), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n318), .A2(new_n319), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT33), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n670), .A2(KEYINPUT99), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  AND2_X1   g486(.A1(new_n670), .A2(KEYINPUT99), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n672), .B(new_n674), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n325), .A2(G902), .ZN(new_n676));
  AOI22_X1  g490(.A1(new_n675), .A2(new_n676), .B1(new_n325), .B2(new_n320), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n677), .B1(new_n272), .B2(new_n278), .ZN(new_n678));
  INV_X1    g492(.A(new_n289), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n678), .A2(new_n532), .A3(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n668), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(KEYINPUT34), .B(G104), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(KEYINPUT100), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n682), .B(new_n684), .ZN(G6));
  NOR3_X1   g499(.A1(new_n507), .A2(new_n522), .A3(new_n459), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n458), .B1(new_n528), .B2(new_n530), .ZN(new_n687));
  OAI211_X1 g501(.A(new_n456), .B(new_n679), .C1(new_n686), .C2(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n336), .A2(new_n272), .A3(new_n278), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n668), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g505(.A(KEYINPUT35), .B(G107), .Z(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G9));
  NOR2_X1   g507(.A1(new_n635), .A2(KEYINPUT36), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n625), .A2(new_n630), .A3(new_n694), .ZN(new_n695));
  OAI22_X1  g509(.A1(new_n636), .A2(new_n637), .B1(KEYINPUT36), .B2(new_n635), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n695), .A2(new_n696), .A3(new_n644), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(KEYINPUT101), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n642), .A2(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n533), .A2(new_n660), .A3(new_n700), .ZN(new_n701));
  XOR2_X1   g515(.A(KEYINPUT37), .B(G110), .Z(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(G12));
  NAND2_X1  g517(.A1(new_n532), .A2(new_n700), .ZN(new_n704));
  INV_X1    g518(.A(G900), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n283), .B1(new_n288), .B2(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n336), .A2(new_n272), .A3(new_n278), .A4(new_n707), .ZN(new_n708));
  NOR3_X1   g522(.A1(new_n666), .A2(new_n704), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n652), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G128), .ZN(G30));
  XOR2_X1   g525(.A(new_n706), .B(KEYINPUT39), .Z(new_n712));
  NAND2_X1  g526(.A1(new_n455), .A2(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT104), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n713), .A2(new_n714), .ZN(new_n717));
  OAI21_X1  g531(.A(KEYINPUT40), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n595), .A2(new_n563), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n581), .B1(new_n603), .B2(new_n606), .ZN(new_n720));
  OAI211_X1 g534(.A(new_n719), .B(new_n287), .C1(new_n563), .C2(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(G472), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n722), .B1(new_n650), .B2(new_n651), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n523), .A2(new_n531), .ZN(new_n724));
  XNOR2_X1  g538(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(KEYINPUT102), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n724), .B(new_n726), .ZN(new_n727));
  NOR3_X1   g541(.A1(new_n700), .A2(new_n457), .A3(new_n335), .ZN(new_n728));
  AND4_X1   g542(.A1(new_n279), .A2(new_n723), .A3(new_n727), .A4(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(new_n717), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT40), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n730), .A2(new_n731), .A3(new_n715), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n718), .A2(new_n729), .A3(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT105), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n733), .B(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G143), .ZN(G45));
  AND3_X1   g550(.A1(new_n724), .A2(new_n700), .A3(new_n456), .ZN(new_n737));
  AOI211_X1 g551(.A(new_n677), .B(new_n706), .C1(new_n272), .C2(new_n278), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n737), .A2(new_n455), .A3(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n652), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G146), .ZN(G48));
  AOI21_X1  g556(.A(new_n339), .B1(new_n443), .B2(new_n340), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n443), .A2(KEYINPUT106), .ZN(new_n744));
  INV_X1    g558(.A(new_n744), .ZN(new_n745));
  OAI21_X1  g559(.A(G469), .B1(new_n443), .B2(KEYINPUT106), .ZN(new_n746));
  OAI211_X1 g560(.A(new_n653), .B(new_n743), .C1(new_n745), .C2(new_n746), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n747), .A2(new_n680), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n652), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(KEYINPUT41), .B(G113), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n749), .B(new_n750), .ZN(G15));
  NOR3_X1   g565(.A1(new_n747), .A2(new_n688), .A3(new_n689), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(new_n652), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G116), .ZN(G18));
  NAND2_X1  g568(.A1(new_n662), .A2(new_n665), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n661), .A2(new_n287), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT106), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n340), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n755), .B1(new_n758), .B2(new_n744), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n652), .A2(new_n337), .A3(new_n737), .A4(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G119), .ZN(G21));
  AOI21_X1  g575(.A(new_n547), .B1(new_n720), .B2(KEYINPUT28), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n590), .B1(new_n762), .B2(new_n563), .ZN(new_n763));
  XOR2_X1   g577(.A(new_n587), .B(KEYINPUT107), .Z(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  AND2_X1   g579(.A1(new_n658), .A2(new_n765), .ZN(new_n766));
  AND3_X1   g580(.A1(new_n532), .A2(new_n279), .A3(new_n336), .ZN(new_n767));
  OAI211_X1 g581(.A(new_n679), .B(new_n743), .C1(new_n745), .C2(new_n746), .ZN(new_n768));
  INV_X1    g582(.A(new_n768), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n766), .A2(new_n653), .A3(new_n767), .A4(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G122), .ZN(G24));
  NAND3_X1  g585(.A1(new_n658), .A2(new_n765), .A3(new_n700), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n436), .A2(new_n424), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT12), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n436), .A2(KEYINPUT12), .A3(new_n424), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n452), .A2(new_n426), .ZN(new_n778));
  AOI22_X1  g592(.A1(new_n447), .A2(new_n777), .B1(new_n778), .B2(new_n429), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n757), .B1(new_n779), .B2(G902), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n780), .A2(G469), .A3(new_n744), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n738), .A2(new_n781), .A3(new_n532), .A4(new_n743), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n772), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(new_n194), .ZN(G27));
  INV_X1    g598(.A(KEYINPUT108), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n454), .A2(new_n785), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n446), .A2(new_n453), .A3(KEYINPUT108), .A4(G469), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n786), .A2(new_n444), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n665), .A2(new_n456), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n724), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n788), .A2(new_n738), .A3(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n652), .A2(new_n792), .A3(new_n653), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT42), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n652), .A2(new_n792), .A3(KEYINPUT42), .A4(new_n653), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G131), .ZN(G33));
  NAND2_X1  g612(.A1(new_n268), .A2(new_n271), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n277), .A2(KEYINPUT20), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n799), .B1(new_n800), .B2(new_n276), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT109), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n801), .A2(new_n802), .A3(new_n336), .A4(new_n707), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n708), .A2(KEYINPUT109), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n803), .A2(new_n804), .A3(new_n788), .A4(new_n790), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n611), .A2(new_n805), .A3(new_n646), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(new_n409), .ZN(G36));
  INV_X1    g621(.A(KEYINPUT112), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n446), .A2(new_n453), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT45), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n340), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(KEYINPUT110), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n446), .A2(new_n453), .A3(KEYINPUT45), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n811), .A2(KEYINPUT110), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n663), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT46), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n662), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g632(.A(KEYINPUT111), .B1(new_n816), .B2(new_n817), .ZN(new_n819));
  INV_X1    g633(.A(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n816), .A2(KEYINPUT111), .A3(new_n817), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n818), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n665), .A2(new_n712), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n808), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(new_n818), .ZN(new_n825));
  INV_X1    g639(.A(new_n821), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n825), .B1(new_n826), .B2(new_n819), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n827), .A2(KEYINPUT112), .A3(new_n665), .A4(new_n712), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT44), .ZN(new_n829));
  INV_X1    g643(.A(new_n677), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n801), .A2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT113), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  XOR2_X1   g647(.A(new_n833), .B(KEYINPUT43), .Z(new_n834));
  INV_X1    g648(.A(new_n660), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(new_n700), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n829), .B1(new_n834), .B2(new_n836), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n833), .B(KEYINPUT43), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n838), .A2(KEYINPUT44), .A3(new_n835), .A4(new_n700), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n724), .A2(new_n457), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n837), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n824), .A2(new_n828), .A3(new_n841), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n842), .B(G137), .ZN(G39));
  OAI21_X1  g657(.A(KEYINPUT47), .B1(new_n822), .B2(new_n339), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT47), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n827), .A2(new_n845), .A3(new_n665), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n738), .A2(new_n646), .A3(new_n840), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n844), .A2(new_n611), .A3(new_n846), .A4(new_n847), .ZN(new_n848));
  XNOR2_X1  g662(.A(new_n848), .B(G140), .ZN(G42));
  NAND4_X1  g663(.A1(new_n781), .A2(new_n790), .A3(new_n662), .A4(new_n283), .ZN(new_n850));
  OR2_X1    g664(.A1(new_n834), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n652), .A2(new_n653), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT48), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n853), .B(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n658), .A2(new_n765), .A3(new_n653), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n856), .A2(new_n282), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n838), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n858), .A2(new_n532), .A3(new_n759), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n723), .A2(new_n646), .A3(new_n850), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(new_n678), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n855), .A2(new_n859), .A3(new_n280), .A4(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n860), .A2(new_n801), .A3(new_n677), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n781), .A2(new_n743), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n727), .A2(new_n864), .A3(new_n456), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n865), .B(KEYINPUT120), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n866), .A2(new_n858), .A3(KEYINPUT50), .ZN(new_n867));
  AOI21_X1  g681(.A(KEYINPUT50), .B1(new_n866), .B2(new_n858), .ZN(new_n868));
  OAI221_X1 g682(.A(new_n863), .B1(new_n772), .B2(new_n851), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n844), .A2(new_n846), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n781), .A2(new_n339), .A3(new_n662), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n858), .A2(new_n840), .ZN(new_n873));
  INV_X1    g687(.A(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n869), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n862), .B1(new_n875), .B2(KEYINPUT51), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT54), .ZN(new_n877));
  INV_X1    g691(.A(new_n772), .ZN(new_n878));
  INV_X1    g692(.A(new_n782), .ZN(new_n879));
  AOI22_X1  g693(.A1(new_n878), .A2(new_n879), .B1(new_n652), .B2(new_n709), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n786), .A2(new_n444), .A3(new_n787), .ZN(new_n881));
  NOR4_X1   g695(.A1(new_n642), .A2(new_n698), .A3(new_n339), .A4(new_n706), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n532), .A2(new_n882), .A3(new_n279), .A4(new_n336), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  AOI22_X1  g698(.A1(new_n652), .A2(new_n740), .B1(new_n723), .B2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT52), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n880), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT118), .ZN(new_n888));
  INV_X1    g702(.A(new_n722), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n889), .B1(new_n588), .B2(new_n594), .ZN(new_n890));
  AOI211_X1 g704(.A(new_n457), .B(new_n335), .C1(new_n523), .C2(new_n531), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n788), .A2(new_n891), .A3(new_n279), .A4(new_n882), .ZN(new_n892));
  OAI22_X1  g706(.A1(new_n611), .A2(new_n739), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(new_n708), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n737), .A2(new_n455), .A3(new_n894), .ZN(new_n895));
  OAI22_X1  g709(.A1(new_n611), .A2(new_n895), .B1(new_n772), .B2(new_n782), .ZN(new_n896));
  OAI21_X1  g710(.A(KEYINPUT52), .B1(new_n893), .B2(new_n896), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n887), .A2(new_n888), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n888), .B1(new_n887), .B2(new_n897), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n759), .A2(new_n337), .A3(new_n737), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n767), .A2(new_n759), .A3(new_n679), .ZN(new_n902));
  OAI22_X1  g716(.A1(new_n611), .A2(new_n901), .B1(new_n902), .B2(new_n856), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n681), .A2(new_n653), .A3(new_n759), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n690), .A2(new_n759), .A3(new_n653), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n611), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g720(.A(KEYINPUT114), .B1(new_n903), .B2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT115), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n680), .A2(new_n908), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n678), .A2(new_n532), .A3(KEYINPUT115), .A4(new_n679), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n911), .A2(new_n660), .A3(new_n667), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n328), .A2(new_n330), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n801), .A2(KEYINPUT116), .A3(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT116), .ZN(new_n915));
  INV_X1    g729(.A(new_n913), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n915), .B1(new_n279), .B2(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n688), .B1(new_n914), .B2(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n660), .A2(new_n918), .A3(new_n667), .ZN(new_n919));
  AND3_X1   g733(.A1(new_n912), .A2(new_n701), .A3(new_n919), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n652), .B1(new_n752), .B2(new_n748), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT114), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n921), .A2(new_n760), .A3(new_n770), .A4(new_n922), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n907), .A2(new_n920), .A3(new_n655), .A4(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n806), .B1(new_n795), .B2(new_n796), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n801), .A2(KEYINPUT117), .A3(new_n916), .A4(new_n707), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n724), .A2(new_n457), .A3(new_n699), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT117), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n916), .A2(new_n707), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n928), .B1(new_n279), .B2(new_n929), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n926), .A2(new_n455), .A3(new_n927), .A4(new_n930), .ZN(new_n931));
  OAI22_X1  g745(.A1(new_n611), .A2(new_n931), .B1(new_n772), .B2(new_n791), .ZN(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n925), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n924), .A2(new_n934), .ZN(new_n935));
  XNOR2_X1  g749(.A(KEYINPUT119), .B(KEYINPUT53), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n900), .A2(new_n935), .A3(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT53), .ZN(new_n939));
  AND2_X1   g753(.A1(new_n907), .A2(new_n923), .ZN(new_n940));
  AOI211_X1 g754(.A(new_n932), .B(new_n806), .C1(new_n795), .C2(new_n796), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n912), .A2(new_n701), .A3(new_n919), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n611), .A2(new_n646), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(new_n648), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n852), .A2(KEYINPUT78), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n942), .B1(new_n946), .B2(new_n533), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n940), .A2(new_n941), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n887), .A2(new_n897), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n939), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n877), .B1(new_n938), .B2(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n949), .A2(KEYINPUT118), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n887), .A2(new_n897), .A3(new_n888), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n936), .B1(new_n955), .B2(new_n948), .ZN(new_n956));
  NOR3_X1   g770(.A1(new_n903), .A2(new_n906), .A3(new_n939), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n957), .A2(new_n655), .A3(new_n920), .ZN(new_n958));
  NOR3_X1   g772(.A1(new_n958), .A2(new_n934), .A3(new_n949), .ZN(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n956), .A2(new_n877), .A3(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n876), .A2(new_n952), .A3(new_n961), .ZN(new_n962));
  OAI21_X1  g776(.A(KEYINPUT121), .B1(new_n875), .B2(KEYINPUT51), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT121), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT51), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n873), .B1(new_n870), .B2(new_n871), .ZN(new_n966));
  OAI211_X1 g780(.A(new_n964), .B(new_n965), .C1(new_n966), .C2(new_n869), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n963), .A2(new_n967), .ZN(new_n968));
  OAI22_X1  g782(.A1(new_n962), .A2(new_n968), .B1(G952), .B2(G953), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n781), .A2(new_n662), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n970), .B(KEYINPUT49), .Z(new_n971));
  NOR4_X1   g785(.A1(new_n727), .A2(new_n646), .A3(new_n789), .A4(new_n831), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n971), .A2(new_n890), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n969), .A2(new_n973), .ZN(G75));
  AND4_X1   g788(.A1(new_n655), .A2(new_n907), .A3(new_n920), .A4(new_n923), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n975), .A2(new_n953), .A3(new_n941), .A4(new_n954), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n959), .B1(new_n976), .B2(new_n936), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n977), .A2(new_n287), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n978), .A2(G210), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT56), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n524), .B(new_n527), .Z(new_n981));
  XNOR2_X1  g795(.A(new_n981), .B(KEYINPUT55), .ZN(new_n982));
  AND3_X1   g796(.A1(new_n979), .A2(new_n980), .A3(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n982), .B1(new_n979), .B2(new_n980), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n218), .A2(G952), .ZN(new_n985));
  NOR3_X1   g799(.A1(new_n983), .A2(new_n984), .A3(new_n985), .ZN(G51));
  AOI21_X1  g800(.A(new_n937), .B1(new_n900), .B2(new_n935), .ZN(new_n987));
  OAI21_X1  g801(.A(KEYINPUT54), .B1(new_n987), .B2(new_n959), .ZN(new_n988));
  INV_X1    g802(.A(KEYINPUT122), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n988), .A2(new_n989), .A3(new_n961), .ZN(new_n990));
  OAI211_X1 g804(.A(KEYINPUT122), .B(KEYINPUT54), .C1(new_n987), .C2(new_n959), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n341), .B(KEYINPUT57), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n990), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n993), .A2(new_n661), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n814), .A2(new_n815), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n978), .A2(new_n995), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n985), .B1(new_n994), .B2(new_n996), .ZN(G54));
  AND2_X1   g811(.A1(KEYINPUT58), .A2(G475), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n978), .A2(new_n998), .ZN(new_n999));
  OAI21_X1  g813(.A(KEYINPUT123), .B1(new_n999), .B2(new_n265), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n985), .B1(new_n999), .B2(new_n265), .ZN(new_n1001));
  INV_X1    g815(.A(KEYINPUT123), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n978), .A2(new_n1002), .A3(new_n275), .A4(new_n998), .ZN(new_n1003));
  AND3_X1   g817(.A1(new_n1000), .A2(new_n1001), .A3(new_n1003), .ZN(G60));
  NAND2_X1  g818(.A1(G478), .A2(G902), .ZN(new_n1005));
  XOR2_X1   g819(.A(new_n1005), .B(KEYINPUT59), .Z(new_n1006));
  INV_X1    g820(.A(new_n1006), .ZN(new_n1007));
  NOR3_X1   g821(.A1(new_n987), .A2(KEYINPUT54), .A3(new_n959), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n1007), .B1(new_n1008), .B2(new_n951), .ZN(new_n1009));
  INV_X1    g823(.A(new_n675), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n985), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NAND4_X1  g825(.A1(new_n990), .A2(new_n675), .A3(new_n991), .A4(new_n1007), .ZN(new_n1012));
  AND2_X1   g826(.A1(new_n1011), .A2(new_n1012), .ZN(G63));
  NAND2_X1  g827(.A1(G217), .A2(G902), .ZN(new_n1014));
  XNOR2_X1  g828(.A(new_n1014), .B(KEYINPUT60), .ZN(new_n1015));
  INV_X1    g829(.A(new_n1015), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n1016), .B1(new_n987), .B2(new_n959), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n985), .B1(new_n1017), .B2(new_n639), .ZN(new_n1018));
  INV_X1    g832(.A(KEYINPUT124), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n1015), .B1(new_n956), .B2(new_n960), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n695), .A2(new_n696), .ZN(new_n1021));
  INV_X1    g835(.A(new_n1021), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n1019), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1023));
  NOR4_X1   g837(.A1(new_n977), .A2(KEYINPUT124), .A3(new_n1021), .A4(new_n1015), .ZN(new_n1024));
  OAI21_X1  g838(.A(new_n1018), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g839(.A(KEYINPUT61), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  OAI211_X1 g841(.A(KEYINPUT61), .B(new_n1018), .C1(new_n1023), .C2(new_n1024), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n1027), .A2(new_n1028), .ZN(G66));
  OAI21_X1  g843(.A(G953), .B1(new_n286), .B2(new_n484), .ZN(new_n1030));
  OAI21_X1  g844(.A(new_n1030), .B1(new_n975), .B2(G953), .ZN(new_n1031));
  XNOR2_X1  g845(.A(new_n1031), .B(KEYINPUT125), .ZN(new_n1032));
  INV_X1    g846(.A(G898), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n524), .B1(new_n1033), .B2(G953), .ZN(new_n1034));
  XNOR2_X1  g848(.A(new_n1032), .B(new_n1034), .ZN(G69));
  AOI21_X1  g849(.A(new_n218), .B1(G227), .B2(G900), .ZN(new_n1036));
  OAI21_X1  g850(.A(new_n573), .B1(KEYINPUT30), .B2(new_n555), .ZN(new_n1037));
  XOR2_X1   g851(.A(new_n1037), .B(KEYINPUT126), .Z(new_n1038));
  AND2_X1   g852(.A1(new_n202), .A2(new_n207), .ZN(new_n1039));
  XOR2_X1   g853(.A(new_n1038), .B(new_n1039), .Z(new_n1040));
  AOI21_X1  g854(.A(new_n1040), .B1(G900), .B2(G953), .ZN(new_n1041));
  INV_X1    g855(.A(new_n1041), .ZN(new_n1042));
  NAND4_X1  g856(.A1(new_n824), .A2(new_n828), .A3(new_n943), .A4(new_n767), .ZN(new_n1043));
  NAND3_X1  g857(.A1(new_n1043), .A2(new_n848), .A3(new_n925), .ZN(new_n1044));
  AOI21_X1  g858(.A(new_n896), .B1(new_n652), .B2(new_n740), .ZN(new_n1045));
  AOI21_X1  g859(.A(KEYINPUT127), .B1(new_n842), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g860(.A(new_n1046), .ZN(new_n1047));
  NAND3_X1  g861(.A1(new_n842), .A2(KEYINPUT127), .A3(new_n1045), .ZN(new_n1048));
  AOI21_X1  g862(.A(new_n1044), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g863(.A(new_n1042), .B1(new_n1049), .B2(new_n218), .ZN(new_n1050));
  INV_X1    g864(.A(new_n1040), .ZN(new_n1051));
  OR2_X1    g865(.A1(new_n733), .A2(KEYINPUT105), .ZN(new_n1052));
  NAND2_X1  g866(.A1(new_n733), .A2(KEYINPUT105), .ZN(new_n1053));
  NAND3_X1  g867(.A1(new_n1052), .A2(new_n1053), .A3(new_n1045), .ZN(new_n1054));
  INV_X1    g868(.A(KEYINPUT62), .ZN(new_n1055));
  NAND2_X1  g869(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g870(.A1(new_n735), .A2(KEYINPUT62), .A3(new_n1045), .ZN(new_n1057));
  NAND2_X1  g871(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NOR2_X1   g872(.A1(new_n716), .A2(new_n717), .ZN(new_n1059));
  OAI211_X1 g873(.A(new_n914), .B(new_n917), .C1(new_n801), .C2(new_n677), .ZN(new_n1060));
  NAND4_X1  g874(.A1(new_n946), .A2(new_n1059), .A3(new_n840), .A4(new_n1060), .ZN(new_n1061));
  AND2_X1   g875(.A1(new_n842), .A2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g876(.A1(new_n1058), .A2(new_n1062), .A3(new_n848), .ZN(new_n1063));
  AOI21_X1  g877(.A(new_n1051), .B1(new_n1063), .B2(new_n218), .ZN(new_n1064));
  OAI21_X1  g878(.A(new_n1036), .B1(new_n1050), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g879(.A1(new_n1063), .A2(new_n218), .ZN(new_n1066));
  NAND2_X1  g880(.A1(new_n1066), .A2(new_n1040), .ZN(new_n1067));
  INV_X1    g881(.A(new_n1044), .ZN(new_n1068));
  INV_X1    g882(.A(new_n1048), .ZN(new_n1069));
  OAI211_X1 g883(.A(new_n1068), .B(new_n218), .C1(new_n1046), .C2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g884(.A1(new_n1070), .A2(new_n1041), .ZN(new_n1071));
  INV_X1    g885(.A(new_n1036), .ZN(new_n1072));
  NAND3_X1  g886(.A1(new_n1067), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1073));
  NAND2_X1  g887(.A1(new_n1065), .A2(new_n1073), .ZN(G72));
  INV_X1    g888(.A(new_n595), .ZN(new_n1075));
  NAND2_X1  g889(.A1(new_n1075), .A2(new_n564), .ZN(new_n1076));
  OAI211_X1 g890(.A(new_n1068), .B(new_n975), .C1(new_n1046), .C2(new_n1069), .ZN(new_n1077));
  NAND2_X1  g891(.A1(G472), .A2(G902), .ZN(new_n1078));
  XOR2_X1   g892(.A(new_n1078), .B(KEYINPUT63), .Z(new_n1079));
  AOI21_X1  g893(.A(new_n1076), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1080));
  NAND4_X1  g894(.A1(new_n1058), .A2(new_n1062), .A3(new_n848), .A4(new_n975), .ZN(new_n1081));
  AOI21_X1  g895(.A(new_n719), .B1(new_n1081), .B2(new_n1079), .ZN(new_n1082));
  NOR2_X1   g896(.A1(new_n1075), .A2(new_n563), .ZN(new_n1083));
  INV_X1    g897(.A(new_n578), .ZN(new_n1084));
  OAI21_X1  g898(.A(new_n1079), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g899(.A(new_n1085), .B1(new_n938), .B2(new_n950), .ZN(new_n1086));
  NOR4_X1   g900(.A1(new_n1080), .A2(new_n1082), .A3(new_n985), .A4(new_n1086), .ZN(G57));
endmodule


