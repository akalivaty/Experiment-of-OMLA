

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U547 ( .A1(n720), .A2(n709), .ZN(n512) );
  INV_X1 U548 ( .A(KEYINPUT26), .ZN(n616) );
  XNOR2_X1 U549 ( .A(n617), .B(n616), .ZN(n619) );
  INV_X1 U550 ( .A(KEYINPUT102), .ZN(n621) );
  XNOR2_X1 U551 ( .A(n622), .B(n621), .ZN(n629) );
  NAND2_X1 U552 ( .A1(n671), .A2(n670), .ZN(n715) );
  NAND2_X1 U553 ( .A1(n710), .A2(n512), .ZN(n711) );
  NOR2_X1 U554 ( .A1(G651), .A2(n574), .ZN(n771) );
  XOR2_X1 U555 ( .A(KEYINPUT0), .B(G543), .Z(n574) );
  NAND2_X1 U556 ( .A1(n771), .A2(G47), .ZN(n515) );
  NOR2_X1 U557 ( .A1(G543), .A2(G651), .ZN(n513) );
  XNOR2_X1 U558 ( .A(n513), .B(KEYINPUT64), .ZN(n775) );
  NAND2_X1 U559 ( .A1(G85), .A2(n775), .ZN(n514) );
  NAND2_X1 U560 ( .A1(n515), .A2(n514), .ZN(n519) );
  XNOR2_X1 U561 ( .A(G651), .B(KEYINPUT65), .ZN(n520) );
  NOR2_X1 U562 ( .A1(G543), .A2(n520), .ZN(n516) );
  XOR2_X1 U563 ( .A(KEYINPUT1), .B(n516), .Z(n770) );
  NAND2_X1 U564 ( .A1(n770), .A2(G60), .ZN(n517) );
  XOR2_X1 U565 ( .A(KEYINPUT66), .B(n517), .Z(n518) );
  NOR2_X1 U566 ( .A1(n519), .A2(n518), .ZN(n522) );
  NOR2_X1 U567 ( .A1(n574), .A2(n520), .ZN(n774) );
  NAND2_X1 U568 ( .A1(n774), .A2(G72), .ZN(n521) );
  NAND2_X1 U569 ( .A1(n522), .A2(n521), .ZN(G290) );
  INV_X1 U570 ( .A(G2105), .ZN(n526) );
  AND2_X1 U571 ( .A1(n526), .A2(G2104), .ZN(n876) );
  NAND2_X1 U572 ( .A1(G102), .A2(n876), .ZN(n525) );
  OR2_X1 U573 ( .A1(G2104), .A2(G2105), .ZN(n523) );
  XNOR2_X2 U574 ( .A(KEYINPUT17), .B(n523), .ZN(n877) );
  NAND2_X1 U575 ( .A1(G138), .A2(n877), .ZN(n524) );
  NAND2_X1 U576 ( .A1(n525), .A2(n524), .ZN(n530) );
  NOR2_X1 U577 ( .A1(G2104), .A2(n526), .ZN(n871) );
  NAND2_X1 U578 ( .A1(G126), .A2(n871), .ZN(n528) );
  AND2_X1 U579 ( .A1(G2104), .A2(G2105), .ZN(n872) );
  NAND2_X1 U580 ( .A1(G114), .A2(n872), .ZN(n527) );
  NAND2_X1 U581 ( .A1(n528), .A2(n527), .ZN(n529) );
  NOR2_X1 U582 ( .A1(n530), .A2(n529), .ZN(G164) );
  NAND2_X1 U583 ( .A1(n877), .A2(G137), .ZN(n533) );
  NAND2_X1 U584 ( .A1(G101), .A2(n876), .ZN(n531) );
  XOR2_X1 U585 ( .A(KEYINPUT23), .B(n531), .Z(n532) );
  NAND2_X1 U586 ( .A1(n533), .A2(n532), .ZN(n537) );
  NAND2_X1 U587 ( .A1(G125), .A2(n871), .ZN(n535) );
  NAND2_X1 U588 ( .A1(G113), .A2(n872), .ZN(n534) );
  NAND2_X1 U589 ( .A1(n535), .A2(n534), .ZN(n536) );
  NOR2_X1 U590 ( .A1(n537), .A2(n536), .ZN(G160) );
  NAND2_X1 U591 ( .A1(n770), .A2(G65), .ZN(n539) );
  NAND2_X1 U592 ( .A1(G91), .A2(n775), .ZN(n538) );
  NAND2_X1 U593 ( .A1(n539), .A2(n538), .ZN(n542) );
  NAND2_X1 U594 ( .A1(n771), .A2(G53), .ZN(n540) );
  XOR2_X1 U595 ( .A(KEYINPUT68), .B(n540), .Z(n541) );
  NOR2_X1 U596 ( .A1(n542), .A2(n541), .ZN(n544) );
  NAND2_X1 U597 ( .A1(n774), .A2(G78), .ZN(n543) );
  NAND2_X1 U598 ( .A1(n544), .A2(n543), .ZN(G299) );
  NAND2_X1 U599 ( .A1(G64), .A2(n770), .ZN(n546) );
  NAND2_X1 U600 ( .A1(G52), .A2(n771), .ZN(n545) );
  NAND2_X1 U601 ( .A1(n546), .A2(n545), .ZN(n551) );
  NAND2_X1 U602 ( .A1(G77), .A2(n774), .ZN(n548) );
  NAND2_X1 U603 ( .A1(G90), .A2(n775), .ZN(n547) );
  NAND2_X1 U604 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U605 ( .A(KEYINPUT9), .B(n549), .Z(n550) );
  NOR2_X1 U606 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U607 ( .A(KEYINPUT67), .B(n552), .ZN(G301) );
  INV_X1 U608 ( .A(G301), .ZN(G171) );
  NAND2_X1 U609 ( .A1(G63), .A2(n770), .ZN(n554) );
  NAND2_X1 U610 ( .A1(G51), .A2(n771), .ZN(n553) );
  NAND2_X1 U611 ( .A1(n554), .A2(n553), .ZN(n556) );
  XOR2_X1 U612 ( .A(KEYINPUT6), .B(KEYINPUT75), .Z(n555) );
  XNOR2_X1 U613 ( .A(n556), .B(n555), .ZN(n564) );
  XOR2_X1 U614 ( .A(KEYINPUT4), .B(KEYINPUT74), .Z(n558) );
  NAND2_X1 U615 ( .A1(G89), .A2(n775), .ZN(n557) );
  XNOR2_X1 U616 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U617 ( .A(KEYINPUT73), .B(n559), .ZN(n561) );
  NAND2_X1 U618 ( .A1(G76), .A2(n774), .ZN(n560) );
  NAND2_X1 U619 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U620 ( .A(KEYINPUT5), .B(n562), .Z(n563) );
  NOR2_X1 U621 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U622 ( .A(n565), .B(KEYINPUT7), .Z(n566) );
  XNOR2_X1 U623 ( .A(KEYINPUT76), .B(n566), .ZN(G168) );
  XOR2_X1 U624 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U625 ( .A1(G75), .A2(n774), .ZN(n568) );
  NAND2_X1 U626 ( .A1(G88), .A2(n775), .ZN(n567) );
  NAND2_X1 U627 ( .A1(n568), .A2(n567), .ZN(n572) );
  NAND2_X1 U628 ( .A1(G62), .A2(n770), .ZN(n570) );
  NAND2_X1 U629 ( .A1(G50), .A2(n771), .ZN(n569) );
  NAND2_X1 U630 ( .A1(n570), .A2(n569), .ZN(n571) );
  NOR2_X1 U631 ( .A1(n572), .A2(n571), .ZN(G166) );
  INV_X1 U632 ( .A(G166), .ZN(G303) );
  NAND2_X1 U633 ( .A1(G49), .A2(n771), .ZN(n573) );
  XNOR2_X1 U634 ( .A(n573), .B(KEYINPUT80), .ZN(n579) );
  NAND2_X1 U635 ( .A1(G87), .A2(n574), .ZN(n576) );
  NAND2_X1 U636 ( .A1(G74), .A2(G651), .ZN(n575) );
  NAND2_X1 U637 ( .A1(n576), .A2(n575), .ZN(n577) );
  NOR2_X1 U638 ( .A1(n770), .A2(n577), .ZN(n578) );
  NAND2_X1 U639 ( .A1(n579), .A2(n578), .ZN(G288) );
  NAND2_X1 U640 ( .A1(n775), .A2(G86), .ZN(n580) );
  XNOR2_X1 U641 ( .A(n580), .B(KEYINPUT82), .ZN(n589) );
  NAND2_X1 U642 ( .A1(G73), .A2(n774), .ZN(n581) );
  XOR2_X1 U643 ( .A(KEYINPUT2), .B(n581), .Z(n582) );
  XNOR2_X1 U644 ( .A(n582), .B(KEYINPUT83), .ZN(n584) );
  NAND2_X1 U645 ( .A1(G48), .A2(n771), .ZN(n583) );
  NAND2_X1 U646 ( .A1(n584), .A2(n583), .ZN(n587) );
  NAND2_X1 U647 ( .A1(G61), .A2(n770), .ZN(n585) );
  XNOR2_X1 U648 ( .A(KEYINPUT81), .B(n585), .ZN(n586) );
  NOR2_X1 U649 ( .A1(n587), .A2(n586), .ZN(n588) );
  NAND2_X1 U650 ( .A1(n589), .A2(n588), .ZN(G305) );
  XNOR2_X1 U651 ( .A(G1986), .B(G290), .ZN(n927) );
  NOR2_X1 U652 ( .A1(G164), .A2(G1384), .ZN(n592) );
  NAND2_X1 U653 ( .A1(G160), .A2(G40), .ZN(n590) );
  NOR2_X1 U654 ( .A1(n592), .A2(n590), .ZN(n739) );
  NAND2_X1 U655 ( .A1(n927), .A2(n739), .ZN(n728) );
  XOR2_X1 U656 ( .A(KEYINPUT96), .B(n590), .Z(n591) );
  NAND2_X1 U657 ( .A1(n592), .A2(n591), .ZN(n656) );
  NAND2_X1 U658 ( .A1(G8), .A2(n656), .ZN(n720) );
  INV_X1 U659 ( .A(G299), .ZN(n631) );
  INV_X1 U660 ( .A(KEYINPUT98), .ZN(n593) );
  XNOR2_X1 U661 ( .A(n593), .B(n656), .ZN(n638) );
  NAND2_X1 U662 ( .A1(G2072), .A2(n638), .ZN(n594) );
  XNOR2_X1 U663 ( .A(n594), .B(KEYINPUT27), .ZN(n596) );
  XOR2_X1 U664 ( .A(KEYINPUT100), .B(G1956), .Z(n994) );
  NOR2_X1 U665 ( .A1(n638), .A2(n994), .ZN(n595) );
  NOR2_X1 U666 ( .A1(n596), .A2(n595), .ZN(n630) );
  NOR2_X1 U667 ( .A1(n631), .A2(n630), .ZN(n598) );
  XNOR2_X1 U668 ( .A(KEYINPUT28), .B(KEYINPUT101), .ZN(n597) );
  XNOR2_X1 U669 ( .A(n598), .B(n597), .ZN(n635) );
  NAND2_X1 U670 ( .A1(n770), .A2(G66), .ZN(n600) );
  NAND2_X1 U671 ( .A1(G92), .A2(n775), .ZN(n599) );
  NAND2_X1 U672 ( .A1(n600), .A2(n599), .ZN(n604) );
  NAND2_X1 U673 ( .A1(G79), .A2(n774), .ZN(n602) );
  NAND2_X1 U674 ( .A1(G54), .A2(n771), .ZN(n601) );
  NAND2_X1 U675 ( .A1(n602), .A2(n601), .ZN(n603) );
  NOR2_X1 U676 ( .A1(n604), .A2(n603), .ZN(n606) );
  XNOR2_X1 U677 ( .A(KEYINPUT71), .B(KEYINPUT15), .ZN(n605) );
  XNOR2_X1 U678 ( .A(n606), .B(n605), .ZN(n925) );
  NAND2_X1 U679 ( .A1(n770), .A2(G56), .ZN(n607) );
  XOR2_X1 U680 ( .A(KEYINPUT14), .B(n607), .Z(n613) );
  NAND2_X1 U681 ( .A1(G81), .A2(n775), .ZN(n608) );
  XNOR2_X1 U682 ( .A(n608), .B(KEYINPUT12), .ZN(n610) );
  NAND2_X1 U683 ( .A1(G68), .A2(n774), .ZN(n609) );
  NAND2_X1 U684 ( .A1(n610), .A2(n609), .ZN(n611) );
  XOR2_X1 U685 ( .A(KEYINPUT13), .B(n611), .Z(n612) );
  NOR2_X1 U686 ( .A1(n613), .A2(n612), .ZN(n615) );
  NAND2_X1 U687 ( .A1(n771), .A2(G43), .ZN(n614) );
  NAND2_X1 U688 ( .A1(n615), .A2(n614), .ZN(n942) );
  INV_X1 U689 ( .A(n656), .ZN(n640) );
  AND2_X1 U690 ( .A1(n640), .A2(G1996), .ZN(n617) );
  NAND2_X1 U691 ( .A1(n656), .A2(G1341), .ZN(n618) );
  NAND2_X1 U692 ( .A1(n619), .A2(n618), .ZN(n620) );
  NOR2_X1 U693 ( .A1(n942), .A2(n620), .ZN(n623) );
  NOR2_X1 U694 ( .A1(n925), .A2(n623), .ZN(n622) );
  NAND2_X1 U695 ( .A1(n925), .A2(n623), .ZN(n627) );
  NAND2_X1 U696 ( .A1(G2067), .A2(n638), .ZN(n625) );
  NAND2_X1 U697 ( .A1(G1348), .A2(n656), .ZN(n624) );
  NAND2_X1 U698 ( .A1(n625), .A2(n624), .ZN(n626) );
  NAND2_X1 U699 ( .A1(n627), .A2(n626), .ZN(n628) );
  NAND2_X1 U700 ( .A1(n629), .A2(n628), .ZN(n633) );
  NAND2_X1 U701 ( .A1(n631), .A2(n630), .ZN(n632) );
  NAND2_X1 U702 ( .A1(n633), .A2(n632), .ZN(n634) );
  NAND2_X1 U703 ( .A1(n635), .A2(n634), .ZN(n637) );
  XNOR2_X1 U704 ( .A(KEYINPUT103), .B(KEYINPUT29), .ZN(n636) );
  XNOR2_X1 U705 ( .A(n637), .B(n636), .ZN(n645) );
  INV_X1 U706 ( .A(n638), .ZN(n639) );
  XOR2_X1 U707 ( .A(G2078), .B(KEYINPUT25), .Z(n905) );
  NOR2_X1 U708 ( .A1(n639), .A2(n905), .ZN(n642) );
  NOR2_X1 U709 ( .A1(n640), .A2(G1961), .ZN(n641) );
  NOR2_X1 U710 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U711 ( .A(KEYINPUT99), .B(n643), .ZN(n646) );
  NAND2_X1 U712 ( .A1(n646), .A2(G171), .ZN(n644) );
  NAND2_X1 U713 ( .A1(n645), .A2(n644), .ZN(n655) );
  NOR2_X1 U714 ( .A1(G171), .A2(n646), .ZN(n651) );
  NOR2_X1 U715 ( .A1(G1966), .A2(n720), .ZN(n667) );
  NOR2_X1 U716 ( .A1(G2084), .A2(n656), .ZN(n664) );
  NOR2_X1 U717 ( .A1(n667), .A2(n664), .ZN(n647) );
  NAND2_X1 U718 ( .A1(G8), .A2(n647), .ZN(n648) );
  XNOR2_X1 U719 ( .A(KEYINPUT30), .B(n648), .ZN(n649) );
  NOR2_X1 U720 ( .A1(n649), .A2(G168), .ZN(n650) );
  NOR2_X1 U721 ( .A1(n651), .A2(n650), .ZN(n652) );
  XOR2_X1 U722 ( .A(n652), .B(KEYINPUT31), .Z(n653) );
  XNOR2_X1 U723 ( .A(KEYINPUT104), .B(n653), .ZN(n654) );
  NAND2_X1 U724 ( .A1(n655), .A2(n654), .ZN(n665) );
  NAND2_X1 U725 ( .A1(n665), .A2(G286), .ZN(n661) );
  NOR2_X1 U726 ( .A1(G2090), .A2(n656), .ZN(n658) );
  NOR2_X1 U727 ( .A1(G1971), .A2(n720), .ZN(n657) );
  NOR2_X1 U728 ( .A1(n658), .A2(n657), .ZN(n659) );
  NAND2_X1 U729 ( .A1(n659), .A2(G303), .ZN(n660) );
  NAND2_X1 U730 ( .A1(n661), .A2(n660), .ZN(n662) );
  NAND2_X1 U731 ( .A1(n662), .A2(G8), .ZN(n663) );
  XNOR2_X1 U732 ( .A(KEYINPUT32), .B(n663), .ZN(n671) );
  NAND2_X1 U733 ( .A1(G8), .A2(n664), .ZN(n669) );
  INV_X1 U734 ( .A(n665), .ZN(n666) );
  NOR2_X1 U735 ( .A1(n667), .A2(n666), .ZN(n668) );
  NAND2_X1 U736 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U737 ( .A1(G1976), .A2(G288), .ZN(n708) );
  NOR2_X1 U738 ( .A1(G1971), .A2(G303), .ZN(n672) );
  NOR2_X1 U739 ( .A1(n708), .A2(n672), .ZN(n936) );
  NAND2_X1 U740 ( .A1(n715), .A2(n936), .ZN(n673) );
  NAND2_X1 U741 ( .A1(G1976), .A2(G288), .ZN(n932) );
  NAND2_X1 U742 ( .A1(n673), .A2(n932), .ZN(n674) );
  NOR2_X1 U743 ( .A1(n720), .A2(n674), .ZN(n675) );
  NOR2_X1 U744 ( .A1(KEYINPUT33), .A2(n675), .ZN(n712) );
  XOR2_X1 U745 ( .A(G1981), .B(G305), .Z(n928) );
  NAND2_X1 U746 ( .A1(G105), .A2(n876), .ZN(n676) );
  XOR2_X1 U747 ( .A(KEYINPUT38), .B(n676), .Z(n682) );
  NAND2_X1 U748 ( .A1(n871), .A2(G129), .ZN(n677) );
  XOR2_X1 U749 ( .A(KEYINPUT91), .B(n677), .Z(n679) );
  NAND2_X1 U750 ( .A1(n872), .A2(G117), .ZN(n678) );
  NAND2_X1 U751 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U752 ( .A(KEYINPUT92), .B(n680), .ZN(n681) );
  NOR2_X1 U753 ( .A1(n682), .A2(n681), .ZN(n684) );
  NAND2_X1 U754 ( .A1(n877), .A2(G141), .ZN(n683) );
  NAND2_X1 U755 ( .A1(n684), .A2(n683), .ZN(n883) );
  NAND2_X1 U756 ( .A1(G1996), .A2(n883), .ZN(n685) );
  XNOR2_X1 U757 ( .A(KEYINPUT93), .B(n685), .ZN(n694) );
  NAND2_X1 U758 ( .A1(G119), .A2(n871), .ZN(n687) );
  NAND2_X1 U759 ( .A1(G131), .A2(n877), .ZN(n686) );
  NAND2_X1 U760 ( .A1(n687), .A2(n686), .ZN(n691) );
  NAND2_X1 U761 ( .A1(G107), .A2(n872), .ZN(n689) );
  NAND2_X1 U762 ( .A1(G95), .A2(n876), .ZN(n688) );
  NAND2_X1 U763 ( .A1(n689), .A2(n688), .ZN(n690) );
  OR2_X1 U764 ( .A1(n691), .A2(n690), .ZN(n868) );
  NAND2_X1 U765 ( .A1(G1991), .A2(n868), .ZN(n692) );
  XOR2_X1 U766 ( .A(KEYINPUT90), .B(n692), .Z(n693) );
  NOR2_X1 U767 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U768 ( .A(KEYINPUT94), .B(n695), .ZN(n961) );
  XNOR2_X1 U769 ( .A(KEYINPUT95), .B(n739), .ZN(n696) );
  NOR2_X1 U770 ( .A1(n961), .A2(n696), .ZN(n731) );
  INV_X1 U771 ( .A(n731), .ZN(n707) );
  XNOR2_X1 U772 ( .A(G2067), .B(KEYINPUT37), .ZN(n736) );
  NAND2_X1 U773 ( .A1(G104), .A2(n876), .ZN(n698) );
  NAND2_X1 U774 ( .A1(G140), .A2(n877), .ZN(n697) );
  NAND2_X1 U775 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U776 ( .A(KEYINPUT34), .B(n699), .ZN(n704) );
  NAND2_X1 U777 ( .A1(G128), .A2(n871), .ZN(n701) );
  NAND2_X1 U778 ( .A1(G116), .A2(n872), .ZN(n700) );
  NAND2_X1 U779 ( .A1(n701), .A2(n700), .ZN(n702) );
  XOR2_X1 U780 ( .A(n702), .B(KEYINPUT35), .Z(n703) );
  NOR2_X1 U781 ( .A1(n704), .A2(n703), .ZN(n705) );
  XOR2_X1 U782 ( .A(KEYINPUT36), .B(n705), .Z(n706) );
  XNOR2_X1 U783 ( .A(KEYINPUT89), .B(n706), .ZN(n886) );
  NOR2_X1 U784 ( .A1(n736), .A2(n886), .ZN(n964) );
  NAND2_X1 U785 ( .A1(n739), .A2(n964), .ZN(n734) );
  AND2_X1 U786 ( .A1(n707), .A2(n734), .ZN(n724) );
  AND2_X1 U787 ( .A1(n928), .A2(n724), .ZN(n710) );
  NAND2_X1 U788 ( .A1(n708), .A2(KEYINPUT33), .ZN(n709) );
  NOR2_X1 U789 ( .A1(n712), .A2(n711), .ZN(n726) );
  NOR2_X1 U790 ( .A1(G2090), .A2(G303), .ZN(n713) );
  NAND2_X1 U791 ( .A1(G8), .A2(n713), .ZN(n714) );
  NAND2_X1 U792 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U793 ( .A1(n716), .A2(n720), .ZN(n722) );
  NOR2_X1 U794 ( .A1(G1981), .A2(G305), .ZN(n717) );
  XNOR2_X1 U795 ( .A(n717), .B(KEYINPUT97), .ZN(n718) );
  XNOR2_X1 U796 ( .A(KEYINPUT24), .B(n718), .ZN(n719) );
  OR2_X1 U797 ( .A1(n720), .A2(n719), .ZN(n721) );
  NAND2_X1 U798 ( .A1(n722), .A2(n721), .ZN(n723) );
  AND2_X1 U799 ( .A1(n724), .A2(n723), .ZN(n725) );
  OR2_X1 U800 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U801 ( .A1(n728), .A2(n727), .ZN(n742) );
  NOR2_X1 U802 ( .A1(G1996), .A2(n883), .ZN(n957) );
  NOR2_X1 U803 ( .A1(G1986), .A2(G290), .ZN(n729) );
  NOR2_X1 U804 ( .A1(G1991), .A2(n868), .ZN(n966) );
  NOR2_X1 U805 ( .A1(n729), .A2(n966), .ZN(n730) );
  NOR2_X1 U806 ( .A1(n731), .A2(n730), .ZN(n732) );
  NOR2_X1 U807 ( .A1(n957), .A2(n732), .ZN(n733) );
  XNOR2_X1 U808 ( .A(KEYINPUT39), .B(n733), .ZN(n735) );
  NAND2_X1 U809 ( .A1(n735), .A2(n734), .ZN(n737) );
  NAND2_X1 U810 ( .A1(n736), .A2(n886), .ZN(n970) );
  NAND2_X1 U811 ( .A1(n737), .A2(n970), .ZN(n738) );
  NAND2_X1 U812 ( .A1(n739), .A2(n738), .ZN(n740) );
  XOR2_X1 U813 ( .A(KEYINPUT105), .B(n740), .Z(n741) );
  NAND2_X1 U814 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U815 ( .A(n743), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U816 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U817 ( .A(G132), .ZN(G219) );
  INV_X1 U818 ( .A(G82), .ZN(G220) );
  INV_X1 U819 ( .A(G57), .ZN(G237) );
  XOR2_X1 U820 ( .A(KEYINPUT10), .B(KEYINPUT69), .Z(n745) );
  NAND2_X1 U821 ( .A1(G7), .A2(G661), .ZN(n744) );
  XNOR2_X1 U822 ( .A(n745), .B(n744), .ZN(G223) );
  INV_X1 U823 ( .A(G223), .ZN(n821) );
  NAND2_X1 U824 ( .A1(n821), .A2(G567), .ZN(n746) );
  XOR2_X1 U825 ( .A(KEYINPUT11), .B(n746), .Z(G234) );
  INV_X1 U826 ( .A(G860), .ZN(n755) );
  OR2_X1 U827 ( .A1(n942), .A2(n755), .ZN(n747) );
  XNOR2_X1 U828 ( .A(KEYINPUT70), .B(n747), .ZN(G153) );
  NAND2_X1 U829 ( .A1(G171), .A2(G868), .ZN(n750) );
  INV_X1 U830 ( .A(G868), .ZN(n748) );
  NAND2_X1 U831 ( .A1(n925), .A2(n748), .ZN(n749) );
  NAND2_X1 U832 ( .A1(n750), .A2(n749), .ZN(n751) );
  XOR2_X1 U833 ( .A(KEYINPUT72), .B(n751), .Z(G284) );
  XNOR2_X1 U834 ( .A(KEYINPUT77), .B(G868), .ZN(n752) );
  NOR2_X1 U835 ( .A1(G286), .A2(n752), .ZN(n754) );
  NOR2_X1 U836 ( .A1(G868), .A2(G299), .ZN(n753) );
  NOR2_X1 U837 ( .A1(n754), .A2(n753), .ZN(G297) );
  NAND2_X1 U838 ( .A1(n755), .A2(G559), .ZN(n756) );
  NAND2_X1 U839 ( .A1(n756), .A2(n925), .ZN(n757) );
  XNOR2_X1 U840 ( .A(n757), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U841 ( .A1(G868), .A2(n942), .ZN(n760) );
  NAND2_X1 U842 ( .A1(G868), .A2(n925), .ZN(n758) );
  NOR2_X1 U843 ( .A1(G559), .A2(n758), .ZN(n759) );
  NOR2_X1 U844 ( .A1(n760), .A2(n759), .ZN(G282) );
  NAND2_X1 U845 ( .A1(n871), .A2(G123), .ZN(n761) );
  XNOR2_X1 U846 ( .A(n761), .B(KEYINPUT18), .ZN(n763) );
  NAND2_X1 U847 ( .A1(G111), .A2(n872), .ZN(n762) );
  NAND2_X1 U848 ( .A1(n763), .A2(n762), .ZN(n767) );
  NAND2_X1 U849 ( .A1(G99), .A2(n876), .ZN(n765) );
  NAND2_X1 U850 ( .A1(G135), .A2(n877), .ZN(n764) );
  NAND2_X1 U851 ( .A1(n765), .A2(n764), .ZN(n766) );
  NOR2_X1 U852 ( .A1(n767), .A2(n766), .ZN(n965) );
  XNOR2_X1 U853 ( .A(n965), .B(G2096), .ZN(n769) );
  INV_X1 U854 ( .A(G2100), .ZN(n768) );
  NAND2_X1 U855 ( .A1(n769), .A2(n768), .ZN(G156) );
  NAND2_X1 U856 ( .A1(G67), .A2(n770), .ZN(n773) );
  NAND2_X1 U857 ( .A1(G55), .A2(n771), .ZN(n772) );
  NAND2_X1 U858 ( .A1(n773), .A2(n772), .ZN(n779) );
  NAND2_X1 U859 ( .A1(G80), .A2(n774), .ZN(n777) );
  NAND2_X1 U860 ( .A1(G93), .A2(n775), .ZN(n776) );
  NAND2_X1 U861 ( .A1(n777), .A2(n776), .ZN(n778) );
  NOR2_X1 U862 ( .A1(n779), .A2(n778), .ZN(n792) );
  NAND2_X1 U863 ( .A1(G559), .A2(n925), .ZN(n780) );
  XOR2_X1 U864 ( .A(n942), .B(n780), .Z(n789) );
  XOR2_X1 U865 ( .A(n789), .B(KEYINPUT78), .Z(n781) );
  NOR2_X1 U866 ( .A1(G860), .A2(n781), .ZN(n782) );
  XOR2_X1 U867 ( .A(KEYINPUT79), .B(n782), .Z(n783) );
  XNOR2_X1 U868 ( .A(n792), .B(n783), .ZN(G145) );
  XNOR2_X1 U869 ( .A(KEYINPUT19), .B(G288), .ZN(n788) );
  XNOR2_X1 U870 ( .A(G166), .B(n792), .ZN(n786) );
  XNOR2_X1 U871 ( .A(G299), .B(G305), .ZN(n784) );
  XNOR2_X1 U872 ( .A(n784), .B(G290), .ZN(n785) );
  XNOR2_X1 U873 ( .A(n786), .B(n785), .ZN(n787) );
  XNOR2_X1 U874 ( .A(n788), .B(n787), .ZN(n890) );
  XNOR2_X1 U875 ( .A(n890), .B(n789), .ZN(n790) );
  NAND2_X1 U876 ( .A1(n790), .A2(G868), .ZN(n791) );
  XNOR2_X1 U877 ( .A(n791), .B(KEYINPUT84), .ZN(n794) );
  OR2_X1 U878 ( .A1(G868), .A2(n792), .ZN(n793) );
  NAND2_X1 U879 ( .A1(n794), .A2(n793), .ZN(G295) );
  NAND2_X1 U880 ( .A1(G2078), .A2(G2084), .ZN(n797) );
  XNOR2_X1 U881 ( .A(KEYINPUT85), .B(KEYINPUT20), .ZN(n795) );
  XNOR2_X1 U882 ( .A(n795), .B(KEYINPUT86), .ZN(n796) );
  XNOR2_X1 U883 ( .A(n797), .B(n796), .ZN(n798) );
  NAND2_X1 U884 ( .A1(n798), .A2(G2090), .ZN(n800) );
  XOR2_X1 U885 ( .A(KEYINPUT87), .B(KEYINPUT21), .Z(n799) );
  XNOR2_X1 U886 ( .A(n800), .B(n799), .ZN(n801) );
  NAND2_X1 U887 ( .A1(G2072), .A2(n801), .ZN(G158) );
  XNOR2_X1 U888 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U889 ( .A1(G120), .A2(G69), .ZN(n802) );
  NOR2_X1 U890 ( .A1(G237), .A2(n802), .ZN(n803) );
  XNOR2_X1 U891 ( .A(KEYINPUT88), .B(n803), .ZN(n804) );
  NAND2_X1 U892 ( .A1(n804), .A2(G108), .ZN(n827) );
  NAND2_X1 U893 ( .A1(n827), .A2(G567), .ZN(n809) );
  NOR2_X1 U894 ( .A1(G220), .A2(G219), .ZN(n805) );
  XOR2_X1 U895 ( .A(KEYINPUT22), .B(n805), .Z(n806) );
  NOR2_X1 U896 ( .A1(G218), .A2(n806), .ZN(n807) );
  NAND2_X1 U897 ( .A1(G96), .A2(n807), .ZN(n828) );
  NAND2_X1 U898 ( .A1(n828), .A2(G2106), .ZN(n808) );
  NAND2_X1 U899 ( .A1(n809), .A2(n808), .ZN(n829) );
  NAND2_X1 U900 ( .A1(G483), .A2(G661), .ZN(n810) );
  NOR2_X1 U901 ( .A1(n829), .A2(n810), .ZN(n824) );
  NAND2_X1 U902 ( .A1(n824), .A2(G36), .ZN(G176) );
  XNOR2_X1 U903 ( .A(G2430), .B(G2454), .ZN(n819) );
  XNOR2_X1 U904 ( .A(KEYINPUT106), .B(G2435), .ZN(n817) );
  XOR2_X1 U905 ( .A(G2451), .B(G2427), .Z(n812) );
  XNOR2_X1 U906 ( .A(G2438), .B(G2446), .ZN(n811) );
  XNOR2_X1 U907 ( .A(n812), .B(n811), .ZN(n813) );
  XOR2_X1 U908 ( .A(n813), .B(G2443), .Z(n815) );
  XNOR2_X1 U909 ( .A(G1341), .B(G1348), .ZN(n814) );
  XNOR2_X1 U910 ( .A(n815), .B(n814), .ZN(n816) );
  XNOR2_X1 U911 ( .A(n817), .B(n816), .ZN(n818) );
  XNOR2_X1 U912 ( .A(n819), .B(n818), .ZN(n820) );
  NAND2_X1 U913 ( .A1(n820), .A2(G14), .ZN(n895) );
  XNOR2_X1 U914 ( .A(KEYINPUT107), .B(n895), .ZN(G401) );
  NAND2_X1 U915 ( .A1(G2106), .A2(n821), .ZN(G217) );
  AND2_X1 U916 ( .A1(G15), .A2(G2), .ZN(n822) );
  NAND2_X1 U917 ( .A1(G661), .A2(n822), .ZN(G259) );
  NAND2_X1 U918 ( .A1(G3), .A2(G1), .ZN(n823) );
  XNOR2_X1 U919 ( .A(KEYINPUT108), .B(n823), .ZN(n825) );
  NAND2_X1 U920 ( .A1(n825), .A2(n824), .ZN(n826) );
  XOR2_X1 U921 ( .A(KEYINPUT109), .B(n826), .Z(G188) );
  NOR2_X1 U922 ( .A1(n828), .A2(n827), .ZN(G325) );
  XOR2_X1 U923 ( .A(KEYINPUT110), .B(G325), .Z(G261) );
  INV_X1 U925 ( .A(G120), .ZN(G236) );
  INV_X1 U926 ( .A(G108), .ZN(G238) );
  INV_X1 U927 ( .A(G96), .ZN(G221) );
  INV_X1 U928 ( .A(G69), .ZN(G235) );
  INV_X1 U929 ( .A(n829), .ZN(G319) );
  XOR2_X1 U930 ( .A(KEYINPUT111), .B(G2090), .Z(n831) );
  XNOR2_X1 U931 ( .A(G2078), .B(G2072), .ZN(n830) );
  XNOR2_X1 U932 ( .A(n831), .B(n830), .ZN(n832) );
  XOR2_X1 U933 ( .A(n832), .B(G2100), .Z(n834) );
  XNOR2_X1 U934 ( .A(G2067), .B(G2084), .ZN(n833) );
  XNOR2_X1 U935 ( .A(n834), .B(n833), .ZN(n838) );
  XOR2_X1 U936 ( .A(G2096), .B(G2678), .Z(n836) );
  XNOR2_X1 U937 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n835) );
  XNOR2_X1 U938 ( .A(n836), .B(n835), .ZN(n837) );
  XOR2_X1 U939 ( .A(n838), .B(n837), .Z(G227) );
  XOR2_X1 U940 ( .A(G1976), .B(G1981), .Z(n840) );
  XNOR2_X1 U941 ( .A(G1966), .B(G1961), .ZN(n839) );
  XNOR2_X1 U942 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U943 ( .A(n841), .B(KEYINPUT41), .Z(n843) );
  XNOR2_X1 U944 ( .A(G1971), .B(G1986), .ZN(n842) );
  XNOR2_X1 U945 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U946 ( .A(G2474), .B(G1956), .Z(n845) );
  XNOR2_X1 U947 ( .A(G1996), .B(G1991), .ZN(n844) );
  XNOR2_X1 U948 ( .A(n845), .B(n844), .ZN(n846) );
  XNOR2_X1 U949 ( .A(n847), .B(n846), .ZN(G229) );
  NAND2_X1 U950 ( .A1(n871), .A2(G124), .ZN(n848) );
  XNOR2_X1 U951 ( .A(n848), .B(KEYINPUT44), .ZN(n850) );
  NAND2_X1 U952 ( .A1(G112), .A2(n872), .ZN(n849) );
  NAND2_X1 U953 ( .A1(n850), .A2(n849), .ZN(n854) );
  NAND2_X1 U954 ( .A1(G100), .A2(n876), .ZN(n852) );
  NAND2_X1 U955 ( .A1(G136), .A2(n877), .ZN(n851) );
  NAND2_X1 U956 ( .A1(n852), .A2(n851), .ZN(n853) );
  NOR2_X1 U957 ( .A1(n854), .A2(n853), .ZN(G162) );
  XOR2_X1 U958 ( .A(KEYINPUT114), .B(KEYINPUT113), .Z(n856) );
  XNOR2_X1 U959 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n855) );
  XNOR2_X1 U960 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U961 ( .A(G162), .B(n965), .Z(n858) );
  XNOR2_X1 U962 ( .A(G164), .B(G160), .ZN(n857) );
  XNOR2_X1 U963 ( .A(n858), .B(n857), .ZN(n859) );
  XNOR2_X1 U964 ( .A(n860), .B(n859), .ZN(n870) );
  NAND2_X1 U965 ( .A1(G103), .A2(n876), .ZN(n862) );
  NAND2_X1 U966 ( .A1(G139), .A2(n877), .ZN(n861) );
  NAND2_X1 U967 ( .A1(n862), .A2(n861), .ZN(n867) );
  NAND2_X1 U968 ( .A1(G127), .A2(n871), .ZN(n864) );
  NAND2_X1 U969 ( .A1(G115), .A2(n872), .ZN(n863) );
  NAND2_X1 U970 ( .A1(n864), .A2(n863), .ZN(n865) );
  XOR2_X1 U971 ( .A(KEYINPUT47), .B(n865), .Z(n866) );
  NOR2_X1 U972 ( .A1(n867), .A2(n866), .ZN(n952) );
  XNOR2_X1 U973 ( .A(n868), .B(n952), .ZN(n869) );
  XNOR2_X1 U974 ( .A(n870), .B(n869), .ZN(n888) );
  NAND2_X1 U975 ( .A1(G130), .A2(n871), .ZN(n874) );
  NAND2_X1 U976 ( .A1(G118), .A2(n872), .ZN(n873) );
  NAND2_X1 U977 ( .A1(n874), .A2(n873), .ZN(n875) );
  XNOR2_X1 U978 ( .A(KEYINPUT112), .B(n875), .ZN(n882) );
  NAND2_X1 U979 ( .A1(G106), .A2(n876), .ZN(n879) );
  NAND2_X1 U980 ( .A1(G142), .A2(n877), .ZN(n878) );
  NAND2_X1 U981 ( .A1(n879), .A2(n878), .ZN(n880) );
  XOR2_X1 U982 ( .A(n880), .B(KEYINPUT45), .Z(n881) );
  NOR2_X1 U983 ( .A1(n882), .A2(n881), .ZN(n884) );
  XNOR2_X1 U984 ( .A(n884), .B(n883), .ZN(n885) );
  XOR2_X1 U985 ( .A(n886), .B(n885), .Z(n887) );
  XNOR2_X1 U986 ( .A(n888), .B(n887), .ZN(n889) );
  NOR2_X1 U987 ( .A1(G37), .A2(n889), .ZN(G395) );
  XNOR2_X1 U988 ( .A(G286), .B(n890), .ZN(n892) );
  XNOR2_X1 U989 ( .A(G171), .B(n925), .ZN(n891) );
  XNOR2_X1 U990 ( .A(n892), .B(n891), .ZN(n893) );
  XNOR2_X1 U991 ( .A(n893), .B(n942), .ZN(n894) );
  NOR2_X1 U992 ( .A1(G37), .A2(n894), .ZN(G397) );
  NAND2_X1 U993 ( .A1(G319), .A2(n895), .ZN(n898) );
  NOR2_X1 U994 ( .A1(G227), .A2(G229), .ZN(n896) );
  XNOR2_X1 U995 ( .A(KEYINPUT49), .B(n896), .ZN(n897) );
  NOR2_X1 U996 ( .A1(n898), .A2(n897), .ZN(n900) );
  NOR2_X1 U997 ( .A1(G395), .A2(G397), .ZN(n899) );
  NAND2_X1 U998 ( .A1(n900), .A2(n899), .ZN(G225) );
  INV_X1 U999 ( .A(G225), .ZN(G308) );
  XOR2_X1 U1000 ( .A(G2090), .B(G35), .Z(n916) );
  XOR2_X1 U1001 ( .A(G2067), .B(G26), .Z(n901) );
  XNOR2_X1 U1002 ( .A(KEYINPUT117), .B(n901), .ZN(n903) );
  XNOR2_X1 U1003 ( .A(G33), .B(G2072), .ZN(n902) );
  NOR2_X1 U1004 ( .A1(n903), .A2(n902), .ZN(n904) );
  XNOR2_X1 U1005 ( .A(KEYINPUT118), .B(n904), .ZN(n909) );
  XNOR2_X1 U1006 ( .A(G1996), .B(G32), .ZN(n907) );
  XNOR2_X1 U1007 ( .A(n905), .B(G27), .ZN(n906) );
  NOR2_X1 U1008 ( .A1(n907), .A2(n906), .ZN(n908) );
  NAND2_X1 U1009 ( .A1(n909), .A2(n908), .ZN(n912) );
  XOR2_X1 U1010 ( .A(G1991), .B(G25), .Z(n910) );
  NAND2_X1 U1011 ( .A1(n910), .A2(G28), .ZN(n911) );
  NOR2_X1 U1012 ( .A1(n912), .A2(n911), .ZN(n913) );
  XNOR2_X1 U1013 ( .A(n913), .B(KEYINPUT53), .ZN(n914) );
  XNOR2_X1 U1014 ( .A(n914), .B(KEYINPUT119), .ZN(n915) );
  NAND2_X1 U1015 ( .A1(n916), .A2(n915), .ZN(n919) );
  XNOR2_X1 U1016 ( .A(G34), .B(G2084), .ZN(n917) );
  XNOR2_X1 U1017 ( .A(KEYINPUT54), .B(n917), .ZN(n918) );
  NOR2_X1 U1018 ( .A1(n919), .A2(n918), .ZN(n921) );
  XOR2_X1 U1019 ( .A(KEYINPUT55), .B(KEYINPUT116), .Z(n975) );
  XOR2_X1 U1020 ( .A(KEYINPUT120), .B(n975), .Z(n920) );
  XNOR2_X1 U1021 ( .A(n921), .B(n920), .ZN(n923) );
  INV_X1 U1022 ( .A(G29), .ZN(n922) );
  NAND2_X1 U1023 ( .A1(n923), .A2(n922), .ZN(n924) );
  NAND2_X1 U1024 ( .A1(n924), .A2(G11), .ZN(n951) );
  XNOR2_X1 U1025 ( .A(KEYINPUT56), .B(G16), .ZN(n948) );
  XOR2_X1 U1026 ( .A(n925), .B(G1348), .Z(n926) );
  NOR2_X1 U1027 ( .A1(n927), .A2(n926), .ZN(n946) );
  XNOR2_X1 U1028 ( .A(G1966), .B(G168), .ZN(n929) );
  NAND2_X1 U1029 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1030 ( .A(KEYINPUT57), .B(n930), .ZN(n941) );
  NAND2_X1 U1031 ( .A1(G1971), .A2(G303), .ZN(n931) );
  NAND2_X1 U1032 ( .A1(n932), .A2(n931), .ZN(n934) );
  XNOR2_X1 U1033 ( .A(G1961), .B(G301), .ZN(n933) );
  NOR2_X1 U1034 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1035 ( .A1(n936), .A2(n935), .ZN(n939) );
  XOR2_X1 U1036 ( .A(G1956), .B(G299), .Z(n937) );
  XNOR2_X1 U1037 ( .A(KEYINPUT121), .B(n937), .ZN(n938) );
  NOR2_X1 U1038 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1039 ( .A1(n941), .A2(n940), .ZN(n944) );
  XNOR2_X1 U1040 ( .A(G1341), .B(n942), .ZN(n943) );
  NOR2_X1 U1041 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1042 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1043 ( .A1(n948), .A2(n947), .ZN(n949) );
  XOR2_X1 U1044 ( .A(KEYINPUT122), .B(n949), .Z(n950) );
  NOR2_X1 U1045 ( .A1(n951), .A2(n950), .ZN(n979) );
  XOR2_X1 U1046 ( .A(G2072), .B(n952), .Z(n954) );
  XOR2_X1 U1047 ( .A(G164), .B(G2078), .Z(n953) );
  NOR2_X1 U1048 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1049 ( .A(KEYINPUT50), .B(n955), .ZN(n960) );
  XOR2_X1 U1050 ( .A(G2090), .B(G162), .Z(n956) );
  NOR2_X1 U1051 ( .A1(n957), .A2(n956), .ZN(n958) );
  XOR2_X1 U1052 ( .A(KEYINPUT51), .B(n958), .Z(n959) );
  NAND2_X1 U1053 ( .A1(n960), .A2(n959), .ZN(n973) );
  XNOR2_X1 U1054 ( .A(G2084), .B(G160), .ZN(n962) );
  NAND2_X1 U1055 ( .A1(n962), .A2(n961), .ZN(n963) );
  NOR2_X1 U1056 ( .A1(n964), .A2(n963), .ZN(n968) );
  NOR2_X1 U1057 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1058 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1059 ( .A(KEYINPUT115), .B(n969), .ZN(n971) );
  NAND2_X1 U1060 ( .A1(n971), .A2(n970), .ZN(n972) );
  NOR2_X1 U1061 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1062 ( .A(KEYINPUT52), .B(n974), .ZN(n976) );
  NAND2_X1 U1063 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1064 ( .A1(n977), .A2(G29), .ZN(n978) );
  NAND2_X1 U1065 ( .A1(n979), .A2(n978), .ZN(n1008) );
  XOR2_X1 U1066 ( .A(G1986), .B(G24), .Z(n983) );
  XNOR2_X1 U1067 ( .A(G1971), .B(G22), .ZN(n981) );
  XNOR2_X1 U1068 ( .A(G23), .B(G1976), .ZN(n980) );
  NOR2_X1 U1069 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1070 ( .A1(n983), .A2(n982), .ZN(n985) );
  XNOR2_X1 U1071 ( .A(KEYINPUT125), .B(KEYINPUT58), .ZN(n984) );
  XNOR2_X1 U1072 ( .A(n985), .B(n984), .ZN(n989) );
  XNOR2_X1 U1073 ( .A(G1966), .B(G21), .ZN(n987) );
  XNOR2_X1 U1074 ( .A(G5), .B(G1961), .ZN(n986) );
  NOR2_X1 U1075 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1076 ( .A1(n989), .A2(n988), .ZN(n1002) );
  XOR2_X1 U1077 ( .A(G1981), .B(G6), .Z(n990) );
  XNOR2_X1 U1078 ( .A(KEYINPUT123), .B(n990), .ZN(n992) );
  XNOR2_X1 U1079 ( .A(G19), .B(G1341), .ZN(n991) );
  NOR2_X1 U1080 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1081 ( .A(KEYINPUT124), .B(n993), .ZN(n996) );
  XNOR2_X1 U1082 ( .A(n994), .B(G20), .ZN(n995) );
  NAND2_X1 U1083 ( .A1(n996), .A2(n995), .ZN(n999) );
  XOR2_X1 U1084 ( .A(KEYINPUT59), .B(G1348), .Z(n997) );
  XNOR2_X1 U1085 ( .A(G4), .B(n997), .ZN(n998) );
  NOR2_X1 U1086 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XOR2_X1 U1087 ( .A(n1000), .B(KEYINPUT60), .Z(n1001) );
  NOR2_X1 U1088 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XOR2_X1 U1089 ( .A(KEYINPUT127), .B(n1003), .Z(n1005) );
  XOR2_X1 U1090 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n1004) );
  XNOR2_X1 U1091 ( .A(n1005), .B(n1004), .ZN(n1006) );
  NOR2_X1 U1092 ( .A1(G16), .A2(n1006), .ZN(n1007) );
  NOR2_X1 U1093 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1094 ( .A(n1009), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1095 ( .A(G311), .ZN(G150) );
endmodule

