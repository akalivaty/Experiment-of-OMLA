//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 1 1 1 0 0 1 1 1 1 0 0 0 1 1 0 0 1 1 0 1 1 0 1 1 0 1 1 1 1 1 0 1 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:23 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n599, new_n601, new_n602, new_n603,
    new_n604, new_n605, new_n606, new_n607, new_n608, new_n609, new_n610,
    new_n611, new_n612, new_n613, new_n614, new_n615, new_n616, new_n617,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n850, new_n851, new_n852, new_n853, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT72), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT71), .ZN(new_n189));
  INV_X1    g003(.A(G131), .ZN(new_n190));
  INV_X1    g004(.A(G137), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G134), .ZN(new_n192));
  INV_X1    g006(.A(G134), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G137), .ZN(new_n194));
  AOI21_X1  g008(.A(new_n190), .B1(new_n192), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT11), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n197), .B1(new_n193), .B2(G137), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n191), .A2(KEYINPUT11), .A3(G134), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n198), .A2(new_n199), .A3(new_n190), .A4(new_n194), .ZN(new_n200));
  AND2_X1   g014(.A1(new_n200), .A2(KEYINPUT64), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n200), .A2(KEYINPUT64), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n196), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT67), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  XNOR2_X1  g019(.A(G143), .B(G146), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT1), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n206), .A2(new_n207), .A3(G128), .ZN(new_n208));
  INV_X1    g022(.A(G128), .ZN(new_n209));
  INV_X1    g023(.A(G146), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n209), .A2(new_n210), .A3(G143), .ZN(new_n211));
  INV_X1    g025(.A(G143), .ZN(new_n212));
  OAI211_X1 g026(.A(new_n212), .B(G146), .C1(new_n209), .C2(KEYINPUT1), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n208), .A2(new_n211), .A3(new_n213), .ZN(new_n214));
  AOI21_X1  g028(.A(KEYINPUT11), .B1(new_n191), .B2(G134), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n191), .A2(G134), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT64), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n217), .A2(new_n218), .A3(new_n190), .A4(new_n199), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n200), .A2(KEYINPUT64), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n221), .A2(KEYINPUT67), .A3(new_n196), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n205), .A2(new_n214), .A3(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT66), .ZN(new_n224));
  INV_X1    g038(.A(G113), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(KEYINPUT2), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT2), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G113), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  XNOR2_X1  g043(.A(G116), .B(G119), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n229), .A2(new_n230), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n224), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  OR2_X1    g048(.A1(new_n229), .A2(new_n230), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n235), .A2(KEYINPUT66), .A3(new_n231), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n198), .A2(new_n199), .A3(new_n194), .ZN(new_n238));
  AOI21_X1  g052(.A(KEYINPUT65), .B1(new_n238), .B2(G131), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n238), .A2(KEYINPUT65), .A3(G131), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n221), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(KEYINPUT0), .A2(G128), .ZN(new_n243));
  OR2_X1    g057(.A1(KEYINPUT0), .A2(G128), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n206), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  AND2_X1   g059(.A1(new_n206), .A2(new_n243), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n237), .B1(new_n242), .B2(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n221), .A2(new_n214), .A3(new_n196), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n238), .A2(G131), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT65), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  AOI22_X1  g067(.A1(new_n253), .A2(new_n240), .B1(new_n219), .B2(new_n220), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n250), .B1(new_n254), .B2(new_n247), .ZN(new_n255));
  AOI22_X1  g069(.A1(new_n223), .A2(new_n249), .B1(new_n255), .B2(new_n237), .ZN(new_n256));
  XOR2_X1   g070(.A(KEYINPUT69), .B(KEYINPUT28), .Z(new_n257));
  OAI21_X1  g071(.A(KEYINPUT70), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n253), .A2(new_n240), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n247), .B1(new_n259), .B2(new_n221), .ZN(new_n260));
  AND3_X1   g074(.A1(new_n221), .A2(new_n214), .A3(new_n196), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n237), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(KEYINPUT67), .B1(new_n221), .B2(new_n196), .ZN(new_n263));
  AOI211_X1 g077(.A(new_n204), .B(new_n195), .C1(new_n219), .C2(new_n220), .ZN(new_n264));
  INV_X1    g078(.A(new_n214), .ZN(new_n265));
  NOR3_X1   g079(.A1(new_n263), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  AND2_X1   g080(.A1(new_n234), .A2(new_n236), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n267), .B1(new_n254), .B2(new_n247), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n262), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT70), .ZN(new_n270));
  INV_X1    g084(.A(new_n257), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n223), .A2(new_n249), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT28), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n258), .A2(new_n272), .A3(new_n275), .ZN(new_n276));
  NOR2_X1   g090(.A1(G237), .A2(G953), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(G210), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n278), .B(G101), .ZN(new_n279));
  XNOR2_X1  g093(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n279), .B(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n276), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT30), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n242), .A2(new_n248), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n284), .B1(new_n223), .B2(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n285), .A2(new_n284), .A3(new_n250), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n237), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n281), .B1(new_n266), .B2(new_n268), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT68), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n273), .A2(KEYINPUT68), .A3(new_n281), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n289), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT31), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n289), .A2(new_n292), .A3(KEYINPUT31), .A4(new_n293), .ZN(new_n297));
  AOI22_X1  g111(.A1(new_n189), .A2(new_n283), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n276), .A2(KEYINPUT71), .A3(new_n282), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n188), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n283), .A2(new_n189), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n296), .A2(new_n297), .ZN(new_n302));
  AND4_X1   g116(.A1(new_n188), .A2(new_n301), .A3(new_n299), .A4(new_n302), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n187), .B1(new_n300), .B2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT32), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n301), .A2(new_n302), .A3(new_n299), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(KEYINPUT72), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n298), .A2(new_n188), .A3(new_n299), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n310), .A2(KEYINPUT32), .A3(new_n187), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n289), .A2(new_n273), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(new_n282), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT29), .ZN(new_n314));
  OAI211_X1 g128(.A(new_n313), .B(new_n314), .C1(new_n282), .C2(new_n276), .ZN(new_n315));
  INV_X1    g129(.A(new_n275), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n266), .A2(new_n260), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n273), .B1(new_n317), .B2(new_n267), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n316), .B1(new_n318), .B2(KEYINPUT28), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n282), .A2(new_n314), .ZN(new_n320));
  AOI21_X1  g134(.A(G902), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n315), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G472), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n306), .A2(new_n311), .A3(new_n323), .ZN(new_n324));
  XNOR2_X1  g138(.A(G125), .B(G140), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(KEYINPUT16), .ZN(new_n326));
  INV_X1    g140(.A(G125), .ZN(new_n327));
  OR3_X1    g141(.A1(new_n327), .A2(KEYINPUT16), .A3(G140), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n329), .A2(new_n210), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n330), .B1(new_n210), .B2(new_n325), .ZN(new_n331));
  OAI21_X1  g145(.A(KEYINPUT23), .B1(new_n209), .B2(G119), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT75), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n209), .A2(G119), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  NOR2_X1   g149(.A1(KEYINPUT75), .A2(KEYINPUT23), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n335), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n337), .A2(G110), .ZN(new_n338));
  XOR2_X1   g152(.A(KEYINPUT24), .B(G110), .Z(new_n339));
  XNOR2_X1  g153(.A(new_n339), .B(KEYINPUT73), .ZN(new_n340));
  XNOR2_X1  g154(.A(G119), .B(G128), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n331), .B1(new_n338), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n340), .A2(new_n341), .ZN(new_n344));
  XOR2_X1   g158(.A(new_n344), .B(KEYINPUT74), .Z(new_n345));
  NAND2_X1  g159(.A1(new_n337), .A2(G110), .ZN(new_n346));
  XOR2_X1   g160(.A(new_n346), .B(KEYINPUT76), .Z(new_n347));
  XNOR2_X1  g161(.A(new_n329), .B(new_n210), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n343), .B1(new_n345), .B2(new_n349), .ZN(new_n350));
  XNOR2_X1  g164(.A(KEYINPUT22), .B(G137), .ZN(new_n351));
  INV_X1    g165(.A(G221), .ZN(new_n352));
  INV_X1    g166(.A(G234), .ZN(new_n353));
  NOR3_X1   g167(.A1(new_n352), .A2(new_n353), .A3(G953), .ZN(new_n354));
  XOR2_X1   g168(.A(new_n351), .B(new_n354), .Z(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n350), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(G902), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n343), .B(new_n355), .C1(new_n345), .C2(new_n349), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT25), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n357), .A2(KEYINPUT25), .A3(new_n358), .A4(new_n359), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(G217), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n365), .B1(G234), .B2(new_n358), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n357), .A2(new_n359), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n366), .A2(G902), .ZN(new_n369));
  XOR2_X1   g183(.A(new_n369), .B(KEYINPUT77), .Z(new_n370));
  NOR2_X1   g184(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(KEYINPUT78), .B1(new_n367), .B2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT78), .ZN(new_n374));
  AOI211_X1 g188(.A(new_n374), .B(new_n371), .C1(new_n364), .C2(new_n366), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  AND3_X1   g191(.A1(new_n277), .A2(G143), .A3(G214), .ZN(new_n378));
  AOI21_X1  g192(.A(G143), .B1(new_n277), .B2(G214), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT89), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n382), .A2(KEYINPUT18), .A3(G131), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n325), .B(new_n210), .ZN(new_n384));
  NAND2_X1  g198(.A1(KEYINPUT18), .A2(G131), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n385), .B1(new_n380), .B2(new_n381), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n383), .B(new_n384), .C1(new_n386), .C2(new_n382), .ZN(new_n387));
  OAI211_X1 g201(.A(KEYINPUT17), .B(G131), .C1(new_n378), .C2(new_n379), .ZN(new_n388));
  XNOR2_X1  g202(.A(new_n380), .B(new_n190), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n388), .B1(new_n389), .B2(KEYINPUT17), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n387), .B1(new_n390), .B2(new_n348), .ZN(new_n391));
  XNOR2_X1  g205(.A(G113), .B(G122), .ZN(new_n392));
  INV_X1    g206(.A(G104), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n392), .B(new_n393), .ZN(new_n394));
  XNOR2_X1  g208(.A(new_n325), .B(KEYINPUT19), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n330), .B1(new_n210), .B2(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n394), .B1(new_n396), .B2(new_n389), .ZN(new_n397));
  AOI22_X1  g211(.A1(new_n391), .A2(new_n394), .B1(new_n387), .B2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(G475), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n398), .A2(new_n399), .A3(new_n358), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT90), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n398), .A2(KEYINPUT90), .A3(new_n399), .A4(new_n358), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n402), .A2(KEYINPUT20), .A3(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n394), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(KEYINPUT91), .ZN(new_n406));
  AOI21_X1  g220(.A(G902), .B1(new_n391), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n407), .B1(new_n406), .B2(new_n391), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(G475), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT20), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n400), .A2(new_n401), .A3(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n404), .A2(new_n409), .A3(new_n411), .ZN(new_n412));
  XNOR2_X1  g226(.A(G128), .B(G143), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n413), .B(G134), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n414), .B(KEYINPUT93), .ZN(new_n415));
  INV_X1    g229(.A(G116), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n416), .A2(G122), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n416), .A2(G122), .ZN(new_n419));
  AND2_X1   g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(G107), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n419), .A2(KEYINPUT14), .ZN(new_n423));
  XOR2_X1   g237(.A(new_n423), .B(KEYINPUT94), .Z(new_n424));
  OAI21_X1  g238(.A(new_n418), .B1(new_n419), .B2(KEYINPUT14), .ZN(new_n425));
  OAI21_X1  g239(.A(G107), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n415), .A2(new_n422), .A3(new_n426), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n420), .B(new_n421), .ZN(new_n428));
  XOR2_X1   g242(.A(KEYINPUT92), .B(KEYINPUT13), .Z(new_n429));
  NAND3_X1  g243(.A1(new_n429), .A2(G128), .A3(new_n212), .ZN(new_n430));
  INV_X1    g244(.A(new_n413), .ZN(new_n431));
  OAI211_X1 g245(.A(new_n430), .B(G134), .C1(new_n429), .C2(new_n431), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n428), .B(new_n432), .C1(G134), .C2(new_n431), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n427), .A2(new_n433), .ZN(new_n434));
  XOR2_X1   g248(.A(KEYINPUT9), .B(G234), .Z(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  NOR3_X1   g250(.A1(new_n436), .A2(new_n365), .A3(G953), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n434), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n427), .A2(new_n433), .A3(new_n437), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n439), .A2(KEYINPUT95), .A3(new_n440), .ZN(new_n441));
  OR3_X1    g255(.A1(new_n434), .A2(KEYINPUT95), .A3(new_n438), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n441), .A2(new_n442), .A3(new_n358), .ZN(new_n443));
  INV_X1    g257(.A(G478), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n444), .A2(KEYINPUT15), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n443), .B(new_n445), .ZN(new_n446));
  OR2_X1    g260(.A1(new_n412), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(G953), .ZN(new_n448));
  INV_X1    g262(.A(G952), .ZN(new_n449));
  AND2_X1   g263(.A1(new_n449), .A2(KEYINPUT96), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n449), .A2(KEYINPUT96), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n448), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n452), .B1(G234), .B2(G237), .ZN(new_n453));
  NAND2_X1  g267(.A1(G234), .A2(G237), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n454), .A2(G902), .A3(G953), .ZN(new_n455));
  XOR2_X1   g269(.A(new_n455), .B(KEYINPUT97), .Z(new_n456));
  XNOR2_X1  g270(.A(KEYINPUT21), .B(G898), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n457), .B(KEYINPUT98), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n453), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n447), .A2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(G469), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n393), .A2(G107), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n421), .A2(G104), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT81), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n465), .B(G101), .C1(new_n464), .C2(new_n463), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT79), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n463), .B1(new_n467), .B2(KEYINPUT3), .ZN(new_n468));
  XNOR2_X1  g282(.A(KEYINPUT79), .B(KEYINPUT3), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n468), .B(new_n462), .C1(new_n469), .C2(new_n463), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n466), .B1(new_n470), .B2(G101), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n471), .B(new_n265), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(new_n242), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT12), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n472), .A2(KEYINPUT12), .A3(new_n242), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT82), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n471), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n393), .A2(G107), .ZN(new_n480));
  AND2_X1   g294(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(G101), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n483), .A2(new_n484), .A3(new_n462), .A4(new_n468), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n485), .A2(KEYINPUT82), .A3(new_n466), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n479), .A2(KEYINPUT10), .A3(new_n214), .A4(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n470), .A2(G101), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n488), .A2(KEYINPUT80), .A3(KEYINPUT4), .A4(new_n485), .ZN(new_n489));
  NAND2_X1  g303(.A1(KEYINPUT80), .A2(KEYINPUT4), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n470), .A2(G101), .A3(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n489), .A2(new_n248), .A3(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT10), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n493), .B1(new_n471), .B2(new_n265), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n487), .A2(new_n492), .A3(new_n254), .A4(new_n494), .ZN(new_n495));
  XNOR2_X1  g309(.A(G110), .B(G140), .ZN(new_n496));
  AND2_X1   g310(.A1(new_n448), .A2(G227), .ZN(new_n497));
  XOR2_X1   g311(.A(new_n496), .B(new_n497), .Z(new_n498));
  AND3_X1   g312(.A1(new_n477), .A2(new_n495), .A3(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n487), .A2(new_n494), .A3(new_n492), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(new_n242), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n498), .B1(new_n501), .B2(new_n495), .ZN(new_n502));
  OAI211_X1 g316(.A(new_n461), .B(new_n358), .C1(new_n499), .C2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n477), .A2(new_n495), .ZN(new_n504));
  INV_X1    g318(.A(new_n498), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n501), .A2(new_n495), .A3(new_n498), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n506), .A2(G469), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(G469), .A2(G902), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n503), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT83), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n352), .B1(new_n435), .B2(new_n358), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  AND3_X1   g327(.A1(new_n510), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n511), .B1(new_n510), .B2(new_n513), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n489), .A2(new_n237), .A3(new_n491), .ZN(new_n517));
  NOR3_X1   g331(.A1(new_n416), .A2(KEYINPUT5), .A3(G119), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n518), .B1(new_n230), .B2(KEYINPUT5), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n232), .B1(G113), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n479), .A2(new_n486), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n517), .A2(new_n521), .ZN(new_n522));
  XOR2_X1   g336(.A(G110), .B(G122), .Z(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n524), .A2(KEYINPUT86), .ZN(new_n525));
  AOI21_X1  g339(.A(KEYINPUT6), .B1(new_n522), .B2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n522), .A2(new_n523), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n522), .A2(KEYINPUT6), .A3(new_n525), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n527), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n248), .A2(G125), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n214), .A2(new_n327), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(G224), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n535), .A2(G953), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  XNOR2_X1  g351(.A(new_n534), .B(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n531), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n537), .A2(KEYINPUT87), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n532), .A2(new_n533), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n537), .A2(KEYINPUT7), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n541), .B(new_n542), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n523), .B(KEYINPUT8), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n520), .B(new_n471), .ZN(new_n545));
  OAI211_X1 g359(.A(new_n529), .B(new_n543), .C1(new_n544), .C2(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n539), .A2(new_n358), .A3(new_n546), .ZN(new_n547));
  OAI21_X1  g361(.A(G210), .B1(G237), .B2(G902), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n539), .A2(new_n358), .A3(new_n548), .A4(new_n546), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n550), .A2(new_n551), .A3(KEYINPUT88), .ZN(new_n552));
  OR2_X1    g366(.A1(new_n551), .A2(KEYINPUT88), .ZN(new_n553));
  OAI21_X1  g367(.A(G214), .B1(G237), .B2(G902), .ZN(new_n554));
  XOR2_X1   g368(.A(new_n554), .B(KEYINPUT84), .Z(new_n555));
  XOR2_X1   g369(.A(new_n555), .B(KEYINPUT85), .Z(new_n556));
  NAND3_X1  g370(.A1(new_n552), .A2(new_n553), .A3(new_n556), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n516), .A2(new_n557), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n324), .A2(new_n377), .A3(new_n460), .A4(new_n558), .ZN(new_n559));
  XNOR2_X1  g373(.A(KEYINPUT99), .B(G101), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n559), .B(new_n560), .ZN(G3));
  NOR2_X1   g375(.A1(new_n376), .A2(new_n516), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT100), .ZN(new_n563));
  AOI21_X1  g377(.A(G902), .B1(new_n308), .B2(new_n309), .ZN(new_n564));
  INV_X1    g378(.A(G472), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n563), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n358), .B1(new_n300), .B2(new_n303), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n567), .A2(KEYINPUT100), .A3(G472), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n562), .A2(new_n566), .A3(new_n568), .A4(new_n304), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n555), .B1(new_n550), .B2(new_n551), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  NOR3_X1   g385(.A1(new_n569), .A2(new_n459), .A3(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n412), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT33), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n441), .A2(new_n442), .A3(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n439), .A2(KEYINPUT33), .A3(new_n440), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n575), .A2(G478), .A3(new_n358), .A4(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n443), .A2(new_n444), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n573), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n572), .A2(new_n581), .ZN(new_n582));
  XOR2_X1   g396(.A(KEYINPUT34), .B(G104), .Z(new_n583));
  XNOR2_X1  g397(.A(new_n582), .B(new_n583), .ZN(G6));
  NAND2_X1  g398(.A1(new_n573), .A2(new_n446), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n572), .A2(new_n586), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n587), .B(new_n421), .ZN(new_n588));
  XNOR2_X1  g402(.A(KEYINPUT101), .B(KEYINPUT35), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n588), .B(new_n589), .ZN(G9));
  NAND4_X1  g404(.A1(new_n558), .A2(new_n566), .A3(new_n568), .A4(new_n304), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n356), .A2(KEYINPUT36), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n350), .B(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n370), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n367), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n460), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n591), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(KEYINPUT37), .B(G110), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n598), .B(new_n599), .ZN(G12));
  AOI21_X1  g414(.A(KEYINPUT32), .B1(new_n310), .B2(new_n187), .ZN(new_n601));
  INV_X1    g415(.A(new_n187), .ZN(new_n602));
  AOI211_X1 g416(.A(new_n305), .B(new_n602), .C1(new_n308), .C2(new_n309), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n516), .B1(new_n604), .B2(new_n323), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT103), .ZN(new_n606));
  XNOR2_X1  g420(.A(KEYINPUT102), .B(G900), .ZN(new_n607));
  AND2_X1   g421(.A1(new_n456), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n608), .A2(new_n453), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n586), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n611), .A2(new_n571), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n605), .A2(new_n606), .A3(new_n596), .A4(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n516), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n324), .A2(new_n614), .A3(new_n596), .A4(new_n612), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(KEYINPUT103), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(G128), .ZN(G30));
  NAND2_X1  g432(.A1(new_n318), .A2(new_n282), .ZN(new_n619));
  XOR2_X1   g433(.A(new_n619), .B(KEYINPUT105), .Z(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n294), .ZN(new_n621));
  AND2_X1   g435(.A1(new_n621), .A2(KEYINPUT106), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n358), .B1(new_n621), .B2(KEYINPUT106), .ZN(new_n623));
  OAI21_X1  g437(.A(G472), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n604), .A2(new_n624), .ZN(new_n625));
  XOR2_X1   g439(.A(new_n609), .B(KEYINPUT39), .Z(new_n626));
  NAND2_X1  g440(.A1(new_n614), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(KEYINPUT40), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n552), .A2(new_n553), .ZN(new_n629));
  XNOR2_X1  g443(.A(KEYINPUT104), .B(KEYINPUT38), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n412), .A2(new_n446), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n632), .A2(new_n555), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n625), .A2(new_n628), .A3(new_n631), .A4(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n596), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n635), .B1(new_n627), .B2(KEYINPUT40), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(new_n212), .ZN(G45));
  NOR3_X1   g452(.A1(new_n573), .A2(new_n580), .A3(new_n609), .ZN(new_n639));
  AND3_X1   g453(.A1(new_n639), .A2(KEYINPUT107), .A3(new_n570), .ZN(new_n640));
  AOI21_X1  g454(.A(KEYINPUT107), .B1(new_n639), .B2(new_n570), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n642), .A2(new_n324), .A3(new_n614), .A4(new_n596), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(G146), .ZN(G48));
  OR2_X1    g458(.A1(new_n499), .A2(new_n502), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n358), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(G469), .ZN(new_n647));
  AND2_X1   g461(.A1(new_n647), .A2(new_n503), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n513), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n649), .A2(new_n571), .ZN(new_n650));
  AND4_X1   g464(.A1(new_n324), .A2(new_n377), .A3(new_n581), .A4(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n459), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(KEYINPUT41), .B(G113), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G15));
  AOI21_X1  g469(.A(new_n376), .B1(new_n604), .B2(new_n323), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n585), .A2(new_n459), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n656), .A2(KEYINPUT108), .A3(new_n650), .A4(new_n657), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n324), .A2(new_n377), .A3(new_n650), .A4(new_n657), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT108), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G116), .ZN(G18));
  INV_X1    g477(.A(new_n597), .ZN(new_n664));
  AND3_X1   g478(.A1(new_n324), .A2(new_n664), .A3(new_n650), .ZN(new_n665));
  XOR2_X1   g479(.A(new_n665), .B(G119), .Z(G21));
  OR2_X1    g480(.A1(new_n319), .A2(new_n281), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n602), .B1(new_n667), .B2(new_n302), .ZN(new_n668));
  OAI21_X1  g482(.A(KEYINPUT109), .B1(new_n564), .B2(new_n565), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT109), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n567), .A2(new_n670), .A3(G472), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n668), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n367), .A2(new_n372), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(KEYINPUT110), .ZN(new_n674));
  AND2_X1   g488(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n632), .A2(new_n459), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n675), .A2(new_n650), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G122), .ZN(G24));
  NAND4_X1  g492(.A1(new_n672), .A2(new_n596), .A3(new_n639), .A4(new_n650), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G125), .ZN(G27));
  AOI21_X1  g494(.A(new_n555), .B1(new_n552), .B2(new_n553), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n510), .A2(new_n513), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  AND4_X1   g497(.A1(KEYINPUT42), .A2(new_n681), .A3(new_n639), .A4(new_n683), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n324), .A2(new_n674), .A3(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT111), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n324), .A2(new_n684), .A3(KEYINPUT111), .A4(new_n674), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT42), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n681), .A2(new_n683), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n324), .A2(new_n377), .A3(new_n639), .A4(new_n691), .ZN(new_n692));
  AOI22_X1  g506(.A1(new_n687), .A2(new_n688), .B1(new_n689), .B2(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(new_n190), .ZN(G33));
  NAND2_X1  g508(.A1(new_n324), .A2(new_n377), .ZN(new_n695));
  NOR3_X1   g509(.A1(new_n695), .A2(new_n611), .A3(new_n690), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(new_n193), .ZN(G36));
  NAND2_X1  g511(.A1(new_n506), .A2(new_n507), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT45), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n506), .A2(KEYINPUT45), .A3(new_n507), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n700), .A2(G469), .A3(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n702), .A2(KEYINPUT46), .A3(new_n509), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(new_n503), .ZN(new_n704));
  AOI21_X1  g518(.A(KEYINPUT46), .B1(new_n702), .B2(new_n509), .ZN(new_n705));
  OR2_X1    g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n706), .A2(new_n513), .A3(new_n626), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(KEYINPUT112), .ZN(new_n708));
  INV_X1    g522(.A(new_n681), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n566), .A2(new_n568), .A3(new_n304), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n573), .A2(new_n579), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT43), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n710), .A2(new_n596), .A3(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT44), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n709), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  OAI211_X1 g530(.A(new_n708), .B(new_n716), .C1(new_n715), .C2(new_n714), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G137), .ZN(G39));
  NAND2_X1  g532(.A1(new_n706), .A2(new_n513), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(KEYINPUT47), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT47), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n706), .A2(new_n721), .A3(new_n513), .ZN(new_n722));
  AND3_X1   g536(.A1(new_n720), .A2(new_n639), .A3(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(new_n324), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n377), .A2(new_n709), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n723), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT113), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n723), .A2(KEYINPUT113), .A3(new_n724), .A4(new_n725), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G140), .ZN(G42));
  INV_X1    g545(.A(KEYINPUT50), .ZN(new_n732));
  INV_X1    g546(.A(new_n649), .ZN(new_n733));
  AND2_X1   g547(.A1(new_n713), .A2(new_n453), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n675), .A2(new_n555), .A3(new_n733), .A4(new_n734), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n732), .B1(new_n735), .B2(new_n631), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  NOR3_X1   g551(.A1(new_n735), .A2(new_n732), .A3(new_n631), .ZN(new_n738));
  OAI21_X1  g552(.A(KEYINPUT116), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(new_n738), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT116), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n740), .A2(new_n741), .A3(new_n736), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n604), .A2(new_n624), .A3(new_n733), .A4(new_n681), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n377), .A2(new_n453), .ZN(new_n744));
  NOR3_X1   g558(.A1(new_n743), .A2(new_n579), .A3(new_n744), .ZN(new_n745));
  AND3_X1   g559(.A1(new_n734), .A2(new_n733), .A3(new_n681), .ZN(new_n746));
  AND2_X1   g560(.A1(new_n672), .A2(new_n596), .ZN(new_n747));
  AOI22_X1  g561(.A1(new_n745), .A2(new_n573), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  AND3_X1   g562(.A1(new_n675), .A2(new_n681), .A3(new_n734), .ZN(new_n749));
  INV_X1    g563(.A(new_n720), .ZN(new_n750));
  INV_X1    g564(.A(new_n722), .ZN(new_n751));
  INV_X1    g565(.A(new_n648), .ZN(new_n752));
  OAI22_X1  g566(.A1(new_n750), .A2(new_n751), .B1(new_n513), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n749), .A2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT115), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n749), .A2(new_n753), .A3(KEYINPUT115), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n739), .A2(new_n742), .A3(new_n748), .A4(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT51), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n760), .B1(new_n749), .B2(new_n753), .ZN(new_n762));
  OAI211_X1 g576(.A(new_n748), .B(new_n762), .C1(new_n737), .C2(new_n738), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n743), .A2(new_n744), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n452), .B1(new_n764), .B2(new_n581), .ZN(new_n765));
  AND2_X1   g579(.A1(new_n324), .A2(new_n674), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n746), .A2(new_n766), .ZN(new_n767));
  XOR2_X1   g581(.A(KEYINPUT117), .B(KEYINPUT48), .Z(new_n768));
  XNOR2_X1  g582(.A(new_n767), .B(new_n768), .ZN(new_n769));
  AND3_X1   g583(.A1(new_n763), .A2(new_n765), .A3(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n675), .A2(new_n650), .A3(new_n734), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n761), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT118), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n679), .A2(new_n643), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n571), .A2(new_n632), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n596), .A2(new_n609), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n625), .A2(new_n683), .A3(new_n776), .A4(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n617), .A2(new_n775), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(KEYINPUT52), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT52), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n617), .A2(new_n775), .A3(new_n781), .A4(new_n778), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n665), .B1(new_n651), .B2(new_n652), .ZN(new_n784));
  AND3_X1   g598(.A1(new_n662), .A2(new_n677), .A3(new_n784), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n691), .A2(new_n639), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(new_n672), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n447), .A2(new_n609), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n324), .A2(new_n788), .A3(new_n614), .A4(new_n681), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n635), .B1(new_n787), .B2(new_n789), .ZN(new_n790));
  NOR3_X1   g604(.A1(new_n693), .A2(new_n696), .A3(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(new_n710), .ZN(new_n792));
  NOR3_X1   g606(.A1(new_n557), .A2(new_n573), .A3(new_n580), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n792), .A2(new_n652), .A3(new_n562), .A4(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(new_n559), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n657), .A2(new_n553), .A3(new_n552), .A4(new_n556), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n569), .A2(new_n796), .ZN(new_n797));
  OAI21_X1  g611(.A(KEYINPUT114), .B1(new_n598), .B2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT114), .ZN(new_n799));
  OAI221_X1 g613(.A(new_n799), .B1(new_n591), .B2(new_n597), .C1(new_n569), .C2(new_n796), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n795), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n785), .A2(new_n791), .A3(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n783), .A2(new_n802), .A3(KEYINPUT53), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT53), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n780), .A2(new_n782), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n785), .A2(new_n791), .A3(new_n801), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n804), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n803), .A2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT54), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n803), .A2(KEYINPUT54), .A3(new_n807), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n761), .A2(KEYINPUT118), .A3(new_n770), .A4(new_n771), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n774), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n814), .B1(G952), .B2(G953), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n674), .B1(new_n752), .B2(KEYINPUT49), .ZN(new_n816));
  AOI211_X1 g630(.A(new_n512), .B(new_n816), .C1(KEYINPUT49), .C2(new_n752), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n625), .A2(new_n631), .A3(new_n711), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n817), .A2(new_n556), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n815), .A2(new_n819), .ZN(G75));
  INV_X1    g634(.A(KEYINPUT120), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n821), .B1(new_n808), .B2(G902), .ZN(new_n822));
  AOI211_X1 g636(.A(KEYINPUT120), .B(new_n358), .C1(new_n803), .C2(new_n807), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n549), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n531), .B(KEYINPUT119), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n825), .B(KEYINPUT55), .ZN(new_n826));
  INV_X1    g640(.A(new_n538), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n826), .B(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(new_n828), .ZN(new_n829));
  XOR2_X1   g643(.A(KEYINPUT121), .B(KEYINPUT56), .Z(new_n830));
  NAND3_X1  g644(.A1(new_n824), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n448), .A2(G952), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n808), .A2(G210), .A3(G902), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n828), .B1(new_n834), .B2(KEYINPUT56), .ZN(new_n835));
  AND3_X1   g649(.A1(new_n831), .A2(new_n833), .A3(new_n835), .ZN(G51));
  AOI21_X1  g650(.A(KEYINPUT53), .B1(new_n783), .B2(new_n802), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n805), .A2(new_n806), .A3(new_n804), .ZN(new_n838));
  OAI21_X1  g652(.A(G902), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(KEYINPUT120), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n808), .A2(new_n821), .A3(G902), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(new_n702), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n509), .A2(KEYINPUT57), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n810), .A2(new_n811), .A3(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n509), .A2(KEYINPUT57), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n645), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n832), .B1(new_n844), .B2(new_n848), .ZN(G54));
  OAI211_X1 g663(.A(KEYINPUT58), .B(G475), .C1(new_n822), .C2(new_n823), .ZN(new_n850));
  INV_X1    g664(.A(new_n398), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n842), .A2(KEYINPUT58), .A3(G475), .A4(new_n398), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n852), .A2(new_n853), .A3(new_n833), .ZN(G60));
  NAND2_X1  g668(.A1(G478), .A2(G902), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n855), .B(KEYINPUT59), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n810), .A2(new_n811), .A3(new_n856), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n575), .A2(new_n576), .ZN(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n857), .A2(new_n859), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n860), .A2(new_n861), .A3(new_n832), .ZN(G63));
  XOR2_X1   g676(.A(KEYINPUT122), .B(KEYINPUT61), .Z(new_n863));
  NAND2_X1  g677(.A1(G217), .A2(G902), .ZN(new_n864));
  XOR2_X1   g678(.A(new_n864), .B(KEYINPUT60), .Z(new_n865));
  NAND3_X1  g679(.A1(new_n808), .A2(new_n593), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(new_n833), .ZN(new_n867));
  AOI22_X1  g681(.A1(new_n808), .A2(new_n865), .B1(new_n359), .B2(new_n357), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n863), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(KEYINPUT123), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n867), .A2(new_n868), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(KEYINPUT61), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT123), .ZN(new_n873));
  OAI211_X1 g687(.A(new_n873), .B(new_n863), .C1(new_n867), .C2(new_n868), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n870), .A2(new_n872), .A3(new_n874), .ZN(G66));
  AND2_X1   g689(.A1(new_n785), .A2(new_n801), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n876), .A2(G953), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n458), .A2(new_n535), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n878), .A2(new_n448), .ZN(new_n879));
  OAI21_X1  g693(.A(KEYINPUT124), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n880), .B1(KEYINPUT124), .B2(new_n879), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n825), .B1(G898), .B2(new_n448), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n881), .B(new_n882), .ZN(G69));
  NAND2_X1  g697(.A1(G227), .A2(G900), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n617), .A2(new_n775), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n708), .A2(new_n766), .A3(new_n776), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(KEYINPUT126), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n730), .A2(new_n717), .A3(new_n885), .A4(new_n887), .ZN(new_n888));
  OR2_X1    g702(.A1(new_n886), .A2(KEYINPUT126), .ZN(new_n889));
  INV_X1    g703(.A(new_n693), .ZN(new_n890));
  INV_X1    g704(.A(new_n696), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n448), .B1(new_n888), .B2(new_n892), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n448), .A2(G900), .ZN(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(new_n895));
  AND3_X1   g709(.A1(new_n893), .A2(KEYINPUT127), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g710(.A(KEYINPUT127), .B1(new_n893), .B2(new_n895), .ZN(new_n897));
  OR2_X1    g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n286), .A2(new_n288), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n899), .B(KEYINPUT125), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n900), .B(new_n395), .Z(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  OAI211_X1 g716(.A(G953), .B(new_n884), .C1(new_n898), .C2(new_n902), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n885), .B1(new_n636), .B2(new_n634), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n904), .B(KEYINPUT62), .Z(new_n905));
  AND2_X1   g719(.A1(new_n730), .A2(new_n717), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n656), .B1(new_n581), .B2(new_n586), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n907), .A2(new_n627), .A3(new_n709), .ZN(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  AND3_X1   g723(.A1(new_n905), .A2(new_n906), .A3(new_n909), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n902), .B1(new_n910), .B2(G953), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n901), .B1(new_n896), .B2(new_n897), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n884), .A2(G953), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n903), .A2(new_n914), .ZN(G72));
  NAND4_X1  g729(.A1(new_n905), .A2(new_n876), .A3(new_n906), .A4(new_n909), .ZN(new_n916));
  NAND2_X1  g730(.A1(G472), .A2(G902), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n917), .B(KEYINPUT63), .Z(new_n918));
  NAND2_X1  g732(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n919), .A2(new_n281), .A3(new_n312), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n313), .A2(new_n294), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n808), .A2(new_n918), .A3(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n888), .A2(new_n892), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n923), .A2(new_n801), .A3(new_n785), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n924), .A2(new_n918), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n312), .A2(new_n281), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n832), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  AND3_X1   g741(.A1(new_n920), .A2(new_n922), .A3(new_n927), .ZN(G57));
endmodule


