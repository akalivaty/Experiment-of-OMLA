

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737;

  XNOR2_X1 U374 ( .A(n533), .B(n532), .ZN(n582) );
  INV_X2 U375 ( .A(G953), .ZN(n712) );
  NOR2_X2 U376 ( .A1(G953), .A2(G237), .ZN(n500) );
  AND2_X4 U377 ( .A1(n425), .A2(n607), .ZN(n696) );
  AND2_X2 U378 ( .A1(n582), .A2(n575), .ZN(n586) );
  XNOR2_X2 U379 ( .A(n580), .B(KEYINPUT35), .ZN(n733) );
  XOR2_X1 U380 ( .A(n521), .B(KEYINPUT99), .Z(n663) );
  NAND2_X2 U381 ( .A1(n519), .A2(n526), .ZN(n630) );
  INV_X1 U382 ( .A(G113), .ZN(n369) );
  XNOR2_X1 U383 ( .A(n688), .B(n372), .ZN(n691) );
  NAND2_X1 U384 ( .A1(n556), .A2(n381), .ZN(n721) );
  NOR2_X1 U385 ( .A1(n584), .A2(n734), .ZN(n368) );
  XOR2_X1 U386 ( .A(KEYINPUT103), .B(n583), .Z(n731) );
  NOR2_X1 U387 ( .A1(n736), .A2(n735), .ZN(n411) );
  AND2_X1 U388 ( .A1(n589), .A2(n577), .ZN(n370) );
  XNOR2_X1 U389 ( .A(n389), .B(n450), .ZN(n533) );
  OR2_X1 U390 ( .A1(n690), .A2(G902), .ZN(n389) );
  INV_X1 U391 ( .A(n697), .ZN(n698) );
  XNOR2_X1 U392 ( .A(n690), .B(n689), .ZN(n372) );
  XNOR2_X1 U393 ( .A(n720), .B(n449), .ZN(n690) );
  XNOR2_X1 U394 ( .A(n703), .B(n408), .ZN(n476) );
  XNOR2_X1 U395 ( .A(n446), .B(n445), .ZN(n703) );
  XNOR2_X1 U396 ( .A(n459), .B(n458), .ZN(n475) );
  XNOR2_X1 U397 ( .A(n463), .B(n409), .ZN(n408) );
  INV_X1 U398 ( .A(n444), .ZN(n446) );
  XNOR2_X1 U399 ( .A(n369), .B(G116), .ZN(n459) );
  XNOR2_X1 U400 ( .A(KEYINPUT3), .B(G119), .ZN(n458) );
  XNOR2_X1 U401 ( .A(KEYINPUT76), .B(G110), .ZN(n445) );
  XNOR2_X1 U402 ( .A(G104), .B(G107), .ZN(n444) );
  INV_X1 U403 ( .A(n643), .ZN(n713) );
  XOR2_X2 U404 ( .A(n587), .B(KEYINPUT88), .Z(n589) );
  XNOR2_X2 U405 ( .A(n379), .B(G143), .ZN(n469) );
  XNOR2_X2 U406 ( .A(G128), .B(KEYINPUT64), .ZN(n379) );
  XNOR2_X1 U407 ( .A(n422), .B(n359), .ZN(n585) );
  OR2_X1 U408 ( .A1(n612), .A2(G902), .ZN(n422) );
  AND2_X1 U409 ( .A1(n391), .A2(n390), .ZN(n679) );
  XOR2_X1 U410 ( .A(KEYINPUT93), .B(KEYINPUT5), .Z(n461) );
  XNOR2_X1 U411 ( .A(n469), .B(G134), .ZN(n487) );
  AND2_X1 U412 ( .A1(n412), .A2(n410), .ZN(n549) );
  NOR2_X1 U413 ( .A1(n548), .A2(n413), .ZN(n412) );
  XNOR2_X1 U414 ( .A(n411), .B(KEYINPUT46), .ZN(n410) );
  XNOR2_X1 U415 ( .A(n388), .B(n487), .ZN(n457) );
  XNOR2_X1 U416 ( .A(n504), .B(n364), .ZN(n388) );
  XNOR2_X1 U417 ( .A(n414), .B(n365), .ZN(n364) );
  INV_X1 U418 ( .A(KEYINPUT4), .ZN(n414) );
  XOR2_X1 U419 ( .A(KEYINPUT68), .B(G140), .Z(n442) );
  XNOR2_X1 U420 ( .A(KEYINPUT23), .B(n719), .ZN(n433) );
  XNOR2_X1 U421 ( .A(n434), .B(n430), .ZN(n384) );
  INV_X1 U422 ( .A(KEYINPUT90), .ZN(n430) );
  XNOR2_X1 U423 ( .A(G119), .B(G110), .ZN(n426) );
  XOR2_X1 U424 ( .A(KEYINPUT9), .B(G107), .Z(n489) );
  XNOR2_X1 U425 ( .A(G116), .B(G122), .ZN(n488) );
  XNOR2_X1 U426 ( .A(KEYINPUT96), .B(KEYINPUT7), .ZN(n490) );
  XOR2_X1 U427 ( .A(KEYINPUT98), .B(KEYINPUT97), .Z(n491) );
  XNOR2_X1 U428 ( .A(G113), .B(G122), .ZN(n498) );
  INV_X1 U429 ( .A(KEYINPUT70), .ZN(n409) );
  XNOR2_X1 U430 ( .A(n457), .B(n443), .ZN(n720) );
  XNOR2_X1 U431 ( .A(n442), .B(KEYINPUT89), .ZN(n443) );
  AND2_X1 U432 ( .A1(n687), .A2(G210), .ZN(n421) );
  OR2_X1 U433 ( .A1(n527), .A2(n484), .ZN(n485) );
  XNOR2_X1 U434 ( .A(n673), .B(KEYINPUT33), .ZN(n577) );
  XNOR2_X1 U435 ( .A(n572), .B(n571), .ZN(n581) );
  XNOR2_X1 U436 ( .A(KEYINPUT22), .B(KEYINPUT72), .ZN(n571) );
  OR2_X1 U437 ( .A1(n385), .A2(n533), .ZN(n516) );
  XNOR2_X1 U438 ( .A(n515), .B(n386), .ZN(n385) );
  XNOR2_X1 U439 ( .A(n387), .B(KEYINPUT28), .ZN(n386) );
  XNOR2_X1 U440 ( .A(n439), .B(n438), .ZN(n597) );
  XNOR2_X1 U441 ( .A(n437), .B(n354), .ZN(n438) );
  XNOR2_X1 U442 ( .A(n451), .B(KEYINPUT92), .ZN(n591) );
  OR2_X1 U443 ( .A1(n651), .A2(n533), .ZN(n451) );
  XNOR2_X1 U444 ( .A(KEYINPUT100), .B(KEYINPUT6), .ZN(n534) );
  NOR2_X1 U445 ( .A1(n581), .A2(n582), .ZN(n596) );
  NAND2_X1 U446 ( .A1(n380), .A2(n713), .ZN(n607) );
  XNOR2_X1 U447 ( .A(n721), .B(n559), .ZN(n380) );
  NOR2_X1 U448 ( .A1(n405), .A2(n681), .ZN(n404) );
  AND2_X1 U449 ( .A1(n712), .A2(n682), .ZN(n399) );
  NAND2_X1 U450 ( .A1(n652), .A2(n651), .ZN(n397) );
  INV_X1 U451 ( .A(KEYINPUT112), .ZN(n396) );
  AND2_X1 U452 ( .A1(n630), .A2(n625), .ZN(n521) );
  XOR2_X1 U453 ( .A(KEYINPUT67), .B(G131), .Z(n504) );
  INV_X1 U454 ( .A(G137), .ZN(n365) );
  XOR2_X1 U455 ( .A(KEYINPUT4), .B(KEYINPUT86), .Z(n472) );
  XNOR2_X1 U456 ( .A(n469), .B(n378), .ZN(n474) );
  XNOR2_X1 U457 ( .A(n470), .B(n468), .ZN(n378) );
  XOR2_X1 U458 ( .A(G137), .B(G128), .Z(n427) );
  XOR2_X1 U459 ( .A(G140), .B(KEYINPUT12), .Z(n502) );
  XOR2_X1 U460 ( .A(G143), .B(G104), .Z(n499) );
  XNOR2_X1 U461 ( .A(n393), .B(n392), .ZN(n391) );
  XNOR2_X1 U462 ( .A(KEYINPUT118), .B(KEYINPUT52), .ZN(n392) );
  NAND2_X1 U463 ( .A1(n353), .A2(n355), .ZN(n393) );
  INV_X1 U464 ( .A(n675), .ZN(n390) );
  INV_X1 U465 ( .A(KEYINPUT106), .ZN(n387) );
  XNOR2_X1 U466 ( .A(n465), .B(n362), .ZN(n423) );
  XNOR2_X1 U467 ( .A(n464), .B(n424), .ZN(n362) );
  XNOR2_X1 U468 ( .A(n475), .B(n407), .ZN(n705) );
  XNOR2_X1 U469 ( .A(KEYINPUT16), .B(G122), .ZN(n407) );
  AND2_X1 U470 ( .A1(n737), .A2(n555), .ZN(n381) );
  XNOR2_X1 U471 ( .A(n549), .B(KEYINPUT48), .ZN(n556) );
  XNOR2_X1 U472 ( .A(n466), .B(n363), .ZN(n467) );
  INV_X1 U473 ( .A(KEYINPUT30), .ZN(n363) );
  XOR2_X1 U474 ( .A(n510), .B(n509), .Z(n520) );
  NOR2_X1 U475 ( .A1(G902), .A2(n608), .ZN(n510) );
  XNOR2_X1 U476 ( .A(n383), .B(n382), .ZN(n697) );
  XNOR2_X1 U477 ( .A(n432), .B(n431), .ZN(n382) );
  XNOR2_X1 U478 ( .A(n433), .B(n384), .ZN(n383) );
  XNOR2_X1 U479 ( .A(n371), .B(n495), .ZN(n693) );
  XNOR2_X1 U480 ( .A(n496), .B(n358), .ZN(n371) );
  XNOR2_X1 U481 ( .A(n447), .B(G146), .ZN(n448) );
  INV_X1 U482 ( .A(n687), .ZN(n416) );
  AND2_X1 U483 ( .A1(n420), .A2(n360), .ZN(n418) );
  NAND2_X1 U484 ( .A1(n696), .A2(n421), .ZN(n420) );
  XNOR2_X1 U485 ( .A(n370), .B(n361), .ZN(n579) );
  XOR2_X1 U486 ( .A(KEYINPUT31), .B(n588), .Z(n635) );
  NOR2_X1 U487 ( .A1(n587), .A2(n657), .ZN(n588) );
  INV_X1 U488 ( .A(n516), .ZN(n518) );
  NAND2_X1 U489 ( .A1(n596), .A2(n357), .ZN(n583) );
  NOR2_X1 U490 ( .A1(n591), .A2(n590), .ZN(n620) );
  AND2_X1 U491 ( .A1(n596), .A2(n376), .ZN(n598) );
  AND2_X1 U492 ( .A1(n595), .A2(n377), .ZN(n376) );
  INV_X1 U493 ( .A(KEYINPUT60), .ZN(n373) );
  XNOR2_X1 U494 ( .A(n367), .B(n366), .ZN(G51) );
  INV_X1 U495 ( .A(KEYINPUT56), .ZN(n366) );
  NAND2_X1 U496 ( .A1(n418), .A2(n415), .ZN(n367) );
  NAND2_X1 U497 ( .A1(n417), .A2(n416), .ZN(n415) );
  NAND2_X1 U498 ( .A1(n403), .A2(n401), .ZN(n683) );
  NAND2_X1 U499 ( .A1(n404), .A2(n402), .ZN(n401) );
  OR2_X1 U500 ( .A1(n676), .A2(n661), .ZN(n353) );
  XOR2_X1 U501 ( .A(KEYINPUT25), .B(KEYINPUT78), .Z(n354) );
  INV_X1 U502 ( .A(n597), .ZN(n377) );
  OR2_X1 U503 ( .A1(n674), .A2(n677), .ZN(n355) );
  AND2_X1 U504 ( .A1(n406), .A2(n647), .ZN(n356) );
  AND2_X1 U505 ( .A1(n655), .A2(n597), .ZN(n357) );
  AND2_X1 U506 ( .A1(G217), .A2(n494), .ZN(n358) );
  XNOR2_X1 U507 ( .A(KEYINPUT94), .B(G472), .ZN(n359) );
  AND2_X1 U508 ( .A1(n419), .A2(n700), .ZN(n360) );
  XNOR2_X1 U509 ( .A(KEYINPUT71), .B(KEYINPUT34), .ZN(n361) );
  XOR2_X1 U510 ( .A(n476), .B(n705), .Z(n477) );
  XNOR2_X1 U511 ( .A(n511), .B(KEYINPUT40), .ZN(n736) );
  NAND2_X1 U512 ( .A1(n643), .A2(n644), .ZN(n606) );
  XNOR2_X2 U513 ( .A(n604), .B(n603), .ZN(n643) );
  XNOR2_X1 U514 ( .A(n368), .B(KEYINPUT44), .ZN(n602) );
  XNOR2_X1 U515 ( .A(n699), .B(n698), .ZN(n701) );
  INV_X1 U516 ( .A(n519), .ZN(n525) );
  XNOR2_X1 U517 ( .A(n497), .B(G478), .ZN(n519) );
  NOR2_X1 U518 ( .A1(n629), .A2(n524), .ZN(n413) );
  XNOR2_X1 U519 ( .A(n374), .B(n373), .ZN(G60) );
  NAND2_X1 U520 ( .A1(n375), .A2(n700), .ZN(n374) );
  XNOR2_X1 U521 ( .A(n610), .B(n609), .ZN(n375) );
  NOR2_X1 U522 ( .A1(n394), .A2(n654), .ZN(n656) );
  XNOR2_X1 U523 ( .A(n397), .B(n395), .ZN(n394) );
  XNOR2_X1 U524 ( .A(n653), .B(n396), .ZN(n395) );
  XNOR2_X2 U525 ( .A(KEYINPUT10), .B(n468), .ZN(n719) );
  XNOR2_X2 U526 ( .A(n398), .B(KEYINPUT0), .ZN(n587) );
  NAND2_X1 U527 ( .A1(n566), .A2(n567), .ZN(n398) );
  XNOR2_X2 U528 ( .A(n538), .B(KEYINPUT19), .ZN(n566) );
  NAND2_X2 U529 ( .A1(n554), .A2(n665), .ZN(n538) );
  NAND2_X1 U530 ( .A1(n400), .A2(n399), .ZN(n403) );
  NAND2_X1 U531 ( .A1(n356), .A2(n648), .ZN(n400) );
  AND2_X1 U532 ( .A1(n648), .A2(n712), .ZN(n402) );
  NAND2_X1 U533 ( .A1(n647), .A2(KEYINPUT120), .ZN(n405) );
  INV_X1 U534 ( .A(n681), .ZN(n406) );
  INV_X1 U535 ( .A(n696), .ZN(n417) );
  OR2_X1 U536 ( .A1(n687), .A2(G210), .ZN(n419) );
  XNOR2_X1 U537 ( .A(n423), .B(n457), .ZN(n612) );
  INV_X1 U538 ( .A(KEYINPUT75), .ZN(n424) );
  INV_X1 U539 ( .A(n487), .ZN(n496) );
  XNOR2_X1 U540 ( .A(n585), .B(n534), .ZN(n595) );
  AND2_X1 U541 ( .A1(n606), .A2(n479), .ZN(n425) );
  INV_X1 U542 ( .A(n639), .ZN(n555) );
  INV_X1 U543 ( .A(KEYINPUT81), .ZN(n640) );
  XNOR2_X1 U544 ( .A(n713), .B(n640), .ZN(n642) );
  XNOR2_X1 U545 ( .A(n476), .B(n448), .ZN(n449) );
  XNOR2_X1 U546 ( .A(n613), .B(KEYINPUT109), .ZN(n614) );
  XNOR2_X1 U547 ( .A(KEYINPUT82), .B(KEYINPUT36), .ZN(n539) );
  XNOR2_X1 U548 ( .A(n615), .B(n614), .ZN(n616) );
  XNOR2_X1 U549 ( .A(n540), .B(n539), .ZN(n541) );
  NAND2_X1 U550 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U551 ( .A1(KEYINPUT2), .A2(KEYINPUT77), .ZN(n559) );
  XNOR2_X1 U552 ( .A(n427), .B(n426), .ZN(n434) );
  XOR2_X1 U553 ( .A(n442), .B(KEYINPUT24), .Z(n432) );
  XOR2_X1 U554 ( .A(KEYINPUT8), .B(KEYINPUT66), .Z(n429) );
  NAND2_X1 U555 ( .A1(G234), .A2(n712), .ZN(n428) );
  XNOR2_X1 U556 ( .A(n429), .B(n428), .ZN(n494) );
  NAND2_X1 U557 ( .A1(n494), .A2(G221), .ZN(n431) );
  XNOR2_X2 U558 ( .A(G125), .B(G146), .ZN(n468) );
  NOR2_X1 U559 ( .A1(G902), .A2(n697), .ZN(n439) );
  XOR2_X1 U560 ( .A(KEYINPUT91), .B(KEYINPUT20), .Z(n436) );
  XNOR2_X1 U561 ( .A(G902), .B(KEYINPUT15), .ZN(n605) );
  NAND2_X1 U562 ( .A1(G234), .A2(n605), .ZN(n435) );
  XNOR2_X1 U563 ( .A(n436), .B(n435), .ZN(n440) );
  NAND2_X1 U564 ( .A1(G217), .A2(n440), .ZN(n437) );
  NAND2_X1 U565 ( .A1(G221), .A2(n440), .ZN(n441) );
  XOR2_X1 U566 ( .A(n441), .B(KEYINPUT21), .Z(n649) );
  NAND2_X1 U567 ( .A1(n377), .A2(n649), .ZN(n651) );
  XOR2_X2 U568 ( .A(KEYINPUT65), .B(G101), .Z(n463) );
  AND2_X1 U569 ( .A1(G227), .A2(n712), .ZN(n447) );
  XNOR2_X1 U570 ( .A(KEYINPUT69), .B(G469), .ZN(n450) );
  XNOR2_X1 U571 ( .A(n591), .B(KEYINPUT104), .ZN(n528) );
  NAND2_X1 U572 ( .A1(G234), .A2(G237), .ZN(n452) );
  XNOR2_X1 U573 ( .A(n452), .B(KEYINPUT14), .ZN(n454) );
  NAND2_X1 U574 ( .A1(n454), .A2(G952), .ZN(n675) );
  NOR2_X1 U575 ( .A1(n675), .A2(G953), .ZN(n453) );
  XNOR2_X1 U576 ( .A(n453), .B(KEYINPUT87), .ZN(n565) );
  NAND2_X1 U577 ( .A1(G902), .A2(n454), .ZN(n562) );
  NOR2_X1 U578 ( .A1(G900), .A2(n562), .ZN(n455) );
  NAND2_X1 U579 ( .A1(G953), .A2(n455), .ZN(n456) );
  NAND2_X1 U580 ( .A1(n565), .A2(n456), .ZN(n513) );
  NAND2_X1 U581 ( .A1(n500), .A2(G210), .ZN(n460) );
  XNOR2_X1 U582 ( .A(n461), .B(n460), .ZN(n462) );
  XOR2_X1 U583 ( .A(n475), .B(n462), .Z(n465) );
  XNOR2_X1 U584 ( .A(n463), .B(G146), .ZN(n464) );
  OR2_X1 U585 ( .A1(G237), .A2(G902), .ZN(n480) );
  NAND2_X1 U586 ( .A1(G214), .A2(n480), .ZN(n665) );
  NAND2_X1 U587 ( .A1(n585), .A2(n665), .ZN(n466) );
  NAND2_X1 U588 ( .A1(n513), .A2(n467), .ZN(n527) );
  XNOR2_X1 U589 ( .A(KEYINPUT38), .B(KEYINPUT74), .ZN(n483) );
  NAND2_X1 U590 ( .A1(G224), .A2(n712), .ZN(n470) );
  XNOR2_X1 U591 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n471) );
  XNOR2_X1 U592 ( .A(n472), .B(n471), .ZN(n473) );
  XOR2_X1 U593 ( .A(n474), .B(n473), .Z(n478) );
  XNOR2_X1 U594 ( .A(n477), .B(n478), .ZN(n684) );
  INV_X1 U595 ( .A(n605), .ZN(n479) );
  NOR2_X1 U596 ( .A1(n684), .A2(n479), .ZN(n482) );
  NAND2_X1 U597 ( .A1(G210), .A2(n480), .ZN(n481) );
  XNOR2_X2 U598 ( .A(n482), .B(n481), .ZN(n554) );
  XOR2_X1 U599 ( .A(n483), .B(n554), .Z(n666) );
  INV_X1 U600 ( .A(n666), .ZN(n484) );
  NOR2_X1 U601 ( .A1(n528), .A2(n485), .ZN(n486) );
  XNOR2_X1 U602 ( .A(n486), .B(KEYINPUT39), .ZN(n557) );
  XNOR2_X1 U603 ( .A(n489), .B(n488), .ZN(n493) );
  XNOR2_X1 U604 ( .A(n491), .B(n490), .ZN(n492) );
  XOR2_X1 U605 ( .A(n493), .B(n492), .Z(n495) );
  NOR2_X1 U606 ( .A1(G902), .A2(n693), .ZN(n497) );
  XNOR2_X1 U607 ( .A(n499), .B(n498), .ZN(n508) );
  NAND2_X1 U608 ( .A1(G214), .A2(n500), .ZN(n501) );
  XNOR2_X1 U609 ( .A(n502), .B(n501), .ZN(n503) );
  XOR2_X1 U610 ( .A(n503), .B(KEYINPUT11), .Z(n506) );
  XNOR2_X1 U611 ( .A(n504), .B(n719), .ZN(n505) );
  XNOR2_X1 U612 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U613 ( .A(n508), .B(n507), .ZN(n608) );
  XNOR2_X1 U614 ( .A(KEYINPUT13), .B(G475), .ZN(n509) );
  INV_X1 U615 ( .A(n520), .ZN(n526) );
  NOR2_X1 U616 ( .A1(n557), .A2(n630), .ZN(n511) );
  NAND2_X1 U617 ( .A1(n520), .A2(n519), .ZN(n669) );
  NAND2_X1 U618 ( .A1(n666), .A2(n665), .ZN(n662) );
  NOR2_X1 U619 ( .A1(n669), .A2(n662), .ZN(n512) );
  XNOR2_X1 U620 ( .A(n512), .B(KEYINPUT41), .ZN(n676) );
  INV_X1 U621 ( .A(n649), .ZN(n568) );
  NAND2_X1 U622 ( .A1(n513), .A2(n597), .ZN(n514) );
  NOR2_X1 U623 ( .A1(n568), .A2(n514), .ZN(n535) );
  AND2_X1 U624 ( .A1(n585), .A2(n535), .ZN(n515) );
  NOR2_X1 U625 ( .A1(n676), .A2(n516), .ZN(n517) );
  XNOR2_X1 U626 ( .A(n517), .B(KEYINPUT42), .ZN(n735) );
  NAND2_X1 U627 ( .A1(n518), .A2(n566), .ZN(n629) );
  INV_X1 U628 ( .A(n630), .ZN(n632) );
  NAND2_X1 U629 ( .A1(n520), .A2(n525), .ZN(n625) );
  INV_X1 U630 ( .A(n625), .ZN(n634) );
  XOR2_X1 U631 ( .A(KEYINPUT80), .B(n663), .Z(n593) );
  INV_X1 U632 ( .A(n593), .ZN(n522) );
  NOR2_X1 U633 ( .A1(KEYINPUT47), .A2(n522), .ZN(n523) );
  XNOR2_X1 U634 ( .A(n523), .B(KEYINPUT73), .ZN(n524) );
  NAND2_X1 U635 ( .A1(n526), .A2(n525), .ZN(n578) );
  NOR2_X1 U636 ( .A1(n528), .A2(n527), .ZN(n529) );
  NAND2_X1 U637 ( .A1(n554), .A2(n529), .ZN(n530) );
  XOR2_X1 U638 ( .A(KEYINPUT105), .B(n530), .Z(n531) );
  NOR2_X1 U639 ( .A1(n578), .A2(n531), .ZN(n628) );
  INV_X1 U640 ( .A(n628), .ZN(n547) );
  INV_X1 U641 ( .A(KEYINPUT1), .ZN(n532) );
  INV_X1 U642 ( .A(n582), .ZN(n652) );
  XOR2_X1 U643 ( .A(KEYINPUT84), .B(n652), .Z(n561) );
  INV_X1 U644 ( .A(n595), .ZN(n576) );
  NAND2_X1 U645 ( .A1(n535), .A2(n576), .ZN(n536) );
  NOR2_X1 U646 ( .A1(n630), .A2(n536), .ZN(n550) );
  XNOR2_X1 U647 ( .A(KEYINPUT107), .B(n550), .ZN(n537) );
  NOR2_X1 U648 ( .A1(n538), .A2(n537), .ZN(n540) );
  NAND2_X1 U649 ( .A1(n561), .A2(n541), .ZN(n638) );
  NAND2_X1 U650 ( .A1(KEYINPUT47), .A2(n629), .ZN(n542) );
  NAND2_X1 U651 ( .A1(n638), .A2(n542), .ZN(n545) );
  NAND2_X1 U652 ( .A1(KEYINPUT47), .A2(n663), .ZN(n543) );
  XNOR2_X1 U653 ( .A(KEYINPUT79), .B(n543), .ZN(n544) );
  NOR2_X1 U654 ( .A1(n545), .A2(n544), .ZN(n546) );
  NAND2_X1 U655 ( .A1(n547), .A2(n546), .ZN(n548) );
  NAND2_X1 U656 ( .A1(n550), .A2(n665), .ZN(n551) );
  NOR2_X1 U657 ( .A1(n582), .A2(n551), .ZN(n552) );
  XNOR2_X1 U658 ( .A(n552), .B(KEYINPUT43), .ZN(n553) );
  NOR2_X1 U659 ( .A1(n554), .A2(n553), .ZN(n639) );
  NOR2_X1 U660 ( .A1(n557), .A2(n625), .ZN(n558) );
  XOR2_X1 U661 ( .A(KEYINPUT108), .B(n558), .Z(n737) );
  NOR2_X1 U662 ( .A1(n377), .A2(n576), .ZN(n560) );
  NAND2_X1 U663 ( .A1(n561), .A2(n560), .ZN(n573) );
  INV_X1 U664 ( .A(n669), .ZN(n570) );
  INV_X1 U665 ( .A(n562), .ZN(n563) );
  NOR2_X1 U666 ( .A1(G898), .A2(n712), .ZN(n707) );
  NAND2_X1 U667 ( .A1(n563), .A2(n707), .ZN(n564) );
  NAND2_X1 U668 ( .A1(n565), .A2(n564), .ZN(n567) );
  NOR2_X1 U669 ( .A1(n568), .A2(n587), .ZN(n569) );
  NAND2_X1 U670 ( .A1(n570), .A2(n569), .ZN(n572) );
  NOR2_X1 U671 ( .A1(n573), .A2(n581), .ZN(n574) );
  XNOR2_X1 U672 ( .A(n574), .B(KEYINPUT32), .ZN(n734) );
  INV_X1 U673 ( .A(n651), .ZN(n575) );
  NAND2_X1 U674 ( .A1(n586), .A2(n576), .ZN(n673) );
  NOR2_X2 U675 ( .A1(n579), .A2(n578), .ZN(n580) );
  INV_X1 U676 ( .A(n585), .ZN(n655) );
  NAND2_X1 U677 ( .A1(n733), .A2(n731), .ZN(n584) );
  NAND2_X1 U678 ( .A1(n586), .A2(n585), .ZN(n657) );
  NAND2_X1 U679 ( .A1(n655), .A2(n589), .ZN(n590) );
  NOR2_X1 U680 ( .A1(n635), .A2(n620), .ZN(n592) );
  XNOR2_X1 U681 ( .A(n592), .B(KEYINPUT95), .ZN(n594) );
  NAND2_X1 U682 ( .A1(n594), .A2(n593), .ZN(n599) );
  XNOR2_X1 U683 ( .A(n598), .B(KEYINPUT101), .ZN(n730) );
  NAND2_X1 U684 ( .A1(n599), .A2(n730), .ZN(n600) );
  XOR2_X1 U685 ( .A(KEYINPUT102), .B(n600), .Z(n601) );
  NAND2_X1 U686 ( .A1(n602), .A2(n601), .ZN(n604) );
  INV_X1 U687 ( .A(KEYINPUT45), .ZN(n603) );
  INV_X1 U688 ( .A(KEYINPUT2), .ZN(n644) );
  NAND2_X1 U689 ( .A1(G475), .A2(n696), .ZN(n610) );
  XNOR2_X1 U690 ( .A(n608), .B(KEYINPUT59), .ZN(n609) );
  NOR2_X1 U691 ( .A1(n712), .A2(G952), .ZN(n611) );
  XOR2_X1 U692 ( .A(n611), .B(KEYINPUT85), .Z(n695) );
  INV_X1 U693 ( .A(n695), .ZN(n700) );
  NAND2_X1 U694 ( .A1(G472), .A2(n696), .ZN(n615) );
  XNOR2_X1 U695 ( .A(n612), .B(KEYINPUT62), .ZN(n613) );
  NAND2_X1 U696 ( .A1(n616), .A2(n700), .ZN(n617) );
  XNOR2_X1 U697 ( .A(n617), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U698 ( .A1(n620), .A2(n632), .ZN(n618) );
  XNOR2_X1 U699 ( .A(n618), .B(KEYINPUT110), .ZN(n619) );
  XNOR2_X1 U700 ( .A(G104), .B(n619), .ZN(G6) );
  XOR2_X1 U701 ( .A(KEYINPUT26), .B(KEYINPUT27), .Z(n622) );
  NAND2_X1 U702 ( .A1(n620), .A2(n634), .ZN(n621) );
  XNOR2_X1 U703 ( .A(n622), .B(n621), .ZN(n624) );
  XOR2_X1 U704 ( .A(G107), .B(KEYINPUT111), .Z(n623) );
  XNOR2_X1 U705 ( .A(n624), .B(n623), .ZN(G9) );
  NOR2_X1 U706 ( .A1(n625), .A2(n629), .ZN(n627) );
  XNOR2_X1 U707 ( .A(G128), .B(KEYINPUT29), .ZN(n626) );
  XNOR2_X1 U708 ( .A(n627), .B(n626), .ZN(G30) );
  XOR2_X1 U709 ( .A(G143), .B(n628), .Z(G45) );
  NOR2_X1 U710 ( .A1(n630), .A2(n629), .ZN(n631) );
  XOR2_X1 U711 ( .A(G146), .B(n631), .Z(G48) );
  NAND2_X1 U712 ( .A1(n635), .A2(n632), .ZN(n633) );
  XNOR2_X1 U713 ( .A(n633), .B(G113), .ZN(G15) );
  NAND2_X1 U714 ( .A1(n635), .A2(n634), .ZN(n636) );
  XNOR2_X1 U715 ( .A(n636), .B(G116), .ZN(G18) );
  XOR2_X1 U716 ( .A(G125), .B(KEYINPUT37), .Z(n637) );
  XNOR2_X1 U717 ( .A(n638), .B(n637), .ZN(G27) );
  XOR2_X1 U718 ( .A(G140), .B(n639), .Z(G42) );
  NOR2_X1 U719 ( .A1(KEYINPUT2), .A2(n721), .ZN(n641) );
  NAND2_X1 U720 ( .A1(n642), .A2(n641), .ZN(n648) );
  NOR2_X1 U721 ( .A1(n721), .A2(n643), .ZN(n645) );
  NOR2_X1 U722 ( .A1(n645), .A2(n644), .ZN(n646) );
  NAND2_X1 U723 ( .A1(n640), .A2(n646), .ZN(n647) );
  NOR2_X1 U724 ( .A1(n377), .A2(n649), .ZN(n650) );
  XOR2_X1 U725 ( .A(KEYINPUT49), .B(n650), .Z(n654) );
  XOR2_X1 U726 ( .A(KEYINPUT50), .B(KEYINPUT113), .Z(n653) );
  NAND2_X1 U727 ( .A1(n656), .A2(n655), .ZN(n658) );
  NAND2_X1 U728 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U729 ( .A(n659), .B(KEYINPUT114), .ZN(n660) );
  XNOR2_X1 U730 ( .A(n660), .B(KEYINPUT51), .ZN(n661) );
  NOR2_X1 U731 ( .A1(n663), .A2(n662), .ZN(n664) );
  XOR2_X1 U732 ( .A(KEYINPUT117), .B(n664), .Z(n672) );
  NOR2_X1 U733 ( .A1(n666), .A2(n665), .ZN(n667) );
  XOR2_X1 U734 ( .A(KEYINPUT115), .B(n667), .Z(n668) );
  NOR2_X1 U735 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U736 ( .A(KEYINPUT116), .B(n670), .ZN(n671) );
  NOR2_X1 U737 ( .A1(n672), .A2(n671), .ZN(n674) );
  XOR2_X1 U738 ( .A(KEYINPUT33), .B(n673), .Z(n677) );
  NOR2_X1 U739 ( .A1(n677), .A2(n676), .ZN(n678) );
  NOR2_X1 U740 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U741 ( .A(n680), .B(KEYINPUT119), .ZN(n681) );
  INV_X1 U742 ( .A(KEYINPUT120), .ZN(n682) );
  XNOR2_X1 U743 ( .A(KEYINPUT53), .B(n683), .ZN(G75) );
  XOR2_X1 U744 ( .A(KEYINPUT83), .B(KEYINPUT55), .Z(n686) );
  XNOR2_X1 U745 ( .A(n684), .B(KEYINPUT54), .ZN(n685) );
  XNOR2_X1 U746 ( .A(n686), .B(n685), .ZN(n687) );
  XOR2_X1 U747 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n689) );
  NAND2_X1 U748 ( .A1(n696), .A2(G469), .ZN(n688) );
  NOR2_X1 U749 ( .A1(n695), .A2(n691), .ZN(G54) );
  NAND2_X1 U750 ( .A1(G478), .A2(n696), .ZN(n692) );
  XNOR2_X1 U751 ( .A(n693), .B(n692), .ZN(n694) );
  NOR2_X1 U752 ( .A1(n695), .A2(n694), .ZN(G63) );
  NAND2_X1 U753 ( .A1(G217), .A2(n696), .ZN(n699) );
  XNOR2_X1 U754 ( .A(n702), .B(KEYINPUT121), .ZN(G66) );
  XOR2_X1 U755 ( .A(n703), .B(G101), .Z(n704) );
  XOR2_X1 U756 ( .A(n705), .B(n704), .Z(n706) );
  NOR2_X1 U757 ( .A1(n707), .A2(n706), .ZN(n717) );
  XOR2_X1 U758 ( .A(KEYINPUT61), .B(KEYINPUT123), .Z(n709) );
  NAND2_X1 U759 ( .A1(G224), .A2(G953), .ZN(n708) );
  XNOR2_X1 U760 ( .A(n709), .B(n708), .ZN(n710) );
  XNOR2_X1 U761 ( .A(KEYINPUT122), .B(n710), .ZN(n711) );
  NAND2_X1 U762 ( .A1(n711), .A2(G898), .ZN(n715) );
  NAND2_X1 U763 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U764 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U765 ( .A(n717), .B(n716), .ZN(n718) );
  XNOR2_X1 U766 ( .A(KEYINPUT124), .B(n718), .ZN(G69) );
  XOR2_X1 U767 ( .A(n720), .B(n719), .Z(n724) );
  XOR2_X1 U768 ( .A(n724), .B(n721), .Z(n722) );
  NOR2_X1 U769 ( .A1(G953), .A2(n722), .ZN(n723) );
  XNOR2_X1 U770 ( .A(KEYINPUT125), .B(n723), .ZN(n728) );
  XNOR2_X1 U771 ( .A(G227), .B(n724), .ZN(n725) );
  NAND2_X1 U772 ( .A1(n725), .A2(G900), .ZN(n726) );
  NAND2_X1 U773 ( .A1(n726), .A2(G953), .ZN(n727) );
  NAND2_X1 U774 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U775 ( .A(n729), .B(KEYINPUT126), .ZN(G72) );
  XNOR2_X1 U776 ( .A(G101), .B(n730), .ZN(G3) );
  XNOR2_X1 U777 ( .A(G110), .B(n731), .ZN(G12) );
  XOR2_X1 U778 ( .A(G122), .B(KEYINPUT127), .Z(n732) );
  XNOR2_X1 U779 ( .A(n733), .B(n732), .ZN(G24) );
  XOR2_X1 U780 ( .A(G119), .B(n734), .Z(G21) );
  XOR2_X1 U781 ( .A(G137), .B(n735), .Z(G39) );
  XOR2_X1 U782 ( .A(n736), .B(G131), .Z(G33) );
  XNOR2_X1 U783 ( .A(G134), .B(n737), .ZN(G36) );
endmodule

