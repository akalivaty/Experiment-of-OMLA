//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 0 0 1 1 1 1 0 1 1 1 1 1 1 1 0 1 1 1 0 1 0 0 0 0 1 0 0 1 0 0 1 0 1 1 1 1 0 1 0 1 1 1 1 1 1 1 1 0 1 0 1 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:48 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n536,
    new_n537, new_n538, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n575, new_n576, new_n577, new_n578,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n591, new_n592, new_n595, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT64), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(G2105), .ZN(new_n458));
  AND2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  OAI21_X1  g035(.A(new_n458), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(G137), .ZN(new_n462));
  INV_X1    g037(.A(G101), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n458), .A2(G2104), .ZN(new_n464));
  OAI22_X1  g039(.A1(new_n461), .A2(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g040(.A(G125), .B1(new_n459), .B2(new_n460), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n458), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n465), .A2(new_n468), .ZN(G160));
  NOR2_X1   g044(.A1(new_n459), .A2(new_n460), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n470), .A2(new_n458), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G124), .ZN(new_n472));
  XOR2_X1   g047(.A(new_n472), .B(KEYINPUT66), .Z(new_n473));
  OAI21_X1  g048(.A(KEYINPUT67), .B1(G100), .B2(G2105), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(new_n475));
  NOR3_X1   g050(.A1(KEYINPUT67), .A2(G100), .A3(G2105), .ZN(new_n476));
  OAI221_X1 g051(.A(G2104), .B1(G112), .B2(new_n458), .C1(new_n475), .C2(new_n476), .ZN(new_n477));
  XNOR2_X1  g052(.A(new_n477), .B(KEYINPUT68), .ZN(new_n478));
  INV_X1    g053(.A(new_n461), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  AND3_X1   g055(.A1(new_n473), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT69), .ZN(new_n482));
  XNOR2_X1  g057(.A(new_n481), .B(new_n482), .ZN(G162));
  OAI21_X1  g058(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(G114), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n484), .B1(new_n485), .B2(G2105), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n486), .B1(new_n471), .B2(G126), .ZN(new_n487));
  INV_X1    g062(.A(G138), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n488), .B1(KEYINPUT70), .B2(KEYINPUT4), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n479), .B(new_n489), .C1(KEYINPUT70), .C2(KEYINPUT4), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT70), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n491), .B(new_n492), .C1(new_n461), .C2(new_n488), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n487), .A2(new_n490), .A3(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(G164));
  INV_X1    g070(.A(G543), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT5), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n496), .B1(new_n497), .B2(KEYINPUT71), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT71), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n499), .A2(KEYINPUT5), .A3(G543), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n501), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n502));
  INV_X1    g077(.A(G651), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g079(.A(KEYINPUT6), .B(G651), .ZN(new_n505));
  AND3_X1   g080(.A1(new_n499), .A2(KEYINPUT5), .A3(G543), .ZN(new_n506));
  AOI21_X1  g081(.A(G543), .B1(new_n499), .B2(KEYINPUT5), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G88), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n505), .A2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G50), .ZN(new_n511));
  OAI22_X1  g086(.A1(new_n508), .A2(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n504), .A2(new_n512), .ZN(G166));
  INV_X1    g088(.A(new_n508), .ZN(new_n514));
  AND2_X1   g089(.A1(new_n514), .A2(G89), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n501), .A2(G63), .A3(G651), .ZN(new_n516));
  NAND3_X1  g091(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n517));
  XNOR2_X1  g092(.A(new_n517), .B(KEYINPUT7), .ZN(new_n518));
  INV_X1    g093(.A(G51), .ZN(new_n519));
  OAI211_X1 g094(.A(new_n516), .B(new_n518), .C1(new_n519), .C2(new_n510), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n515), .A2(new_n520), .ZN(G168));
  AOI22_X1  g096(.A1(new_n501), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n522), .A2(new_n503), .ZN(new_n523));
  INV_X1    g098(.A(G90), .ZN(new_n524));
  INV_X1    g099(.A(G52), .ZN(new_n525));
  OAI22_X1  g100(.A1(new_n508), .A2(new_n524), .B1(new_n510), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n523), .A2(new_n526), .ZN(G171));
  AOI22_X1  g102(.A1(new_n501), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n528), .A2(new_n503), .ZN(new_n529));
  XOR2_X1   g104(.A(KEYINPUT72), .B(G81), .Z(new_n530));
  INV_X1    g105(.A(G43), .ZN(new_n531));
  OAI22_X1  g106(.A1(new_n508), .A2(new_n530), .B1(new_n510), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G860), .ZN(G153));
  NAND4_X1  g109(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g110(.A1(G1), .A2(G3), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT73), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n537), .B(KEYINPUT8), .ZN(new_n538));
  NAND4_X1  g113(.A1(G319), .A2(G483), .A3(G661), .A4(new_n538), .ZN(G188));
  INV_X1    g114(.A(KEYINPUT74), .ZN(new_n540));
  AND3_X1   g115(.A1(new_n501), .A2(new_n540), .A3(new_n505), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n540), .B1(new_n501), .B2(new_n505), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G91), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n501), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n545), .A2(new_n503), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n505), .A2(G53), .A3(G543), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT9), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n544), .A2(new_n546), .A3(new_n548), .ZN(G299));
  INV_X1    g124(.A(G171), .ZN(G301));
  INV_X1    g125(.A(G168), .ZN(G286));
  INV_X1    g126(.A(G166), .ZN(G303));
  INV_X1    g127(.A(G49), .ZN(new_n553));
  OR3_X1    g128(.A1(new_n510), .A2(KEYINPUT75), .A3(new_n553), .ZN(new_n554));
  OAI21_X1  g129(.A(KEYINPUT75), .B1(new_n510), .B2(new_n553), .ZN(new_n555));
  OR2_X1    g130(.A1(new_n501), .A2(G74), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n554), .A2(new_n555), .B1(G651), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n543), .A2(G87), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n557), .A2(new_n558), .ZN(G288));
  NAND2_X1  g134(.A1(new_n508), .A2(KEYINPUT74), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n501), .A2(new_n540), .A3(new_n505), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n560), .A2(G86), .A3(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT76), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n560), .A2(KEYINPUT76), .A3(G86), .A4(new_n561), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n501), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n567));
  INV_X1    g142(.A(G48), .ZN(new_n568));
  OAI22_X1  g143(.A1(new_n567), .A2(new_n503), .B1(new_n568), .B2(new_n510), .ZN(new_n569));
  INV_X1    g144(.A(new_n569), .ZN(new_n570));
  AOI21_X1  g145(.A(KEYINPUT77), .B1(new_n566), .B2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT77), .ZN(new_n572));
  AOI211_X1 g147(.A(new_n572), .B(new_n569), .C1(new_n564), .C2(new_n565), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n571), .A2(new_n573), .ZN(G305));
  AOI22_X1  g149(.A1(new_n501), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n575));
  OR2_X1    g150(.A1(new_n575), .A2(new_n503), .ZN(new_n576));
  INV_X1    g151(.A(new_n510), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n514), .A2(G85), .B1(new_n577), .B2(G47), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n576), .A2(new_n578), .ZN(G290));
  NAND2_X1  g154(.A1(G301), .A2(G868), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n501), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n581));
  INV_X1    g156(.A(G54), .ZN(new_n582));
  OAI22_X1  g157(.A1(new_n581), .A2(new_n503), .B1(new_n582), .B2(new_n510), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n560), .A2(G92), .A3(new_n561), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT10), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND4_X1  g161(.A1(new_n560), .A2(KEYINPUT10), .A3(G92), .A4(new_n561), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n583), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n580), .B1(new_n588), .B2(G868), .ZN(G321));
  XNOR2_X1  g164(.A(G321), .B(KEYINPUT78), .ZN(G284));
  NAND2_X1  g165(.A1(G286), .A2(G868), .ZN(new_n591));
  AND3_X1   g166(.A1(new_n544), .A2(new_n546), .A3(new_n548), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n592), .B2(G868), .ZN(G297));
  OAI21_X1  g168(.A(new_n591), .B1(new_n592), .B2(G868), .ZN(G280));
  INV_X1    g169(.A(G559), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n588), .B1(new_n595), .B2(G860), .ZN(G148));
  OR2_X1    g171(.A1(new_n529), .A2(new_n532), .ZN(new_n597));
  INV_X1    g172(.A(G868), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n586), .A2(new_n587), .ZN(new_n600));
  INV_X1    g175(.A(new_n583), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n602), .A2(G559), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n599), .B1(new_n603), .B2(new_n598), .ZN(G323));
  XNOR2_X1  g179(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g180(.A1(new_n470), .A2(new_n464), .ZN(new_n606));
  XNOR2_X1  g181(.A(KEYINPUT79), .B(KEYINPUT12), .ZN(new_n607));
  XOR2_X1   g182(.A(new_n606), .B(new_n607), .Z(new_n608));
  XOR2_X1   g183(.A(KEYINPUT80), .B(KEYINPUT13), .Z(new_n609));
  XNOR2_X1  g184(.A(new_n608), .B(new_n609), .ZN(new_n610));
  XNOR2_X1  g185(.A(KEYINPUT81), .B(G2100), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT82), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n471), .A2(G123), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n479), .A2(G135), .ZN(new_n615));
  OAI21_X1  g190(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n616));
  INV_X1    g191(.A(G111), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n616), .A2(KEYINPUT83), .B1(new_n617), .B2(G2105), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n618), .B1(KEYINPUT83), .B2(new_n616), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n614), .A2(new_n615), .A3(new_n619), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(G2096), .Z(new_n621));
  OAI211_X1 g196(.A(new_n613), .B(new_n621), .C1(new_n611), .C2(new_n610), .ZN(G156));
  XOR2_X1   g197(.A(KEYINPUT15), .B(G2435), .Z(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(G2438), .ZN(new_n624));
  XNOR2_X1  g199(.A(G2427), .B(G2430), .ZN(new_n625));
  INV_X1    g200(.A(KEYINPUT85), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  OR2_X1    g202(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n624), .A2(new_n627), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n628), .A2(KEYINPUT14), .A3(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(KEYINPUT84), .B(KEYINPUT16), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(G2451), .B(G2454), .Z(new_n633));
  XNOR2_X1  g208(.A(G2443), .B(G2446), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n632), .B(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(G1341), .B(G1348), .Z(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n638), .A2(G14), .ZN(new_n639));
  OR3_X1    g214(.A1(new_n636), .A2(KEYINPUT86), .A3(new_n637), .ZN(new_n640));
  OAI21_X1  g215(.A(KEYINPUT86), .B1(new_n636), .B2(new_n637), .ZN(new_n641));
  AOI21_X1  g216(.A(new_n639), .B1(new_n640), .B2(new_n641), .ZN(G401));
  XNOR2_X1  g217(.A(G2067), .B(G2678), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT87), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2072), .B(G2078), .ZN(new_n645));
  XOR2_X1   g220(.A(G2084), .B(G2090), .Z(new_n646));
  NAND3_X1  g221(.A1(new_n644), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT88), .B(KEYINPUT18), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n644), .A2(new_n646), .ZN(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n645), .B1(new_n651), .B2(KEYINPUT17), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n644), .A2(new_n646), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n645), .A2(KEYINPUT17), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n653), .B1(new_n650), .B2(new_n654), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n649), .B1(new_n652), .B2(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G2096), .B(G2100), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(G227));
  XOR2_X1   g233(.A(G1971), .B(G1976), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT19), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1956), .B(G2474), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1961), .B(G1966), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AND2_X1   g238(.A1(new_n661), .A2(new_n662), .ZN(new_n664));
  NOR3_X1   g239(.A1(new_n660), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n660), .A2(new_n663), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(KEYINPUT20), .Z(new_n667));
  AOI211_X1 g242(.A(new_n665), .B(new_n667), .C1(new_n660), .C2(new_n664), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT89), .ZN(new_n669));
  XOR2_X1   g244(.A(G1981), .B(G1986), .Z(new_n670));
  XNOR2_X1  g245(.A(G1991), .B(G1996), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n669), .B(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(G229));
  NOR2_X1   g251(.A1(G16), .A2(G23), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT93), .ZN(new_n678));
  INV_X1    g253(.A(G16), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n678), .B1(G288), .B2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT33), .B(G1976), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT92), .B(G16), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n684), .A2(G22), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n685), .B1(G166), .B2(new_n684), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(G1971), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n682), .A2(new_n687), .ZN(new_n688));
  AND2_X1   g263(.A1(new_n679), .A2(G6), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n689), .B1(G305), .B2(G16), .ZN(new_n690));
  XOR2_X1   g265(.A(KEYINPUT32), .B(G1981), .Z(new_n691));
  AND2_X1   g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n690), .A2(new_n691), .ZN(new_n693));
  NOR3_X1   g268(.A1(new_n688), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(KEYINPUT34), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n694), .A2(new_n695), .ZN(new_n697));
  INV_X1    g272(.A(G25), .ZN(new_n698));
  OR3_X1    g273(.A1(new_n698), .A2(KEYINPUT90), .A3(G29), .ZN(new_n699));
  OAI21_X1  g274(.A(KEYINPUT90), .B1(new_n698), .B2(G29), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n471), .A2(G119), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n479), .A2(G131), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n458), .A2(G107), .ZN(new_n703));
  OAI21_X1  g278(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n704));
  OAI211_X1 g279(.A(new_n701), .B(new_n702), .C1(new_n703), .C2(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(KEYINPUT91), .ZN(new_n706));
  OR2_X1    g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n705), .A2(new_n706), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(G29), .ZN(new_n711));
  OAI211_X1 g286(.A(new_n699), .B(new_n700), .C1(new_n710), .C2(new_n711), .ZN(new_n712));
  XOR2_X1   g287(.A(KEYINPUT35), .B(G1991), .Z(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n684), .A2(G24), .ZN(new_n715));
  INV_X1    g290(.A(G290), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n715), .B1(new_n716), .B2(new_n684), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(G1986), .Z(new_n718));
  NAND4_X1  g293(.A1(new_n696), .A2(new_n697), .A3(new_n714), .A4(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT36), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n683), .A2(G20), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT23), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(new_n592), .B2(new_n679), .ZN(new_n724));
  INV_X1    g299(.A(G1956), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  NOR2_X1   g301(.A1(G4), .A2(G16), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(new_n588), .B2(G16), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(G1348), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n684), .A2(G19), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(new_n533), .B2(new_n684), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(G1341), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n711), .A2(G26), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT28), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n471), .A2(G128), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n479), .A2(G140), .ZN(new_n736));
  OR2_X1    g311(.A1(G104), .A2(G2105), .ZN(new_n737));
  OAI211_X1 g312(.A(new_n737), .B(G2104), .C1(G116), .C2(new_n458), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n735), .A2(new_n736), .A3(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(new_n739), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n734), .B1(new_n740), .B2(new_n711), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(G2067), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n732), .A2(new_n742), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n728), .A2(G1348), .ZN(new_n744));
  NAND4_X1  g319(.A1(new_n726), .A2(new_n729), .A3(new_n743), .A4(new_n744), .ZN(new_n745));
  NOR2_X1   g320(.A1(G29), .A2(G35), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(G162), .B2(G29), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT29), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n745), .B1(new_n748), .B2(G2090), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G2090), .B2(new_n748), .ZN(new_n750));
  INV_X1    g325(.A(G34), .ZN(new_n751));
  AND2_X1   g326(.A1(new_n751), .A2(KEYINPUT24), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n751), .A2(KEYINPUT24), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n711), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G160), .B2(new_n711), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT95), .Z(new_n756));
  NOR2_X1   g331(.A1(new_n756), .A2(G2084), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n756), .A2(G2084), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n711), .A2(G33), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n458), .A2(G103), .A3(G2104), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT25), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(G139), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n762), .B1(new_n763), .B2(new_n461), .ZN(new_n764));
  OAI21_X1  g339(.A(G127), .B1(new_n459), .B2(new_n460), .ZN(new_n765));
  NAND2_X1  g340(.A1(G115), .A2(G2104), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n458), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n764), .A2(new_n767), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n759), .B1(new_n768), .B2(new_n711), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT94), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n758), .B1(G2072), .B2(new_n770), .ZN(new_n771));
  AOI211_X1 g346(.A(new_n757), .B(new_n771), .C1(G2072), .C2(new_n770), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n711), .A2(G32), .ZN(new_n773));
  NAND3_X1  g348(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT26), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(new_n471), .B2(G129), .ZN(new_n776));
  INV_X1    g351(.A(new_n464), .ZN(new_n777));
  AOI22_X1  g352(.A1(new_n479), .A2(G141), .B1(G105), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT96), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n773), .B1(new_n780), .B2(new_n711), .ZN(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT27), .B(G1996), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(G171), .A2(new_n679), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(G5), .B2(new_n679), .ZN(new_n785));
  INV_X1    g360(.A(G1961), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  AND2_X1   g362(.A1(new_n785), .A2(new_n786), .ZN(new_n788));
  INV_X1    g363(.A(G2078), .ZN(new_n789));
  NAND2_X1  g364(.A1(G164), .A2(G29), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G27), .B2(G29), .ZN(new_n791));
  AOI211_X1 g366(.A(new_n787), .B(new_n788), .C1(new_n789), .C2(new_n791), .ZN(new_n792));
  XNOR2_X1  g367(.A(KEYINPUT31), .B(G11), .ZN(new_n793));
  INV_X1    g368(.A(KEYINPUT30), .ZN(new_n794));
  AND2_X1   g369(.A1(new_n794), .A2(G28), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n711), .B1(new_n794), .B2(G28), .ZN(new_n796));
  OAI221_X1 g371(.A(new_n793), .B1(new_n795), .B2(new_n796), .C1(new_n620), .C2(new_n711), .ZN(new_n797));
  NOR2_X1   g372(.A1(G168), .A2(new_n679), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(new_n679), .B2(G21), .ZN(new_n799));
  INV_X1    g374(.A(G1966), .ZN(new_n800));
  OAI22_X1  g375(.A1(new_n799), .A2(new_n800), .B1(new_n791), .B2(new_n789), .ZN(new_n801));
  AOI211_X1 g376(.A(new_n797), .B(new_n801), .C1(new_n800), .C2(new_n799), .ZN(new_n802));
  NAND4_X1  g377(.A1(new_n772), .A2(new_n783), .A3(new_n792), .A4(new_n802), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT97), .ZN(new_n804));
  NOR3_X1   g379(.A1(new_n721), .A2(new_n750), .A3(new_n804), .ZN(G311));
  INV_X1    g380(.A(G311), .ZN(G150));
  AOI22_X1  g381(.A1(new_n514), .A2(G93), .B1(new_n577), .B2(G55), .ZN(new_n807));
  INV_X1    g382(.A(KEYINPUT98), .ZN(new_n808));
  AND2_X1   g383(.A1(new_n501), .A2(G67), .ZN(new_n809));
  AND2_X1   g384(.A1(G80), .A2(G543), .ZN(new_n810));
  OAI211_X1 g385(.A(new_n808), .B(G651), .C1(new_n809), .C2(new_n810), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n810), .B1(new_n501), .B2(G67), .ZN(new_n812));
  OAI21_X1  g387(.A(KEYINPUT98), .B1(new_n812), .B2(new_n503), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n807), .A2(new_n811), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n814), .A2(G860), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(KEYINPUT37), .Z(new_n816));
  NAND2_X1  g391(.A1(new_n588), .A2(G559), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT38), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n814), .A2(new_n597), .ZN(new_n819));
  NAND4_X1  g394(.A1(new_n533), .A2(new_n811), .A3(new_n813), .A4(new_n807), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n818), .B(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n823), .A2(KEYINPUT39), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT99), .ZN(new_n825));
  INV_X1    g400(.A(G860), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(new_n823), .B2(KEYINPUT39), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n816), .B1(new_n825), .B2(new_n827), .ZN(G145));
  XNOR2_X1  g403(.A(new_n481), .B(KEYINPUT69), .ZN(new_n829));
  INV_X1    g404(.A(G160), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g406(.A1(G162), .A2(G160), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(new_n620), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n620), .B1(new_n831), .B2(new_n832), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AOI22_X1  g412(.A1(G130), .A2(new_n471), .B1(new_n479), .B2(G142), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT100), .ZN(new_n839));
  NOR3_X1   g414(.A1(new_n839), .A2(new_n458), .A3(G118), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n839), .B1(new_n458), .B2(G118), .ZN(new_n841));
  OAI211_X1 g416(.A(new_n841), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n838), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n709), .B(new_n843), .ZN(new_n844));
  OR2_X1    g419(.A1(new_n844), .A2(new_n608), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n608), .ZN(new_n846));
  AND2_X1   g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NOR3_X1   g422(.A1(new_n780), .A2(new_n767), .A3(new_n764), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n494), .B(new_n739), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n768), .A2(new_n779), .ZN(new_n850));
  OR3_X1    g425(.A1(new_n848), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n849), .B1(new_n848), .B2(new_n850), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n847), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n845), .A2(new_n846), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n855), .B1(new_n852), .B2(new_n851), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n837), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(G37), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  OAI21_X1  g434(.A(KEYINPUT101), .B1(new_n847), .B2(new_n853), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT101), .ZN(new_n861));
  NAND4_X1  g436(.A1(new_n855), .A2(new_n861), .A3(new_n852), .A4(new_n851), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n847), .A2(new_n853), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n864), .A2(new_n835), .A3(new_n836), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g441(.A(KEYINPUT102), .B1(new_n859), .B2(new_n866), .ZN(new_n867));
  OR2_X1    g442(.A1(new_n863), .A2(new_n865), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n847), .B(new_n853), .ZN(new_n869));
  AOI21_X1  g444(.A(G37), .B1(new_n869), .B2(new_n837), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT102), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n868), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  AND3_X1   g447(.A1(new_n867), .A2(KEYINPUT40), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(KEYINPUT40), .B1(new_n867), .B2(new_n872), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n873), .A2(new_n874), .ZN(G395));
  NAND2_X1  g450(.A1(new_n814), .A2(new_n598), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n566), .A2(new_n570), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(new_n572), .ZN(new_n878));
  OR3_X1    g453(.A1(new_n504), .A2(new_n512), .A3(KEYINPUT105), .ZN(new_n879));
  OAI21_X1  g454(.A(KEYINPUT105), .B1(new_n504), .B2(new_n512), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n569), .B1(new_n564), .B2(new_n565), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(KEYINPUT77), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n878), .A2(new_n882), .A3(new_n884), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n881), .B1(new_n571), .B2(new_n573), .ZN(new_n886));
  XNOR2_X1  g461(.A(G288), .B(G290), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT106), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND4_X1  g465(.A1(new_n885), .A2(new_n886), .A3(KEYINPUT106), .A4(new_n887), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT107), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n885), .A2(new_n886), .ZN(new_n894));
  INV_X1    g469(.A(new_n887), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n893), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  AOI211_X1 g471(.A(KEYINPUT107), .B(new_n887), .C1(new_n885), .C2(new_n886), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n892), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n898), .B(KEYINPUT42), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n603), .B(new_n821), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n602), .A2(KEYINPUT103), .A3(new_n592), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT103), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n903), .B1(new_n588), .B2(G299), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n588), .A2(G299), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n902), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n901), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n907), .B(KEYINPUT104), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n906), .A2(KEYINPUT41), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT41), .ZN(new_n910));
  NAND4_X1  g485(.A1(new_n902), .A2(new_n904), .A3(new_n910), .A4(new_n905), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n900), .A2(new_n909), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n908), .A2(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n899), .B(new_n913), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n876), .B1(new_n914), .B2(new_n598), .ZN(G295));
  OAI21_X1  g490(.A(new_n876), .B1(new_n914), .B2(new_n598), .ZN(G331));
  AOI21_X1  g491(.A(new_n882), .B1(new_n878), .B2(new_n884), .ZN(new_n917));
  NOR3_X1   g492(.A1(new_n571), .A2(new_n573), .A3(new_n881), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n895), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(KEYINPUT107), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n894), .A2(new_n893), .A3(new_n895), .ZN(new_n921));
  AOI22_X1  g496(.A1(new_n920), .A2(new_n921), .B1(new_n890), .B2(new_n891), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n821), .A2(G171), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n819), .A2(new_n820), .A3(G301), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n923), .A2(G168), .A3(new_n924), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n819), .A2(new_n820), .A3(G301), .ZN(new_n926));
  AOI21_X1  g501(.A(G301), .B1(new_n819), .B2(new_n820), .ZN(new_n927));
  OAI21_X1  g502(.A(G286), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n909), .A2(new_n911), .A3(new_n925), .A4(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n925), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(new_n906), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(KEYINPUT108), .B1(new_n922), .B2(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(G37), .B1(new_n922), .B2(new_n932), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT108), .ZN(new_n935));
  AND2_X1   g510(.A1(new_n929), .A2(new_n931), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n898), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n933), .A2(new_n934), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(KEYINPUT43), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT43), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n933), .A2(new_n934), .A3(new_n937), .A4(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n939), .A2(KEYINPUT109), .A3(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT109), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n938), .A2(new_n943), .A3(KEYINPUT43), .ZN(new_n944));
  AOI21_X1  g519(.A(KEYINPUT44), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n939), .A2(KEYINPUT110), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(new_n941), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT110), .ZN(new_n948));
  OR3_X1    g523(.A1(new_n938), .A2(new_n948), .A3(KEYINPUT43), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n945), .B1(new_n950), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g526(.A(G1384), .ZN(new_n952));
  AOI21_X1  g527(.A(KEYINPUT45), .B1(new_n494), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(G40), .ZN(new_n954));
  NOR3_X1   g529(.A1(new_n465), .A2(new_n468), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n956), .A2(G1996), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(KEYINPUT46), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT125), .ZN(new_n959));
  XNOR2_X1  g534(.A(new_n958), .B(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(G2067), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n739), .B(new_n961), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n962), .B(KEYINPUT112), .ZN(new_n963));
  INV_X1    g538(.A(new_n779), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n956), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n957), .A2(KEYINPUT46), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n960), .A2(new_n967), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n968), .B(KEYINPUT47), .ZN(new_n969));
  INV_X1    g544(.A(G1996), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n963), .A2(new_n970), .ZN(new_n971));
  AOI22_X1  g546(.A1(new_n965), .A2(new_n971), .B1(new_n780), .B2(new_n957), .ZN(new_n972));
  INV_X1    g547(.A(new_n956), .ZN(new_n973));
  AND2_X1   g548(.A1(new_n710), .A2(new_n713), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n710), .A2(new_n713), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n973), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  OR3_X1    g551(.A1(new_n956), .A2(G1986), .A3(G290), .ZN(new_n977));
  XNOR2_X1  g552(.A(new_n977), .B(KEYINPUT48), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n972), .A2(new_n976), .A3(new_n978), .ZN(new_n979));
  XOR2_X1   g554(.A(new_n974), .B(KEYINPUT124), .Z(new_n980));
  AOI22_X1  g555(.A1(new_n980), .A2(new_n972), .B1(new_n961), .B2(new_n740), .ZN(new_n981));
  OAI211_X1 g556(.A(new_n969), .B(new_n979), .C1(new_n956), .C2(new_n981), .ZN(new_n982));
  XOR2_X1   g557(.A(new_n982), .B(KEYINPUT126), .Z(new_n983));
  NAND2_X1  g558(.A1(G303), .A2(G8), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n984), .B(KEYINPUT55), .ZN(new_n985));
  INV_X1    g560(.A(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n953), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n494), .A2(KEYINPUT45), .A3(new_n952), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n987), .A2(new_n988), .A3(new_n955), .ZN(new_n989));
  INV_X1    g564(.A(G1971), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT50), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n494), .A2(new_n994), .A3(new_n952), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n993), .A2(new_n955), .A3(new_n995), .ZN(new_n996));
  OAI22_X1  g571(.A1(new_n992), .A2(KEYINPUT113), .B1(G2090), .B2(new_n996), .ZN(new_n997));
  AND2_X1   g572(.A1(new_n992), .A2(KEYINPUT113), .ZN(new_n998));
  OAI211_X1 g573(.A(G8), .B(new_n986), .C1(new_n997), .C2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n494), .A2(new_n955), .A3(new_n952), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(G8), .ZN(new_n1002));
  INV_X1    g577(.A(new_n1002), .ZN(new_n1003));
  XOR2_X1   g578(.A(KEYINPUT114), .B(G1981), .Z(new_n1004));
  NAND2_X1  g579(.A1(new_n883), .A2(new_n1004), .ZN(new_n1005));
  AND2_X1   g580(.A1(new_n514), .A2(G86), .ZN(new_n1006));
  OAI21_X1  g581(.A(G1981), .B1(new_n569), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1003), .B1(new_n1009), .B2(KEYINPUT49), .ZN(new_n1010));
  AND3_X1   g585(.A1(new_n1005), .A2(KEYINPUT49), .A3(new_n1007), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(G1976), .ZN(new_n1013));
  AOI21_X1  g588(.A(KEYINPUT52), .B1(G288), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(G288), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1002), .B1(new_n1015), .B2(G1976), .ZN(new_n1016));
  MUX2_X1   g591(.A(KEYINPUT52), .B(new_n1014), .S(new_n1016), .Z(new_n1017));
  NOR2_X1   g592(.A1(new_n1012), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1015), .A2(new_n1013), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1005), .B1(new_n1012), .B2(new_n1019), .ZN(new_n1020));
  XOR2_X1   g595(.A(new_n1002), .B(KEYINPUT115), .Z(new_n1021));
  AOI22_X1  g596(.A1(new_n1000), .A2(new_n1018), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  AND2_X1   g597(.A1(new_n999), .A2(new_n1018), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT116), .ZN(new_n1024));
  OR3_X1    g599(.A1(new_n996), .A2(new_n1024), .A3(G2084), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1024), .B1(new_n996), .B2(G2084), .ZN(new_n1026));
  INV_X1    g601(.A(new_n989), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n1025), .B(new_n1026), .C1(G1966), .C2(new_n1027), .ZN(new_n1028));
  AND3_X1   g603(.A1(new_n1028), .A2(G8), .A3(G168), .ZN(new_n1029));
  OAI21_X1  g604(.A(G8), .B1(new_n997), .B2(new_n998), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(new_n985), .ZN(new_n1031));
  AND4_X1   g606(.A1(KEYINPUT63), .A2(new_n1023), .A3(new_n1029), .A4(new_n1031), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n996), .A2(G2090), .ZN(new_n1033));
  OAI21_X1  g608(.A(G8), .B1(new_n992), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(new_n985), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1029), .A2(new_n1035), .A3(new_n999), .A4(new_n1018), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT63), .ZN(new_n1037));
  AND2_X1   g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1022), .B1(new_n1032), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(G8), .ZN(new_n1040));
  NOR2_X1   g615(.A1(G168), .A2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1041), .B1(new_n1028), .B2(G8), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1041), .ZN(new_n1043));
  AOI21_X1  g618(.A(KEYINPUT51), .B1(new_n1043), .B2(KEYINPUT123), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1044), .ZN(new_n1045));
  OR2_X1    g620(.A1(new_n1042), .A2(new_n1045), .ZN(new_n1046));
  AOI22_X1  g621(.A1(new_n1042), .A2(new_n1045), .B1(new_n1041), .B2(new_n1028), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT62), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n989), .A2(G2078), .ZN(new_n1049));
  OR2_X1    g624(.A1(new_n1049), .A2(KEYINPUT53), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n996), .A2(new_n786), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1049), .A2(KEYINPUT53), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1050), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  AND2_X1   g628(.A1(new_n1053), .A2(G171), .ZN(new_n1054));
  AOI22_X1  g629(.A1(new_n1046), .A2(new_n1047), .B1(new_n1048), .B2(new_n1054), .ZN(new_n1055));
  XNOR2_X1  g630(.A(G299), .B(KEYINPUT57), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  XNOR2_X1  g632(.A(KEYINPUT56), .B(G2072), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n989), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n996), .A2(KEYINPUT117), .A3(new_n725), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(KEYINPUT117), .B1(new_n996), .B2(new_n725), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n1057), .B(new_n1061), .C1(new_n1063), .C2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(G1348), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n996), .A2(new_n1067), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n494), .A2(new_n955), .A3(new_n952), .A4(new_n961), .ZN(new_n1069));
  XNOR2_X1  g644(.A(new_n1069), .B(KEYINPUT118), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n602), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1061), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(new_n1056), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1071), .B1(new_n1073), .B2(KEYINPUT119), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1064), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(new_n1062), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1057), .B1(new_n1076), .B2(new_n1061), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT119), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1066), .B1(new_n1074), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1065), .A2(KEYINPUT61), .ZN(new_n1081));
  AND3_X1   g656(.A1(new_n1068), .A2(new_n602), .A3(new_n1070), .ZN(new_n1082));
  OAI21_X1  g657(.A(KEYINPUT60), .B1(new_n1082), .B2(new_n1071), .ZN(new_n1083));
  XOR2_X1   g658(.A(KEYINPUT120), .B(G1996), .Z(new_n1084));
  NAND4_X1  g659(.A1(new_n987), .A2(new_n988), .A3(new_n955), .A4(new_n1084), .ZN(new_n1085));
  XOR2_X1   g660(.A(KEYINPUT58), .B(G1341), .Z(new_n1086));
  NAND2_X1  g661(.A1(new_n1001), .A2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n597), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n1089));
  XNOR2_X1  g664(.A(new_n1088), .B(new_n1089), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n602), .A2(KEYINPUT60), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1068), .A2(new_n1070), .A3(new_n1091), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1081), .A2(new_n1083), .A3(new_n1090), .A4(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT122), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT61), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1095), .B1(new_n1077), .B2(new_n1066), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1093), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  OAI211_X1 g672(.A(KEYINPUT122), .B(new_n1095), .C1(new_n1077), .C2(new_n1066), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1080), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1053), .A2(G171), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT54), .ZN(new_n1101));
  OR3_X1    g676(.A1(new_n1054), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1101), .B1(new_n1054), .B2(new_n1100), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1055), .B1(new_n1099), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1023), .A2(new_n1035), .ZN(new_n1106));
  AND2_X1   g681(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1054), .A2(KEYINPUT62), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1106), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1039), .B1(new_n1105), .B2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n973), .A2(G1986), .A3(G290), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n977), .A2(new_n1111), .ZN(new_n1112));
  XOR2_X1   g687(.A(new_n1112), .B(KEYINPUT111), .Z(new_n1113));
  NAND3_X1  g688(.A1(new_n1113), .A2(new_n972), .A3(new_n976), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n983), .B1(new_n1110), .B2(new_n1114), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g690(.A(G319), .ZN(new_n1117));
  NOR2_X1   g691(.A1(G227), .A2(new_n1117), .ZN(new_n1118));
  AND2_X1   g692(.A1(new_n640), .A2(new_n641), .ZN(new_n1119));
  OAI211_X1 g693(.A(KEYINPUT127), .B(new_n1118), .C1(new_n1119), .C2(new_n639), .ZN(new_n1120));
  INV_X1    g694(.A(KEYINPUT127), .ZN(new_n1121));
  INV_X1    g695(.A(new_n1118), .ZN(new_n1122));
  OAI21_X1  g696(.A(new_n1121), .B1(G401), .B2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g697(.A1(new_n1120), .A2(new_n675), .A3(new_n1123), .ZN(new_n1124));
  AOI21_X1  g698(.A(new_n1124), .B1(new_n867), .B2(new_n872), .ZN(new_n1125));
  AND3_X1   g699(.A1(new_n1125), .A2(new_n944), .A3(new_n942), .ZN(G308));
  NAND3_X1  g700(.A1(new_n1125), .A2(new_n944), .A3(new_n942), .ZN(G225));
endmodule


