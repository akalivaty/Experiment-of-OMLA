//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 0 1 1 0 1 0 0 0 1 1 0 0 1 0 1 0 0 0 0 1 0 0 0 0 0 0 0 1 1 0 0 0 0 0 1 1 1 1 0 0 1 0 0 1 1 1 1 1 1 1 0 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:01 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1274, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(new_n204));
  XOR2_X1   g0004(.A(new_n204), .B(KEYINPUT64), .Z(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0006(.A1(G77), .A2(G244), .B1(G87), .B2(G250), .ZN(new_n207));
  INV_X1    g0007(.A(G116), .ZN(new_n208));
  INV_X1    g0008(.A(G270), .ZN(new_n209));
  OAI21_X1  g0009(.A(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G68), .A2(G238), .ZN(new_n212));
  INV_X1    g0012(.A(G226), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n211), .B(new_n212), .C1(new_n202), .C2(new_n213), .ZN(new_n214));
  AOI211_X1 g0014(.A(new_n210), .B(new_n214), .C1(G97), .C2(G257), .ZN(new_n215));
  AOI21_X1  g0015(.A(new_n215), .B1(G1), .B2(G20), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT1), .Z(new_n217));
  OAI21_X1  g0017(.A(G50), .B1(G58), .B2(G68), .ZN(new_n218));
  INV_X1    g0018(.A(G20), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G13), .ZN(new_n220));
  NOR3_X1   g0020(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(G1), .ZN(new_n222));
  NOR3_X1   g0022(.A1(new_n222), .A2(new_n219), .A3(G13), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n223), .B(G250), .C1(G257), .C2(G264), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT0), .Z(new_n225));
  NOR3_X1   g0025(.A1(new_n217), .A2(new_n221), .A3(new_n225), .ZN(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(KEYINPUT2), .B(G226), .ZN(new_n229));
  XOR2_X1   g0029(.A(new_n228), .B(new_n229), .Z(new_n230));
  XOR2_X1   g0030(.A(G250), .B(G257), .Z(new_n231));
  XNOR2_X1  g0031(.A(G264), .B(G270), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n230), .B(new_n233), .Z(G358));
  XOR2_X1   g0034(.A(G68), .B(G77), .Z(new_n235));
  XNOR2_X1  g0035(.A(G50), .B(G58), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G351));
  NAND3_X1  g0041(.A1(new_n222), .A2(G13), .A3(G20), .ZN(new_n242));
  NOR2_X1   g0042(.A1(new_n242), .A2(G97), .ZN(new_n243));
  INV_X1    g0043(.A(new_n243), .ZN(new_n244));
  INV_X1    g0044(.A(new_n242), .ZN(new_n245));
  NAND3_X1  g0045(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(new_n220), .ZN(new_n247));
  NOR2_X1   g0047(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(G33), .ZN(new_n249));
  OAI21_X1  g0049(.A(new_n248), .B1(G1), .B2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G97), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  NOR2_X1   g0053(.A1(G20), .A2(G33), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G77), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT6), .ZN(new_n258));
  INV_X1    g0058(.A(G107), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n251), .A2(new_n259), .ZN(new_n260));
  NOR2_X1   g0060(.A1(G97), .A2(G107), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n258), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n259), .A2(KEYINPUT6), .A3(G97), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n219), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT74), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n265), .B1(new_n249), .B2(KEYINPUT3), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n249), .A2(KEYINPUT3), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT3), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n268), .A2(KEYINPUT74), .A3(G33), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n266), .A2(new_n267), .A3(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n270), .A2(KEYINPUT7), .A3(new_n219), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT7), .ZN(new_n272));
  XNOR2_X1  g0072(.A(KEYINPUT3), .B(G33), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n272), .B1(new_n273), .B2(G20), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n271), .A2(new_n274), .ZN(new_n275));
  AOI211_X1 g0075(.A(new_n257), .B(new_n264), .C1(new_n275), .C2(G107), .ZN(new_n276));
  INV_X1    g0076(.A(new_n247), .ZN(new_n277));
  OAI211_X1 g0077(.A(new_n244), .B(new_n253), .C1(new_n276), .C2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n268), .A2(G33), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n267), .A2(new_n280), .A3(G244), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT4), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(G33), .A2(G283), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n282), .A2(G1698), .ZN(new_n285));
  NAND4_X1  g0085(.A1(new_n285), .A2(new_n267), .A3(new_n280), .A4(G244), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n283), .A2(new_n284), .A3(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G1698), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n267), .A2(new_n280), .A3(G250), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n288), .B1(new_n289), .B2(KEYINPUT4), .ZN(new_n290));
  OAI21_X1  g0090(.A(KEYINPUT77), .B1(new_n287), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(G33), .A2(G41), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n292), .A2(G1), .A3(G13), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n289), .A2(KEYINPUT4), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(G1698), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT77), .ZN(new_n297));
  AOI22_X1  g0097(.A1(new_n281), .A2(new_n282), .B1(G33), .B2(G283), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n296), .A2(new_n297), .A3(new_n298), .A4(new_n286), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n291), .A2(new_n294), .A3(new_n299), .ZN(new_n300));
  XNOR2_X1  g0100(.A(KEYINPUT5), .B(G41), .ZN(new_n301));
  INV_X1    g0101(.A(G45), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n302), .A2(G1), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n304), .A2(G257), .A3(new_n293), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n301), .A2(G274), .A3(new_n303), .ZN(new_n306));
  AND2_X1   g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n300), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(G200), .ZN(new_n309));
  INV_X1    g0109(.A(G190), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n279), .B(new_n309), .C1(new_n310), .C2(new_n308), .ZN(new_n311));
  AND2_X1   g0111(.A1(new_n300), .A2(new_n307), .ZN(new_n312));
  INV_X1    g0112(.A(G179), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G169), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n308), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n314), .A2(new_n278), .A3(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT19), .ZN(new_n318));
  INV_X1    g0118(.A(G87), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n319), .A2(new_n251), .A3(new_n259), .ZN(new_n320));
  NAND2_X1  g0120(.A1(G33), .A2(G97), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(new_n219), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n318), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  NOR3_X1   g0123(.A1(new_n321), .A2(KEYINPUT19), .A3(G20), .ZN(new_n324));
  INV_X1    g0124(.A(G68), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n267), .A2(new_n280), .A3(new_n219), .ZN(new_n326));
  OAI22_X1  g0126(.A1(new_n323), .A2(new_n324), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT79), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  OAI221_X1 g0129(.A(KEYINPUT79), .B1(new_n326), .B2(new_n325), .C1(new_n323), .C2(new_n324), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n329), .A2(new_n247), .A3(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT15), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(new_n319), .ZN(new_n333));
  NAND2_X1  g0133(.A1(KEYINPUT15), .A2(G87), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(new_n245), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n331), .B(new_n336), .C1(new_n319), .C2(new_n250), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n267), .A2(new_n280), .A3(G238), .A4(new_n288), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT78), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND4_X1  g0140(.A1(new_n273), .A2(KEYINPUT78), .A3(G238), .A4(new_n288), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n249), .A2(new_n208), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n273), .A2(G244), .A3(G1698), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n340), .A2(new_n341), .A3(new_n343), .A4(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(new_n294), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n293), .B(G250), .C1(G1), .C2(new_n302), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n303), .A2(G274), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n346), .A2(new_n350), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n351), .A2(new_n310), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n349), .B1(new_n345), .B2(new_n294), .ZN(new_n353));
  INV_X1    g0153(.A(G200), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  OR3_X1    g0155(.A1(new_n337), .A2(new_n352), .A3(new_n355), .ZN(new_n356));
  AND3_X1   g0156(.A1(new_n311), .A2(new_n317), .A3(new_n356), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n242), .A2(G77), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n333), .A2(new_n219), .A3(G33), .A4(new_n334), .ZN(new_n359));
  NAND2_X1  g0159(.A1(G20), .A2(G77), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT8), .ZN(new_n361));
  INV_X1    g0161(.A(G58), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(KEYINPUT8), .A2(G58), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n363), .A2(new_n254), .A3(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n359), .A2(new_n360), .A3(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n358), .B1(new_n366), .B2(new_n247), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n247), .B1(new_n222), .B2(G20), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(G77), .ZN(new_n369));
  AOI21_X1  g0169(.A(KEYINPUT68), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n367), .A2(KEYINPUT68), .A3(new_n369), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n222), .B1(G41), .B2(G45), .ZN(new_n374));
  INV_X1    g0174(.A(G274), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n293), .A2(new_n374), .ZN(new_n378));
  INV_X1    g0178(.A(G244), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n377), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n267), .A2(new_n280), .A3(G232), .A4(new_n288), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT67), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n273), .A2(KEYINPUT67), .A3(G232), .A4(new_n288), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n273), .A2(G238), .A3(G1698), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n267), .A2(new_n280), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(G107), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n383), .A2(new_n384), .A3(new_n385), .A4(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n380), .B1(new_n388), .B2(new_n294), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n389), .A2(new_n354), .ZN(new_n390));
  OAI21_X1  g0190(.A(KEYINPUT69), .B1(new_n373), .B2(new_n390), .ZN(new_n391));
  OR2_X1    g0191(.A1(new_n389), .A2(new_n354), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT69), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n392), .A2(new_n393), .A3(new_n371), .A4(new_n372), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n389), .A2(G190), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n391), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n366), .A2(new_n247), .ZN(new_n397));
  INV_X1    g0197(.A(new_n358), .ZN(new_n398));
  AND4_X1   g0198(.A1(KEYINPUT68), .A2(new_n397), .A3(new_n398), .A4(new_n369), .ZN(new_n399));
  OAI22_X1  g0199(.A1(new_n399), .A2(new_n370), .B1(new_n389), .B2(G169), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT70), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  OAI221_X1 g0202(.A(KEYINPUT70), .B1(new_n389), .B2(G169), .C1(new_n399), .C2(new_n370), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n389), .A2(new_n313), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n402), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n396), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n363), .A2(new_n364), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n408), .A2(new_n245), .ZN(new_n409));
  INV_X1    g0209(.A(new_n368), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n409), .B1(new_n410), .B2(new_n408), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n362), .A2(new_n325), .ZN(new_n412));
  OAI21_X1  g0212(.A(G20), .B1(new_n412), .B2(new_n201), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n254), .A2(G159), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n386), .A2(KEYINPUT7), .A3(new_n219), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n274), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n415), .B1(new_n417), .B2(G68), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n277), .B1(new_n418), .B2(KEYINPUT16), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT16), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n325), .B1(new_n271), .B2(new_n274), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n420), .B1(new_n421), .B2(new_n415), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n411), .B1(new_n419), .B2(new_n422), .ZN(new_n423));
  OR2_X1    g0223(.A1(G223), .A2(G1698), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n213), .A2(G1698), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n267), .A2(new_n424), .A3(new_n280), .A4(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(G33), .A2(G87), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n293), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(G232), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n378), .A2(new_n429), .ZN(new_n430));
  NOR3_X1   g0230(.A1(new_n428), .A2(new_n430), .A3(new_n376), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(G190), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n426), .A2(new_n427), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(new_n294), .ZN(new_n434));
  INV_X1    g0234(.A(new_n430), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n434), .A2(new_n377), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(G200), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n423), .A2(new_n432), .A3(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT17), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n423), .A2(KEYINPUT17), .A3(new_n432), .A4(new_n437), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n411), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n417), .A2(G68), .ZN(new_n444));
  INV_X1    g0244(.A(new_n415), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n444), .A2(KEYINPUT16), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(new_n247), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n275), .A2(G68), .ZN(new_n448));
  AOI21_X1  g0248(.A(KEYINPUT16), .B1(new_n448), .B2(new_n445), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n443), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n436), .A2(G169), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n431), .A2(G179), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(KEYINPUT18), .B1(new_n450), .B2(new_n453), .ZN(new_n454));
  AND2_X1   g0254(.A1(new_n451), .A2(new_n452), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT18), .ZN(new_n456));
  NOR3_X1   g0256(.A1(new_n423), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT75), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n454), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n450), .A2(KEYINPUT18), .A3(new_n453), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(KEYINPUT75), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n442), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT76), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n457), .A2(new_n458), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n456), .B1(new_n423), .B2(new_n455), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n465), .A2(new_n461), .A3(new_n466), .ZN(new_n467));
  AND2_X1   g0267(.A1(new_n440), .A2(new_n441), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(KEYINPUT76), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n406), .B1(new_n464), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n203), .A2(G20), .ZN(new_n472));
  INV_X1    g0272(.A(G150), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n219), .A2(G33), .ZN(new_n474));
  OAI221_X1 g0274(.A(new_n472), .B1(new_n473), .B2(new_n255), .C1(new_n474), .C2(new_n407), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(new_n247), .ZN(new_n476));
  OAI21_X1  g0276(.A(G50), .B1(new_n219), .B2(G1), .ZN(new_n477));
  XNOR2_X1  g0277(.A(new_n477), .B(KEYINPUT66), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(new_n248), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n476), .B(new_n479), .C1(G50), .C2(new_n242), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT9), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n378), .A2(new_n213), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n273), .A2(G222), .A3(new_n288), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(KEYINPUT65), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n273), .A2(G223), .A3(G1698), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n386), .A2(G77), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT65), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n273), .A2(new_n488), .A3(G222), .A4(new_n288), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n485), .A2(new_n486), .A3(new_n487), .A4(new_n489), .ZN(new_n490));
  AOI211_X1 g0290(.A(new_n376), .B(new_n483), .C1(new_n490), .C2(new_n294), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n482), .B1(new_n491), .B2(G190), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n480), .A2(new_n481), .ZN(new_n493));
  OR2_X1    g0293(.A1(new_n491), .A2(new_n354), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n492), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(KEYINPUT10), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT10), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n492), .A2(new_n497), .A3(new_n493), .A4(new_n494), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n491), .A2(new_n313), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n480), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n491), .A2(G169), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n499), .A2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT13), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n213), .A2(new_n288), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n429), .A2(G1698), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n267), .A2(new_n507), .A3(new_n280), .A4(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(new_n321), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n376), .B1(new_n510), .B2(new_n294), .ZN(new_n511));
  AND3_X1   g0311(.A1(new_n293), .A2(G238), .A3(new_n374), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n506), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n293), .B1(new_n509), .B2(new_n321), .ZN(new_n515));
  NOR4_X1   g0315(.A1(new_n515), .A2(KEYINPUT13), .A3(new_n512), .A4(new_n376), .ZN(new_n516));
  OAI21_X1  g0316(.A(G169), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(KEYINPUT14), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n514), .A2(new_n516), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(G179), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT14), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n521), .B(G169), .C1(new_n514), .C2(new_n516), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n518), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(KEYINPUT73), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT71), .ZN(new_n525));
  AOI211_X1 g0325(.A(G68), .B(new_n242), .C1(new_n525), .C2(KEYINPUT12), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n526), .B1(new_n525), .B2(KEYINPUT12), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT12), .ZN(new_n528));
  OAI211_X1 g0328(.A(KEYINPUT71), .B(new_n528), .C1(new_n242), .C2(G68), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n527), .B(new_n529), .C1(new_n325), .C2(new_n410), .ZN(new_n530));
  XOR2_X1   g0330(.A(new_n530), .B(KEYINPUT72), .Z(new_n531));
  NAND2_X1  g0331(.A1(new_n325), .A2(G20), .ZN(new_n532));
  OAI221_X1 g0332(.A(new_n532), .B1(new_n474), .B2(new_n256), .C1(new_n255), .C2(new_n202), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n247), .ZN(new_n534));
  XNOR2_X1  g0334(.A(new_n534), .B(KEYINPUT11), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n531), .A2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT73), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n518), .A2(new_n520), .A3(new_n537), .A4(new_n522), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n524), .A2(new_n536), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n519), .A2(G190), .ZN(new_n540));
  OAI21_X1  g0340(.A(G200), .B1(new_n514), .B2(new_n516), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n531), .A2(new_n535), .A3(new_n540), .A4(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n505), .A2(new_n543), .ZN(new_n544));
  AND2_X1   g0344(.A1(new_n471), .A2(new_n544), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n248), .B(G116), .C1(G1), .C2(new_n249), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n245), .A2(new_n208), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n246), .A2(new_n220), .B1(G20), .B2(new_n208), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n284), .B(new_n219), .C1(G33), .C2(new_n251), .ZN(new_n549));
  AOI21_X1  g0349(.A(KEYINPUT20), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  AND3_X1   g0350(.A1(new_n548), .A2(KEYINPUT20), .A3(new_n549), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n546), .B(new_n547), .C1(new_n550), .C2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n288), .A2(G257), .ZN(new_n554));
  NAND2_X1  g0354(.A1(G264), .A2(G1698), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n267), .A2(new_n280), .A3(new_n554), .A4(new_n555), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n556), .B(new_n294), .C1(G303), .C2(new_n273), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n304), .A2(G270), .A3(new_n293), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n557), .A2(new_n558), .A3(new_n306), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(G200), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n553), .B(new_n560), .C1(new_n310), .C2(new_n559), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT21), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n559), .A2(G169), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n562), .B1(new_n553), .B2(new_n563), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n552), .A2(KEYINPUT21), .A3(G169), .A4(new_n559), .ZN(new_n565));
  AND4_X1   g0365(.A1(G179), .A2(new_n557), .A3(new_n558), .A4(new_n306), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n552), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n561), .A2(new_n564), .A3(new_n565), .A4(new_n567), .ZN(new_n568));
  OR2_X1    g0368(.A1(new_n568), .A2(KEYINPUT80), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(KEYINPUT80), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n222), .A2(new_n259), .A3(G13), .A4(G20), .ZN(new_n572));
  XNOR2_X1  g0372(.A(new_n572), .B(KEYINPUT25), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n574), .B1(new_n250), .B2(new_n259), .ZN(new_n575));
  INV_X1    g0375(.A(new_n575), .ZN(new_n576));
  AND3_X1   g0376(.A1(new_n304), .A2(G264), .A3(new_n293), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n267), .A2(new_n280), .A3(G250), .A4(new_n288), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT84), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n273), .A2(KEYINPUT84), .A3(G250), .A4(new_n288), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n273), .A2(G257), .A3(G1698), .ZN(new_n582));
  NAND2_X1  g0382(.A1(G33), .A2(G294), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n580), .A2(new_n581), .A3(new_n582), .A4(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n577), .B1(new_n584), .B2(new_n294), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n306), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n354), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n585), .A2(new_n310), .A3(new_n306), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT23), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n590), .B1(new_n219), .B2(G107), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n259), .A2(KEYINPUT23), .A3(G20), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n342), .A2(new_n219), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT81), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT82), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT22), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  OAI21_X1  g0400(.A(KEYINPUT82), .B1(KEYINPUT81), .B2(KEYINPUT22), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g0402(.A(G87), .B1(new_n597), .B2(new_n599), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n602), .B1(new_n326), .B2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  NOR3_X1   g0405(.A1(new_n602), .A2(new_n326), .A3(new_n603), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n596), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(KEYINPUT24), .ZN(new_n608));
  INV_X1    g0408(.A(new_n601), .ZN(new_n609));
  NOR3_X1   g0409(.A1(KEYINPUT81), .A2(KEYINPUT82), .A3(KEYINPUT22), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AND3_X1   g0411(.A1(new_n267), .A2(new_n280), .A3(new_n219), .ZN(new_n612));
  INV_X1    g0412(.A(new_n603), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(new_n604), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT24), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n615), .A2(new_n616), .A3(new_n596), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n608), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(KEYINPUT83), .B1(new_n618), .B2(new_n247), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n616), .B1(new_n615), .B2(new_n596), .ZN(new_n620));
  AOI211_X1 g0420(.A(KEYINPUT24), .B(new_n595), .C1(new_n614), .C2(new_n604), .ZN(new_n621));
  OAI211_X1 g0421(.A(KEYINPUT83), .B(new_n247), .C1(new_n620), .C2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(new_n622), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n576), .B(new_n589), .C1(new_n619), .C2(new_n623), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n331), .B(new_n336), .C1(new_n250), .C2(new_n335), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n351), .A2(new_n315), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n353), .A2(new_n313), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n247), .B1(new_n620), .B2(new_n621), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT83), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n575), .B1(new_n631), .B2(new_n622), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n586), .A2(new_n315), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n633), .B1(G179), .B2(new_n586), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n624), .B(new_n628), .C1(new_n632), .C2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  AND4_X1   g0436(.A1(new_n357), .A2(new_n545), .A3(new_n571), .A4(new_n636), .ZN(G372));
  INV_X1    g0437(.A(new_n628), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n356), .A2(new_n278), .A3(new_n316), .A4(new_n314), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n638), .B1(new_n639), .B2(KEYINPUT26), .ZN(new_n640));
  INV_X1    g0440(.A(new_n317), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n564), .A2(new_n565), .A3(new_n567), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n643), .B1(new_n632), .B2(new_n634), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n641), .B1(new_n644), .B2(new_n624), .ZN(new_n645));
  NOR3_X1   g0445(.A1(new_n337), .A2(new_n352), .A3(new_n355), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n278), .B1(G190), .B2(new_n312), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n646), .B1(new_n647), .B2(new_n309), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT26), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n640), .B1(new_n645), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n545), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT85), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n653), .B1(new_n454), .B2(new_n457), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n460), .A2(new_n466), .A3(KEYINPUT85), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AND3_X1   g0456(.A1(new_n402), .A2(new_n403), .A3(new_n404), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n542), .A2(new_n657), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n658), .A2(new_n539), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n656), .B1(new_n659), .B2(new_n442), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n503), .B1(new_n660), .B2(new_n499), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n652), .A2(new_n661), .ZN(G369));
  INV_X1    g0462(.A(G13), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n663), .A2(G20), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(new_n222), .ZN(new_n665));
  OR2_X1    g0465(.A1(new_n665), .A2(KEYINPUT27), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(KEYINPUT27), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n666), .A2(G213), .A3(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(G343), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n552), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g0471(.A(new_n671), .B(KEYINPUT86), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n672), .B1(new_n569), .B2(new_n570), .ZN(new_n673));
  INV_X1    g0473(.A(new_n672), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n674), .A2(new_n643), .ZN(new_n675));
  OAI21_X1  g0475(.A(G330), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n632), .A2(new_n634), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(new_n670), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n624), .B1(new_n632), .B2(new_n634), .ZN(new_n680));
  INV_X1    g0480(.A(new_n670), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n632), .A2(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n679), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n677), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n644), .A2(new_n624), .A3(new_n681), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(G399));
  INV_X1    g0486(.A(new_n223), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n687), .A2(G41), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n320), .A2(G116), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n689), .A2(G1), .A3(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n691), .B1(new_n218), .B2(new_n689), .ZN(new_n692));
  XNOR2_X1  g0492(.A(new_n692), .B(KEYINPUT28), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n644), .A2(new_n648), .A3(new_n317), .A4(new_n624), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n641), .A2(new_n649), .A3(new_n356), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(new_n640), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(new_n681), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(KEYINPUT29), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT29), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n651), .A2(new_n699), .A3(new_n681), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(G330), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n559), .A2(new_n313), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n308), .A2(new_n351), .A3(new_n586), .A4(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT30), .ZN(new_n705));
  AND3_X1   g0505(.A1(new_n353), .A2(new_n585), .A3(new_n566), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n705), .B1(new_n312), .B2(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n353), .A2(new_n585), .A3(new_n566), .ZN(new_n708));
  NOR3_X1   g0508(.A1(new_n308), .A2(new_n708), .A3(KEYINPUT30), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n704), .B1(new_n707), .B2(new_n709), .ZN(new_n710));
  AND3_X1   g0510(.A1(new_n710), .A2(KEYINPUT31), .A3(new_n670), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(KEYINPUT87), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT87), .ZN(new_n713));
  OAI211_X1 g0513(.A(new_n713), .B(new_n704), .C1(new_n707), .C2(new_n709), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n712), .A2(new_n670), .A3(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT31), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n711), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n636), .A2(new_n357), .A3(new_n571), .A4(new_n681), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n702), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n701), .A2(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n693), .B1(new_n720), .B2(G1), .ZN(G364));
  NAND2_X1  g0521(.A1(new_n664), .A2(G45), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n689), .A2(G1), .A3(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n677), .A2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n673), .ZN(new_n726));
  INV_X1    g0526(.A(new_n675), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n725), .B1(G330), .B2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n219), .A2(G190), .ZN(new_n730));
  NOR2_X1   g0530(.A1(G179), .A2(G200), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(G159), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n219), .B1(new_n731), .B2(G190), .ZN(new_n735));
  OAI22_X1  g0535(.A1(new_n734), .A2(KEYINPUT32), .B1(new_n251), .B2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n354), .A2(G179), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(new_n730), .ZN(new_n738));
  XNOR2_X1  g0538(.A(new_n738), .B(KEYINPUT89), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(new_n259), .ZN(new_n740));
  AOI211_X1 g0540(.A(new_n736), .B(new_n740), .C1(KEYINPUT32), .C2(new_n734), .ZN(new_n741));
  NAND2_X1  g0541(.A1(G20), .A2(G179), .ZN(new_n742));
  XNOR2_X1  g0542(.A(new_n742), .B(KEYINPUT88), .ZN(new_n743));
  AND3_X1   g0543(.A1(new_n743), .A2(new_n310), .A3(G200), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n743), .A2(new_n310), .A3(new_n354), .ZN(new_n746));
  OAI22_X1  g0546(.A1(new_n745), .A2(new_n325), .B1(new_n256), .B2(new_n746), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n743), .A2(G190), .A3(G200), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n747), .B1(G50), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n743), .A2(G190), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(G200), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(G58), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n737), .A2(G20), .A3(G190), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n386), .B1(new_n755), .B2(G87), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n741), .A2(new_n750), .A3(new_n753), .A4(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n735), .ZN(new_n758));
  AOI22_X1  g0558(.A1(new_n749), .A2(G326), .B1(G294), .B2(new_n758), .ZN(new_n759));
  XOR2_X1   g0559(.A(new_n759), .B(KEYINPUT90), .Z(new_n760));
  AOI21_X1  g0560(.A(new_n273), .B1(new_n733), .B2(G329), .ZN(new_n761));
  INV_X1    g0561(.A(G311), .ZN(new_n762));
  INV_X1    g0562(.A(G283), .ZN(new_n763));
  OAI221_X1 g0563(.A(new_n761), .B1(new_n746), .B2(new_n762), .C1(new_n739), .C2(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n764), .B1(G303), .B2(new_n755), .ZN(new_n765));
  XOR2_X1   g0565(.A(KEYINPUT33), .B(G317), .Z(new_n766));
  OAI211_X1 g0566(.A(new_n760), .B(new_n765), .C1(new_n745), .C2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n752), .ZN(new_n768));
  INV_X1    g0568(.A(G322), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n757), .B1(new_n767), .B2(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n220), .B1(G20), .B2(new_n315), .ZN(new_n772));
  NOR2_X1   g0572(.A1(G13), .A2(G33), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(G20), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n772), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n687), .A2(new_n273), .ZN(new_n777));
  OR2_X1    g0577(.A1(new_n218), .A2(G45), .ZN(new_n778));
  OAI211_X1 g0578(.A(new_n777), .B(new_n778), .C1(new_n237), .C2(new_n302), .ZN(new_n779));
  INV_X1    g0579(.A(G355), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n273), .A2(new_n223), .ZN(new_n781));
  OAI221_X1 g0581(.A(new_n779), .B1(G116), .B2(new_n223), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  AOI22_X1  g0582(.A1(new_n771), .A2(new_n772), .B1(new_n776), .B2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n775), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n783), .B1(new_n728), .B2(new_n784), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n729), .B1(new_n723), .B2(new_n785), .ZN(G396));
  INV_X1    g0586(.A(KEYINPUT92), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n681), .B1(new_n371), .B2(new_n372), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n657), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n788), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n396), .A2(new_n405), .A3(new_n790), .ZN(new_n791));
  NAND4_X1  g0591(.A1(new_n402), .A2(new_n403), .A3(new_n404), .A4(new_n788), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(KEYINPUT92), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n789), .A2(new_n791), .A3(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(KEYINPUT93), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND4_X1  g0596(.A1(new_n789), .A2(new_n791), .A3(new_n793), .A4(KEYINPUT93), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n576), .B1(new_n619), .B2(new_n623), .ZN(new_n800));
  INV_X1    g0600(.A(new_n634), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n642), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n624), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n317), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n650), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n670), .B1(new_n806), .B2(new_n640), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n799), .B(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n719), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(new_n723), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n752), .A2(G143), .B1(new_n744), .B2(G150), .ZN(new_n812));
  INV_X1    g0612(.A(G137), .ZN(new_n813));
  INV_X1    g0613(.A(G159), .ZN(new_n814));
  OAI221_X1 g0614(.A(new_n812), .B1(new_n813), .B2(new_n748), .C1(new_n814), .C2(new_n746), .ZN(new_n815));
  INV_X1    g0615(.A(KEYINPUT34), .ZN(new_n816));
  OR2_X1    g0616(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n755), .A2(G50), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n815), .A2(new_n816), .ZN(new_n819));
  INV_X1    g0619(.A(G132), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n273), .B1(new_n735), .B2(new_n362), .C1(new_n820), .C2(new_n732), .ZN(new_n821));
  INV_X1    g0621(.A(new_n739), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n821), .B1(new_n822), .B2(G68), .ZN(new_n823));
  NAND4_X1  g0623(.A1(new_n817), .A2(new_n818), .A3(new_n819), .A4(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n822), .A2(G87), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n825), .B1(new_n762), .B2(new_n732), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT91), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n273), .B(new_n828), .C1(G107), .C2(new_n755), .ZN(new_n829));
  AOI22_X1  g0629(.A1(G294), .A2(new_n752), .B1(new_n749), .B2(G303), .ZN(new_n830));
  OAI22_X1  g0630(.A1(new_n745), .A2(new_n763), .B1(new_n251), .B2(new_n735), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n831), .B1(new_n826), .B2(new_n827), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n829), .A2(new_n830), .A3(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n746), .A2(new_n208), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n824), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n772), .A2(new_n773), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n835), .A2(new_n772), .B1(new_n256), .B2(new_n836), .ZN(new_n837));
  OAI211_X1 g0637(.A(new_n837), .B(new_n724), .C1(new_n774), .C2(new_n798), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n811), .A2(new_n838), .ZN(G384));
  NAND2_X1  g0639(.A1(new_n536), .A2(new_n670), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n543), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n539), .A2(new_n542), .A3(new_n840), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n792), .B(new_n787), .ZN(new_n846));
  AOI21_X1  g0646(.A(KEYINPUT93), .B1(new_n846), .B2(new_n791), .ZN(new_n847));
  INV_X1    g0647(.A(new_n797), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n651), .B(new_n681), .C1(new_n847), .C2(new_n848), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n405), .A2(new_n670), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n845), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT38), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n325), .B1(new_n274), .B2(new_n416), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n420), .B1(new_n854), .B2(new_n415), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n411), .B1(new_n419), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(KEYINPUT94), .B1(new_n856), .B2(new_n668), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n446), .A2(new_n855), .A3(new_n247), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(new_n443), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT94), .ZN(new_n860));
  INV_X1    g0660(.A(new_n668), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  AND2_X1   g0662(.A1(new_n857), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n863), .B1(new_n467), .B2(new_n468), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n450), .B1(new_n453), .B2(new_n861), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT37), .ZN(new_n866));
  AND3_X1   g0666(.A1(new_n865), .A2(new_n866), .A3(new_n438), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n859), .A2(new_n453), .ZN(new_n868));
  NAND4_X1  g0668(.A1(new_n857), .A2(new_n862), .A3(new_n438), .A4(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n867), .B1(KEYINPUT37), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n853), .B1(new_n864), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n869), .A2(KEYINPUT37), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n865), .A2(new_n866), .A3(new_n438), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  OAI211_X1 g0674(.A(KEYINPUT38), .B(new_n874), .C1(new_n462), .C2(new_n863), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n871), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n852), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT39), .ZN(new_n878));
  INV_X1    g0678(.A(new_n655), .ZN(new_n879));
  AOI21_X1  g0679(.A(KEYINPUT85), .B1(new_n460), .B2(new_n466), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n468), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n423), .A2(new_n668), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n865), .A2(new_n438), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(KEYINPUT37), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n873), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT38), .B1(new_n883), .B2(new_n886), .ZN(new_n887));
  NOR3_X1   g0687(.A1(new_n864), .A2(new_n870), .A3(new_n853), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n878), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n539), .A2(new_n670), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n871), .A2(new_n875), .A3(KEYINPUT39), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n654), .A2(new_n655), .A3(new_n668), .ZN(new_n893));
  AND3_X1   g0693(.A1(new_n877), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n701), .A2(new_n545), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(new_n661), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n894), .B(new_n896), .ZN(new_n897));
  AOI22_X1  g0697(.A1(new_n796), .A2(new_n797), .B1(new_n842), .B2(new_n843), .ZN(new_n898));
  NOR2_X1   g0698(.A1(KEYINPUT95), .A2(KEYINPUT31), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n715), .A2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n899), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n712), .A2(new_n670), .A3(new_n714), .A4(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n718), .A2(new_n900), .A3(new_n902), .ZN(new_n903));
  AND2_X1   g0703(.A1(new_n898), .A2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT40), .ZN(new_n905));
  INV_X1    g0705(.A(new_n882), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n906), .B1(new_n656), .B2(new_n468), .ZN(new_n907));
  INV_X1    g0707(.A(new_n886), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n853), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n905), .B1(new_n909), .B2(new_n875), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n876), .A2(new_n898), .A3(new_n903), .ZN(new_n911));
  AOI22_X1  g0711(.A1(new_n904), .A2(new_n910), .B1(new_n911), .B2(new_n905), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n545), .A2(new_n903), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n912), .B(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(G330), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n897), .B(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(new_n222), .B2(new_n664), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n262), .A2(new_n263), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT35), .ZN(new_n919));
  AOI211_X1 g0719(.A(new_n219), .B(new_n220), .C1(new_n918), .C2(new_n919), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n920), .B(G116), .C1(new_n919), .C2(new_n918), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n921), .B(KEYINPUT36), .ZN(new_n922));
  OAI21_X1  g0722(.A(G77), .B1(new_n362), .B2(new_n325), .ZN(new_n923));
  OAI22_X1  g0723(.A1(new_n923), .A2(new_n218), .B1(G50), .B2(new_n325), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n924), .A2(G1), .A3(new_n663), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n917), .A2(new_n922), .A3(new_n925), .ZN(new_n926));
  XOR2_X1   g0726(.A(new_n926), .B(KEYINPUT96), .Z(G367));
  INV_X1    g0727(.A(KEYINPUT104), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n722), .A2(G1), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n720), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT101), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT100), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n677), .A2(new_n933), .A3(new_n683), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n278), .A2(new_n670), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n311), .A2(new_n317), .A3(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT97), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND4_X1  g0739(.A1(new_n311), .A2(new_n317), .A3(KEYINPUT97), .A4(new_n936), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n641), .A2(new_n670), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n942), .A2(KEYINPUT45), .A3(new_n685), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(KEYINPUT45), .B1(new_n942), .B2(new_n685), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n939), .A2(new_n940), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n685), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT99), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(KEYINPUT44), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n950), .A2(KEYINPUT44), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n948), .A2(new_n949), .A3(new_n951), .A4(new_n952), .ZN(new_n953));
  OAI211_X1 g0753(.A(new_n950), .B(KEYINPUT44), .C1(new_n947), .C2(new_n685), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n935), .B1(new_n946), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n942), .A2(new_n685), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT45), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(new_n943), .ZN(new_n960));
  NAND4_X1  g0760(.A1(new_n960), .A2(new_n934), .A3(new_n954), .A4(new_n953), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n956), .A2(new_n961), .ZN(new_n962));
  OAI221_X1 g0762(.A(new_n679), .B1(new_n643), .B2(new_n670), .C1(new_n680), .C2(new_n682), .ZN(new_n963));
  INV_X1    g0763(.A(new_n680), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n643), .A2(new_n670), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  AND3_X1   g0766(.A1(new_n963), .A2(new_n676), .A3(new_n966), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n676), .B1(new_n963), .B2(new_n966), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND4_X1  g0769(.A1(new_n969), .A2(new_n698), .A3(new_n700), .A4(new_n809), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n932), .B1(new_n962), .B2(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n967), .A2(new_n968), .ZN(new_n972));
  NOR3_X1   g0772(.A1(new_n972), .A2(new_n701), .A3(new_n719), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n973), .A2(KEYINPUT101), .A3(new_n961), .A4(new_n956), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n931), .B1(new_n971), .B2(new_n974), .ZN(new_n975));
  XNOR2_X1  g0775(.A(KEYINPUT98), .B(KEYINPUT41), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n688), .B(new_n976), .Z(new_n977));
  OAI21_X1  g0777(.A(new_n930), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n942), .A2(new_n964), .A3(new_n965), .ZN(new_n979));
  OR2_X1    g0779(.A1(new_n979), .A2(KEYINPUT42), .ZN(new_n980));
  AND2_X1   g0780(.A1(new_n947), .A2(new_n678), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n681), .B1(new_n981), .B2(new_n641), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n979), .A2(KEYINPUT42), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n980), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  AND2_X1   g0784(.A1(new_n337), .A2(new_n670), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n628), .B1(new_n646), .B2(new_n985), .ZN(new_n986));
  OR2_X1    g0786(.A1(new_n985), .A2(new_n628), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(KEYINPUT43), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n984), .A2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n684), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(new_n942), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n991), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n984), .A2(new_n993), .A3(new_n990), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n989), .A2(KEYINPUT43), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n997), .B(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n978), .A2(new_n999), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n745), .A2(new_n814), .B1(new_n202), .B2(new_n746), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n735), .A2(new_n325), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n273), .B1(new_n754), .B2(new_n362), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n738), .ZN(new_n1004));
  AOI211_X1 g0804(.A(new_n1002), .B(new_n1003), .C1(G77), .C2(new_n1004), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n1005), .B1(new_n813), .B2(new_n732), .C1(new_n473), .C2(new_n768), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n1001), .B(new_n1006), .C1(G143), .C2(new_n749), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT103), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n386), .B1(new_n735), .B2(new_n259), .C1(new_n251), .C2(new_n738), .ZN(new_n1009));
  INV_X1    g0809(.A(G294), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n745), .A2(new_n1010), .B1(new_n763), .B2(new_n746), .ZN(new_n1011));
  OAI21_X1  g0811(.A(KEYINPUT46), .B1(new_n754), .B2(new_n208), .ZN(new_n1012));
  OR3_X1    g0812(.A1(new_n754), .A2(KEYINPUT46), .A3(new_n208), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n1009), .B(new_n1011), .C1(new_n1012), .C2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(G303), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n768), .A2(new_n1015), .B1(new_n762), .B2(new_n748), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT102), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  AND2_X1   g0818(.A1(new_n1014), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(G317), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1019), .B1(new_n1017), .B2(new_n1016), .C1(new_n1020), .C2(new_n732), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1008), .A2(new_n1021), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT47), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1023), .A2(new_n772), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n777), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n776), .B1(new_n223), .B2(new_n335), .C1(new_n233), .C2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n988), .A2(new_n775), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n1024), .A2(new_n724), .A3(new_n1026), .A4(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n928), .B1(new_n1000), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1028), .ZN(new_n1030));
  AOI211_X1 g0830(.A(KEYINPUT104), .B(new_n1030), .C1(new_n978), .C2(new_n999), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n1032), .ZN(G387));
  NAND2_X1  g0833(.A1(new_n931), .A2(new_n972), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1034), .A2(new_n688), .A3(new_n970), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n768), .A2(new_n202), .B1(new_n325), .B2(new_n746), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(new_n408), .B2(new_n744), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n273), .B1(new_n754), .B2(new_n256), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n335), .A2(new_n735), .B1(new_n732), .B2(new_n473), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n1038), .B(new_n1039), .C1(new_n822), .C2(G97), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1037), .B(new_n1040), .C1(new_n814), .C2(new_n748), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n752), .A2(G317), .B1(new_n744), .B2(G311), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n1042), .B1(new_n1015), .B2(new_n746), .C1(new_n769), .C2(new_n748), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT48), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1044), .B1(new_n763), .B2(new_n735), .C1(new_n1010), .C2(new_n754), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT49), .ZN(new_n1046));
  OR2_X1    g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n273), .B1(new_n733), .B2(G326), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1047), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n738), .A2(new_n208), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1041), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT105), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n230), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1053), .B1(new_n1054), .B2(new_n302), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n408), .A2(new_n202), .ZN(new_n1056));
  AOI211_X1 g0856(.A(G116), .B(new_n320), .C1(new_n1056), .C2(KEYINPUT50), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(G68), .A2(G77), .ZN(new_n1058));
  OR2_X1    g0858(.A1(new_n1056), .A2(KEYINPUT50), .ZN(new_n1059));
  NAND4_X1  g0859(.A1(new_n1057), .A2(new_n302), .A3(new_n1058), .A4(new_n1059), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n230), .A2(KEYINPUT105), .A3(G45), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n1055), .A2(new_n777), .A3(new_n1060), .A4(new_n1061), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1062), .B1(G107), .B2(new_n223), .C1(new_n690), .C2(new_n781), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n1052), .A2(new_n772), .B1(new_n776), .B2(new_n1063), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n1064), .B(new_n724), .C1(new_n683), .C2(new_n784), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1035), .B(new_n1065), .C1(new_n930), .C2(new_n972), .ZN(G393));
  INV_X1    g0866(.A(KEYINPUT109), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n992), .B1(new_n946), .B2(new_n955), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n960), .A2(new_n684), .A3(new_n954), .A4(new_n953), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n1068), .A2(new_n1069), .B1(new_n720), .B2(new_n969), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n689), .B(new_n1070), .C1(new_n971), .C2(new_n974), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1068), .A2(new_n929), .A3(new_n1069), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n768), .A2(new_n814), .B1(new_n473), .B2(new_n748), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT51), .ZN(new_n1074));
  OR2_X1    g0874(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n735), .A2(new_n256), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n273), .B1(new_n754), .B2(new_n325), .ZN(new_n1077));
  AOI211_X1 g0877(.A(new_n1076), .B(new_n1077), .C1(G143), .C2(new_n733), .ZN(new_n1078));
  AND3_X1   g0878(.A1(new_n1075), .A2(new_n825), .A3(new_n1078), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n745), .A2(new_n202), .B1(new_n407), .B2(new_n746), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n1073), .A2(new_n1074), .B1(new_n1080), .B2(KEYINPUT106), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1079), .B(new_n1081), .C1(KEYINPUT106), .C2(new_n1080), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT107), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n735), .A2(new_n208), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n386), .B1(new_n732), .B2(new_n769), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n1085), .B(new_n740), .C1(G283), .C2(new_n755), .ZN(new_n1086));
  XOR2_X1   g0886(.A(new_n1086), .B(KEYINPUT108), .Z(new_n1087));
  OAI22_X1  g0887(.A1(new_n768), .A2(new_n762), .B1(new_n1020), .B2(new_n748), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1088), .B(KEYINPUT52), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n746), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(G294), .A2(new_n1090), .B1(new_n744), .B2(G303), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1087), .A2(new_n1089), .A3(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1083), .B1(new_n1084), .B2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n723), .B1(new_n1093), .B2(new_n772), .ZN(new_n1094));
  OAI221_X1 g0894(.A(new_n776), .B1(new_n251), .B2(new_n223), .C1(new_n240), .C2(new_n1025), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n1094), .B(new_n1095), .C1(new_n784), .C2(new_n942), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1072), .A2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1067), .B1(new_n1071), .B2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1070), .B1(new_n971), .B2(new_n974), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n688), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1097), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1100), .A2(KEYINPUT109), .A3(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1098), .A2(new_n1102), .ZN(G390));
  AOI21_X1  g0903(.A(KEYINPUT39), .B1(new_n909), .B2(new_n875), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n891), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n852), .A2(new_n890), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n890), .B1(new_n909), .B2(new_n875), .ZN(new_n1107));
  AND2_X1   g0907(.A1(new_n696), .A2(new_n681), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n850), .B1(new_n1108), .B2(new_n798), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1107), .B1(new_n1109), .B2(new_n845), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n717), .A2(new_n718), .ZN(new_n1111));
  AND3_X1   g0911(.A1(new_n898), .A2(new_n1111), .A3(G330), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1106), .A2(new_n1110), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n890), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n850), .B1(new_n807), .B2(new_n798), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1114), .B1(new_n1115), .B2(new_n845), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n889), .A2(new_n891), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n851), .B1(new_n799), .B2(new_n697), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(new_n844), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n1116), .A2(new_n1117), .B1(new_n1119), .B2(new_n1107), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n702), .B1(new_n796), .B2(new_n797), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n903), .A2(new_n1121), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1122), .A2(new_n845), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1113), .B1(new_n1120), .B2(new_n1123), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n903), .A2(new_n471), .A3(G330), .A4(new_n544), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n895), .A2(new_n661), .A3(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n844), .B1(new_n903), .B2(new_n1121), .ZN(new_n1127));
  OAI21_X1  g0927(.A(KEYINPUT110), .B1(new_n1112), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1122), .A2(new_n845), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT110), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1118), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1128), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1115), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n844), .B1(new_n719), .B2(new_n798), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1133), .B1(new_n1123), .B2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1126), .B1(new_n1132), .B2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n689), .B1(new_n1124), .B2(new_n1136), .ZN(new_n1137));
  AND3_X1   g0937(.A1(new_n1106), .A2(new_n1110), .A3(new_n1112), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1123), .B1(new_n1106), .B2(new_n1110), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n719), .A2(new_n898), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1130), .B1(new_n1129), .B2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1109), .B1(new_n1127), .B2(KEYINPUT110), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1135), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1126), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1140), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1137), .A2(new_n1147), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n754), .A2(new_n473), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n1149), .B(KEYINPUT112), .ZN(new_n1150));
  XOR2_X1   g0950(.A(new_n1150), .B(KEYINPUT53), .Z(new_n1151));
  OAI21_X1  g0951(.A(new_n1151), .B1(new_n813), .B2(new_n745), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n738), .A2(new_n202), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(KEYINPUT54), .B(G143), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1154), .B(KEYINPUT111), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  OAI22_X1  g0956(.A1(new_n768), .A2(new_n820), .B1(new_n746), .B2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n386), .B1(new_n733), .B2(G125), .ZN(new_n1158));
  INV_X1    g0958(.A(G128), .ZN(new_n1159));
  OAI221_X1 g0959(.A(new_n1158), .B1(new_n814), .B2(new_n735), .C1(new_n748), .C2(new_n1159), .ZN(new_n1160));
  NOR4_X1   g0960(.A1(new_n1152), .A2(new_n1153), .A3(new_n1157), .A4(new_n1160), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(G116), .A2(new_n752), .B1(new_n749), .B2(G283), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1162), .B1(new_n251), .B2(new_n746), .ZN(new_n1163));
  AOI211_X1 g0963(.A(new_n273), .B(new_n1076), .C1(G294), .C2(new_n733), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n1164), .B1(new_n325), .B2(new_n739), .C1(new_n319), .C2(new_n754), .ZN(new_n1165));
  AOI211_X1 g0965(.A(new_n1163), .B(new_n1165), .C1(G107), .C2(new_n744), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n772), .B1(new_n1161), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n836), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1167), .B1(new_n408), .B2(new_n1168), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n723), .B(new_n1169), .C1(new_n1117), .C2(new_n773), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1170), .B1(new_n1124), .B2(new_n929), .ZN(new_n1171));
  AND2_X1   g0971(.A1(new_n1148), .A2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(G378));
  INV_X1    g0973(.A(new_n894), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n505), .A2(KEYINPUT55), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT55), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(new_n499), .B2(new_n504), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n480), .A2(new_n861), .ZN(new_n1178));
  XOR2_X1   g0978(.A(new_n1178), .B(KEYINPUT56), .Z(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  OR3_X1    g0980(.A1(new_n1175), .A2(new_n1177), .A3(new_n1180), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1180), .B1(new_n1175), .B2(new_n1177), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(new_n912), .B2(G330), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n911), .A2(new_n905), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n909), .A2(new_n875), .ZN(new_n1186));
  NAND4_X1  g0986(.A1(new_n1186), .A2(KEYINPUT40), .A3(new_n903), .A4(new_n898), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1185), .A2(new_n1183), .A3(G330), .A4(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1174), .B1(new_n1184), .B2(new_n1189), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1185), .A2(G330), .A3(new_n1187), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1183), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1193), .A2(new_n894), .A3(new_n1188), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1190), .A2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(new_n929), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n1004), .A2(G58), .B1(new_n733), .B2(G283), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1197), .B1(new_n256), .B2(new_n754), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1002), .B1(new_n749), .B2(G116), .ZN(new_n1199));
  XOR2_X1   g0999(.A(new_n1199), .B(KEYINPUT115), .Z(new_n1200));
  AOI211_X1 g1000(.A(new_n1198), .B(new_n1200), .C1(G107), .C2(new_n752), .ZN(new_n1201));
  INV_X1    g1001(.A(G41), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n745), .A2(new_n251), .B1(new_n335), .B2(new_n746), .ZN(new_n1203));
  XOR2_X1   g1003(.A(new_n1203), .B(KEYINPUT114), .Z(new_n1204));
  NAND4_X1  g1004(.A1(new_n1201), .A2(new_n1202), .A3(new_n386), .A4(new_n1204), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(new_n1205), .B(KEYINPUT116), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT58), .ZN(new_n1207));
  OR2_X1    g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n745), .A2(new_n820), .B1(new_n813), .B2(new_n746), .ZN(new_n1210));
  XOR2_X1   g1010(.A(new_n1210), .B(KEYINPUT117), .Z(new_n1211));
  OAI22_X1  g1011(.A1(new_n768), .A2(new_n1159), .B1(new_n473), .B2(new_n735), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(G125), .B2(new_n749), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n1211), .B(new_n1213), .C1(new_n754), .C2(new_n1156), .ZN(new_n1214));
  XOR2_X1   g1014(.A(new_n1214), .B(KEYINPUT59), .Z(new_n1215));
  AOI21_X1  g1015(.A(G41), .B1(new_n733), .B2(G124), .ZN(new_n1216));
  AOI21_X1  g1016(.A(G33), .B1(new_n1004), .B2(G159), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1215), .A2(new_n1216), .A3(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(KEYINPUT3), .A2(G33), .ZN(new_n1219));
  AOI21_X1  g1019(.A(G50), .B1(new_n1219), .B2(new_n1202), .ZN(new_n1220));
  XOR2_X1   g1020(.A(new_n1220), .B(KEYINPUT113), .Z(new_n1221));
  NAND4_X1  g1021(.A1(new_n1208), .A2(new_n1209), .A3(new_n1218), .A4(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n723), .B1(new_n1222), .B2(new_n772), .ZN(new_n1223));
  OAI221_X1 g1023(.A(new_n1223), .B1(G50), .B2(new_n1168), .C1(new_n1183), .C2(new_n774), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1196), .A2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1126), .A2(KEYINPUT118), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT118), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n895), .A2(new_n1227), .A3(new_n661), .A4(new_n1125), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1226), .A2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1230), .B1(new_n1140), .B2(new_n1146), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(new_n1195), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT57), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n689), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1231), .A2(KEYINPUT57), .A3(new_n1195), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1225), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(G375));
  NAND3_X1  g1037(.A1(new_n1132), .A2(new_n1135), .A3(new_n1126), .ZN(new_n1238));
  AND2_X1   g1038(.A1(new_n1146), .A2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n977), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  XNOR2_X1  g1041(.A(new_n1241), .B(KEYINPUT119), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n1159), .A2(new_n732), .B1(new_n735), .B2(new_n202), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n273), .B1(new_n738), .B2(new_n362), .ZN(new_n1244));
  XOR2_X1   g1044(.A(new_n1244), .B(KEYINPUT122), .Z(new_n1245));
  AOI211_X1 g1045(.A(new_n1243), .B(new_n1245), .C1(G159), .C2(new_n755), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n744), .A2(new_n1155), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n749), .A2(G132), .ZN(new_n1248));
  XNOR2_X1  g1048(.A(new_n1248), .B(KEYINPUT121), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(G137), .A2(new_n752), .B1(new_n1090), .B2(G150), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1246), .A2(new_n1247), .A3(new_n1249), .A4(new_n1250), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(G107), .A2(new_n1090), .B1(new_n749), .B2(G294), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1252), .B1(new_n208), .B2(new_n745), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT120), .ZN(new_n1254));
  OR2_X1    g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1256));
  OAI221_X1 g1056(.A(new_n386), .B1(new_n735), .B2(new_n335), .C1(new_n251), .C2(new_n754), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n739), .A2(new_n256), .ZN(new_n1258));
  AOI211_X1 g1058(.A(new_n1257), .B(new_n1258), .C1(G283), .C2(new_n752), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1255), .A2(new_n1256), .A3(new_n1259), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n732), .A2(new_n1015), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1251), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(new_n772), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1263), .B1(G68), .B2(new_n1168), .ZN(new_n1264));
  AOI211_X1 g1064(.A(new_n723), .B(new_n1264), .C1(new_n845), .C2(new_n773), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1265), .B1(new_n1144), .B2(new_n929), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1242), .A2(new_n1266), .ZN(G381));
  NOR2_X1   g1067(.A1(G381), .A2(G384), .ZN(new_n1268));
  NOR3_X1   g1068(.A1(new_n1029), .A2(new_n1031), .A3(G390), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(G393), .A2(G396), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1196), .A2(new_n1148), .A3(new_n1171), .A4(new_n1224), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1271), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1268), .A2(new_n1269), .A3(new_n1270), .A4(new_n1272), .ZN(G407));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n669), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(G407), .A2(G213), .A3(new_n1274), .ZN(G409));
  NOR2_X1   g1075(.A1(new_n1232), .A2(new_n977), .ZN(new_n1276));
  OR2_X1    g1076(.A1(new_n1271), .A2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT123), .ZN(new_n1278));
  OAI211_X1 g1078(.A(new_n1277), .B(new_n1278), .C1(new_n1236), .C2(new_n1172), .ZN(new_n1279));
  AND3_X1   g1079(.A1(new_n1193), .A2(new_n894), .A3(new_n1188), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n894), .B1(new_n1193), .B2(new_n1188), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1229), .B1(new_n1124), .B2(new_n1136), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1233), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1284), .A2(new_n1235), .A3(new_n688), .ZN(new_n1285));
  AND2_X1   g1085(.A1(new_n1196), .A2(new_n1224), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1172), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1271), .A2(new_n1276), .ZN(new_n1288));
  OAI21_X1  g1088(.A(KEYINPUT123), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(G213), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1290), .A2(G343), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT60), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1238), .A2(new_n1293), .ZN(new_n1294));
  OAI211_X1 g1094(.A(new_n688), .B(new_n1294), .C1(new_n1239), .C2(new_n1293), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(new_n1266), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1296), .A2(new_n811), .A3(new_n838), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1295), .A2(G384), .A3(new_n1266), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1299), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1279), .A2(new_n1289), .A3(new_n1292), .A4(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT63), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT124), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1299), .A2(new_n1302), .ZN(new_n1306));
  NOR3_X1   g1106(.A1(new_n1287), .A2(new_n1288), .A3(new_n1291), .ZN(new_n1307));
  AOI21_X1  g1107(.A(KEYINPUT61), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1291), .A2(G2897), .ZN(new_n1309));
  XNOR2_X1  g1109(.A(new_n1299), .B(new_n1309), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1279), .A2(new_n1289), .A3(new_n1292), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1000), .A2(new_n1028), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1312), .A2(G390), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1000), .A2(new_n1098), .A3(new_n1102), .A4(new_n1028), .ZN(new_n1314));
  XOR2_X1   g1114(.A(G393), .B(G396), .Z(new_n1315));
  NAND3_X1  g1115(.A1(new_n1313), .A2(new_n1314), .A3(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(KEYINPUT125), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT125), .ZN(new_n1318));
  NAND4_X1  g1118(.A1(new_n1313), .A2(new_n1314), .A3(new_n1318), .A4(new_n1315), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1317), .A2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1315), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1313), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1321), .B1(new_n1269), .B2(new_n1322), .ZN(new_n1323));
  AOI22_X1  g1123(.A1(new_n1310), .A2(new_n1311), .B1(new_n1320), .B2(new_n1323), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1301), .A2(KEYINPUT124), .A3(new_n1302), .ZN(new_n1325));
  NAND4_X1  g1125(.A1(new_n1305), .A2(new_n1308), .A3(new_n1324), .A4(new_n1325), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT62), .ZN(new_n1327));
  NOR2_X1   g1127(.A1(new_n1299), .A2(new_n1327), .ZN(new_n1328));
  AOI22_X1  g1128(.A1(new_n1301), .A2(new_n1327), .B1(new_n1307), .B2(new_n1328), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT61), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n1309), .ZN(new_n1331));
  XNOR2_X1  g1131(.A(new_n1299), .B(new_n1331), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1330), .B1(new_n1332), .B2(new_n1307), .ZN(new_n1333));
  AND3_X1   g1133(.A1(new_n1320), .A2(KEYINPUT126), .A3(new_n1323), .ZN(new_n1334));
  AOI21_X1  g1134(.A(KEYINPUT126), .B1(new_n1320), .B2(new_n1323), .ZN(new_n1335));
  OAI22_X1  g1135(.A1(new_n1329), .A2(new_n1333), .B1(new_n1334), .B2(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1326), .A2(new_n1336), .ZN(G405));
  NAND2_X1  g1137(.A1(new_n1300), .A2(KEYINPUT127), .ZN(new_n1338));
  NOR2_X1   g1138(.A1(new_n1287), .A2(new_n1272), .ZN(new_n1339));
  AND2_X1   g1139(.A1(new_n1338), .A2(new_n1339), .ZN(new_n1340));
  NOR2_X1   g1140(.A1(new_n1338), .A2(new_n1339), .ZN(new_n1341));
  NOR2_X1   g1141(.A1(new_n1340), .A2(new_n1341), .ZN(new_n1342));
  AND2_X1   g1142(.A1(new_n1320), .A2(new_n1323), .ZN(new_n1343));
  XNOR2_X1  g1143(.A(new_n1342), .B(new_n1343), .ZN(G402));
endmodule


