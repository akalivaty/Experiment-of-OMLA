//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 0 1 1 1 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 1 1 1 0 1 0 0 0 0 0 0 1 0 1 0 1 1 0 1 0 0 0 1 0 1 0 1 0 1 0 1 1 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:16 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n548, new_n550, new_n551,
    new_n552, new_n553, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n600, new_n601, new_n604,
    new_n606, new_n607, new_n608, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1149, new_n1150, new_n1151, new_n1152;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT64), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT65), .Z(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  OAI211_X1 g038(.A(G137), .B(new_n461), .C1(new_n462), .C2(new_n463), .ZN(new_n464));
  AND2_X1   g039(.A1(new_n461), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G101), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT66), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n464), .A2(new_n466), .A3(KEYINPUT66), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n462), .A2(new_n463), .ZN(new_n472));
  INV_X1    g047(.A(G125), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AOI22_X1  g049(.A1(new_n469), .A2(new_n470), .B1(G2105), .B2(new_n474), .ZN(G160));
  XNOR2_X1  g050(.A(KEYINPUT3), .B(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G2105), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n472), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n479), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  AND2_X1   g060(.A1(new_n465), .A2(G102), .ZN(new_n486));
  OAI21_X1  g061(.A(G126), .B1(new_n462), .B2(new_n463), .ZN(new_n487));
  NAND2_X1  g062(.A1(G114), .A2(G2104), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n486), .B1(new_n489), .B2(G2105), .ZN(new_n490));
  OAI211_X1 g065(.A(G138), .B(new_n461), .C1(new_n462), .C2(new_n463), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT4), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n476), .A2(new_n493), .A3(G138), .A4(new_n461), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n490), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G164));
  INV_X1    g072(.A(G651), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT6), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT6), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G651), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G50), .ZN(new_n505));
  INV_X1    g080(.A(new_n502), .ZN(new_n506));
  NAND2_X1  g081(.A1(KEYINPUT67), .A2(KEYINPUT5), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(new_n503), .ZN(new_n508));
  NAND3_X1  g083(.A1(KEYINPUT67), .A2(KEYINPUT5), .A3(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G88), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT68), .ZN(new_n514));
  AND2_X1   g089(.A1(new_n508), .A2(new_n509), .ZN(new_n515));
  INV_X1    g090(.A(G62), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(G75), .A2(G543), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n510), .A2(KEYINPUT68), .A3(G62), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  AND3_X1   g095(.A1(new_n520), .A2(KEYINPUT69), .A3(G651), .ZN(new_n521));
  AOI21_X1  g096(.A(KEYINPUT69), .B1(new_n520), .B2(G651), .ZN(new_n522));
  OAI211_X1 g097(.A(new_n505), .B(new_n513), .C1(new_n521), .C2(new_n522), .ZN(G303));
  INV_X1    g098(.A(G303), .ZN(G166));
  NAND2_X1  g099(.A1(new_n504), .A2(G51), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n510), .A2(G63), .A3(G651), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT7), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n525), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n529), .B1(G89), .B2(new_n512), .ZN(new_n530));
  OR2_X1    g105(.A1(new_n530), .A2(KEYINPUT70), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(KEYINPUT70), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(G168));
  NAND2_X1  g108(.A1(new_n504), .A2(G52), .ZN(new_n534));
  INV_X1    g109(.A(G90), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n534), .B1(new_n535), .B2(new_n511), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n510), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n498), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n536), .A2(new_n538), .ZN(G171));
  NAND2_X1  g114(.A1(new_n504), .A2(G43), .ZN(new_n540));
  INV_X1    g115(.A(G81), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n540), .B1(new_n541), .B2(new_n511), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n510), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n543), .A2(new_n498), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G860), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT71), .ZN(G153));
  AND3_X1   g122(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G36), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT73), .ZN(new_n551));
  XOR2_X1   g126(.A(KEYINPUT72), .B(KEYINPUT8), .Z(new_n552));
  XNOR2_X1  g127(.A(new_n551), .B(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n548), .A2(new_n553), .ZN(G188));
  NAND2_X1  g129(.A1(new_n506), .A2(G543), .ZN(new_n555));
  INV_X1    g130(.A(G53), .ZN(new_n556));
  OAI21_X1  g131(.A(KEYINPUT9), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT9), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n504), .A2(new_n558), .A3(G53), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n510), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n561));
  OR2_X1    g136(.A1(new_n561), .A2(new_n498), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n512), .A2(G91), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n560), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  XOR2_X1   g139(.A(new_n564), .B(KEYINPUT74), .Z(G299));
  INV_X1    g140(.A(G171), .ZN(G301));
  INV_X1    g141(.A(G168), .ZN(G286));
  OR2_X1    g142(.A1(new_n510), .A2(G74), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n568), .A2(G651), .B1(new_n504), .B2(G49), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n512), .A2(G87), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(G288));
  NAND2_X1  g146(.A1(new_n504), .A2(G48), .ZN(new_n572));
  INV_X1    g147(.A(G86), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n573), .B2(new_n511), .ZN(new_n574));
  NAND2_X1  g149(.A1(G73), .A2(G543), .ZN(new_n575));
  XOR2_X1   g150(.A(new_n575), .B(KEYINPUT75), .Z(new_n576));
  NAND2_X1  g151(.A1(new_n510), .A2(G61), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n498), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n574), .A2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(G305));
  NAND2_X1  g155(.A1(new_n504), .A2(G47), .ZN(new_n581));
  INV_X1    g156(.A(G85), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n582), .B2(new_n511), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT76), .ZN(new_n584));
  AND2_X1   g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n583), .A2(new_n584), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n510), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n587));
  OAI22_X1  g162(.A1(new_n585), .A2(new_n586), .B1(new_n498), .B2(new_n587), .ZN(G290));
  NAND2_X1  g163(.A1(G301), .A2(G868), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n512), .A2(G92), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n590), .B(KEYINPUT10), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n510), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n592), .A2(new_n498), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n504), .A2(G54), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n589), .B1(new_n597), .B2(G868), .ZN(G284));
  OAI21_X1  g173(.A(new_n589), .B1(new_n597), .B2(G868), .ZN(G321));
  INV_X1    g174(.A(G868), .ZN(new_n600));
  NAND2_X1  g175(.A1(G299), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n601), .B1(new_n600), .B2(G168), .ZN(G297));
  OAI21_X1  g177(.A(new_n601), .B1(new_n600), .B2(G168), .ZN(G280));
  INV_X1    g178(.A(G559), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n597), .B1(new_n604), .B2(G860), .ZN(G148));
  INV_X1    g180(.A(new_n545), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(new_n600), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n596), .A2(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(new_n600), .ZN(G323));
  XNOR2_X1  g184(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g185(.A1(new_n476), .A2(new_n465), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT12), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT13), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(G2100), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n478), .A2(G123), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n480), .A2(G135), .ZN(new_n616));
  NOR2_X1   g191(.A1(G99), .A2(G2105), .ZN(new_n617));
  OAI21_X1  g192(.A(G2104), .B1(new_n461), .B2(G111), .ZN(new_n618));
  OAI211_X1 g193(.A(new_n615), .B(new_n616), .C1(new_n617), .C2(new_n618), .ZN(new_n619));
  XNOR2_X1  g194(.A(KEYINPUT77), .B(G2096), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n619), .B(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n614), .A2(new_n621), .ZN(G156));
  XNOR2_X1  g197(.A(KEYINPUT15), .B(G2430), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(G2435), .ZN(new_n624));
  XOR2_X1   g199(.A(G2427), .B(G2438), .Z(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(KEYINPUT14), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(KEYINPUT79), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT16), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2451), .B(G2454), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT78), .ZN(new_n631));
  XNOR2_X1  g206(.A(G2443), .B(G2446), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(G1341), .B(G1348), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n629), .B(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(G14), .ZN(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(G401));
  XOR2_X1   g213(.A(G2084), .B(G2090), .Z(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G2067), .B(G2678), .Z(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n642), .A2(new_n643), .A3(KEYINPUT17), .ZN(new_n644));
  XOR2_X1   g219(.A(KEYINPUT80), .B(KEYINPUT18), .Z(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G2072), .B(G2078), .Z(new_n648));
  AOI21_X1  g223(.A(new_n648), .B1(new_n642), .B2(new_n645), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n647), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2096), .B(G2100), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(G227));
  XOR2_X1   g227(.A(G1956), .B(G2474), .Z(new_n653));
  XOR2_X1   g228(.A(G1961), .B(G1966), .Z(new_n654));
  AND2_X1   g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n655), .A2(KEYINPUT81), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1971), .B(G1976), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT19), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n655), .A2(KEYINPUT81), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n656), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(KEYINPUT20), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n653), .A2(new_n654), .ZN(new_n664));
  OR3_X1    g239(.A1(new_n659), .A2(new_n655), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n661), .A2(new_n662), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n659), .A2(new_n664), .ZN(new_n667));
  NAND4_X1  g242(.A1(new_n663), .A2(new_n665), .A3(new_n666), .A4(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G1991), .B(G1996), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1981), .B(G1986), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(G229));
  NAND2_X1  g249(.A1(new_n478), .A2(G119), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n480), .A2(G131), .ZN(new_n676));
  NOR2_X1   g251(.A1(G95), .A2(G2105), .ZN(new_n677));
  OAI21_X1  g252(.A(G2104), .B1(new_n461), .B2(G107), .ZN(new_n678));
  OAI211_X1 g253(.A(new_n675), .B(new_n676), .C1(new_n677), .C2(new_n678), .ZN(new_n679));
  MUX2_X1   g254(.A(G25), .B(new_n679), .S(G29), .Z(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT35), .B(G1991), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(G16), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n683), .A2(G23), .ZN(new_n684));
  INV_X1    g259(.A(G288), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n684), .B1(new_n685), .B2(new_n683), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT33), .ZN(new_n687));
  INV_X1    g262(.A(G1976), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n683), .A2(G22), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n690), .B1(G166), .B2(new_n683), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n689), .B1(G1971), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n683), .A2(G6), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n693), .B1(new_n579), .B2(new_n683), .ZN(new_n694));
  XOR2_X1   g269(.A(KEYINPUT32), .B(G1981), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  OAI211_X1 g271(.A(new_n692), .B(new_n696), .C1(G1971), .C2(new_n691), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n682), .B1(new_n697), .B2(KEYINPUT34), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n683), .A2(G24), .ZN(new_n699));
  INV_X1    g274(.A(G290), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n699), .B1(new_n700), .B2(new_n683), .ZN(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT82), .B(G1986), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT83), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n701), .B(new_n703), .ZN(new_n704));
  OAI211_X1 g279(.A(new_n698), .B(new_n704), .C1(KEYINPUT34), .C2(new_n697), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT36), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n683), .A2(G21), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(G168), .B2(new_n683), .ZN(new_n708));
  XOR2_X1   g283(.A(KEYINPUT90), .B(G1966), .Z(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(G29), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G35), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(G162), .B2(new_n711), .ZN(new_n713));
  MUX2_X1   g288(.A(new_n712), .B(new_n713), .S(KEYINPUT92), .Z(new_n714));
  XOR2_X1   g289(.A(KEYINPUT29), .B(G2090), .Z(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  NOR2_X1   g291(.A1(G164), .A2(new_n711), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(G27), .B2(new_n711), .ZN(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n716), .B1(G2078), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(G160), .A2(G29), .ZN(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT88), .B(KEYINPUT24), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(G34), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(new_n711), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n721), .A2(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n683), .A2(G5), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(G171), .B2(new_n683), .ZN(new_n728));
  AOI22_X1  g303(.A1(new_n726), .A2(G2084), .B1(G1961), .B2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(G2084), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n725), .A2(new_n730), .ZN(new_n731));
  OAI211_X1 g306(.A(new_n729), .B(new_n731), .C1(G1961), .C2(new_n728), .ZN(new_n732));
  OR2_X1    g307(.A1(G29), .A2(G32), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n478), .A2(G129), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n465), .A2(G105), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n480), .A2(G141), .ZN(new_n736));
  NAND3_X1  g311(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT26), .Z(new_n738));
  NAND4_X1  g313(.A1(new_n734), .A2(new_n735), .A3(new_n736), .A4(new_n738), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n733), .B1(new_n739), .B2(new_n711), .ZN(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT27), .B(G1996), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT89), .Z(new_n743));
  NAND2_X1  g318(.A1(new_n719), .A2(G2078), .ZN(new_n744));
  OR2_X1    g319(.A1(new_n740), .A2(new_n741), .ZN(new_n745));
  OR2_X1    g320(.A1(new_n619), .A2(new_n711), .ZN(new_n746));
  INV_X1    g321(.A(KEYINPUT30), .ZN(new_n747));
  AND3_X1   g322(.A1(new_n747), .A2(KEYINPUT91), .A3(G28), .ZN(new_n748));
  AOI21_X1  g323(.A(KEYINPUT91), .B1(new_n747), .B2(G28), .ZN(new_n749));
  OAI221_X1 g324(.A(new_n711), .B1(new_n747), .B2(G28), .C1(new_n748), .C2(new_n749), .ZN(new_n750));
  AND3_X1   g325(.A1(new_n745), .A2(new_n746), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n683), .A2(G19), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(new_n545), .B2(new_n683), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n753), .A2(G1341), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n753), .A2(G1341), .ZN(new_n755));
  NAND4_X1  g330(.A1(new_n744), .A2(new_n751), .A3(new_n754), .A4(new_n755), .ZN(new_n756));
  NOR4_X1   g331(.A1(new_n720), .A2(new_n732), .A3(new_n743), .A4(new_n756), .ZN(new_n757));
  XNOR2_X1  g332(.A(KEYINPUT31), .B(G11), .ZN(new_n758));
  OAI21_X1  g333(.A(KEYINPUT86), .B1(G29), .B2(G33), .ZN(new_n759));
  OR3_X1    g334(.A1(KEYINPUT86), .A2(G29), .A3(G33), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n480), .A2(G139), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT87), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n465), .A2(G103), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT25), .Z(new_n764));
  AOI22_X1  g339(.A1(new_n476), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n765));
  OAI211_X1 g340(.A(new_n762), .B(new_n764), .C1(new_n461), .C2(new_n765), .ZN(new_n766));
  OAI211_X1 g341(.A(new_n759), .B(new_n760), .C1(new_n766), .C2(new_n711), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(G2072), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n683), .A2(G4), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(new_n597), .B2(new_n683), .ZN(new_n770));
  INV_X1    g345(.A(G1348), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  NAND4_X1  g347(.A1(new_n757), .A2(new_n758), .A3(new_n768), .A4(new_n772), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT93), .B(KEYINPUT23), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n683), .A2(G20), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(G299), .B2(G16), .ZN(new_n777));
  INV_X1    g352(.A(G1956), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n711), .A2(G26), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(KEYINPUT85), .Z(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT28), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n478), .A2(G128), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n480), .A2(G140), .ZN(new_n784));
  NOR2_X1   g359(.A1(G104), .A2(G2105), .ZN(new_n785));
  OAI21_X1  g360(.A(G2104), .B1(new_n461), .B2(G116), .ZN(new_n786));
  OAI211_X1 g361(.A(new_n783), .B(new_n784), .C1(new_n785), .C2(new_n786), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT84), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n782), .B1(new_n788), .B2(G29), .ZN(new_n789));
  INV_X1    g364(.A(G2067), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NOR3_X1   g366(.A1(new_n773), .A2(new_n779), .A3(new_n791), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n706), .A2(new_n710), .A3(new_n792), .ZN(G150));
  INV_X1    g368(.A(G150), .ZN(G311));
  AOI22_X1  g369(.A1(new_n510), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n795), .A2(new_n498), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT94), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n512), .A2(G93), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n504), .A2(G55), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n797), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n800), .A2(G860), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(KEYINPUT37), .Z(new_n802));
  NOR2_X1   g377(.A1(new_n596), .A2(new_n604), .ZN(new_n803));
  XNOR2_X1  g378(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  AND3_X1   g380(.A1(new_n797), .A2(new_n798), .A3(new_n799), .ZN(new_n806));
  AOI21_X1  g381(.A(KEYINPUT96), .B1(new_n806), .B2(new_n606), .ZN(new_n807));
  INV_X1    g382(.A(KEYINPUT96), .ZN(new_n808));
  NOR3_X1   g383(.A1(new_n800), .A2(new_n808), .A3(new_n545), .ZN(new_n809));
  AND3_X1   g384(.A1(new_n800), .A2(KEYINPUT95), .A3(new_n545), .ZN(new_n810));
  AOI21_X1  g385(.A(KEYINPUT95), .B1(new_n800), .B2(new_n545), .ZN(new_n811));
  OAI22_X1  g386(.A1(new_n807), .A2(new_n809), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n805), .B(new_n812), .Z(new_n813));
  OAI21_X1  g388(.A(new_n802), .B1(new_n813), .B2(G860), .ZN(G145));
  XOR2_X1   g389(.A(new_n619), .B(G160), .Z(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(new_n484), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n788), .B(new_n766), .Z(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(new_n739), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(new_n612), .Z(new_n819));
  AND3_X1   g394(.A1(new_n490), .A2(KEYINPUT97), .A3(new_n495), .ZN(new_n820));
  AOI21_X1  g395(.A(KEYINPUT97), .B1(new_n490), .B2(new_n495), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(G130), .ZN(new_n823));
  NOR2_X1   g398(.A1(G106), .A2(G2105), .ZN(new_n824));
  OAI21_X1  g399(.A(G2104), .B1(new_n461), .B2(G118), .ZN(new_n825));
  OAI22_X1  g400(.A1(new_n477), .A2(new_n823), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n826), .B1(G142), .B2(new_n480), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n822), .B(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(new_n679), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n819), .A2(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n819), .A2(new_n829), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n816), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(new_n832), .ZN(new_n834));
  INV_X1    g409(.A(new_n816), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n834), .A2(new_n830), .A3(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(G37), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n833), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g414(.A(G299), .B(new_n596), .ZN(new_n840));
  XOR2_X1   g415(.A(KEYINPUT98), .B(KEYINPUT41), .Z(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n842), .B1(KEYINPUT41), .B2(new_n840), .ZN(new_n843));
  AND2_X1   g418(.A1(new_n812), .A2(new_n608), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n812), .A2(new_n608), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n840), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n848), .B1(new_n844), .B2(new_n845), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(KEYINPUT99), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n579), .B(G288), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n700), .B(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(G166), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT100), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT42), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n856), .A2(new_n857), .ZN(new_n859));
  NAND2_X1  g434(.A1(KEYINPUT100), .A2(KEYINPUT42), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n854), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(KEYINPUT99), .B1(new_n843), .B2(new_n846), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n851), .A2(new_n863), .A3(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT99), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n867), .B1(new_n847), .B2(new_n849), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n862), .B1(new_n868), .B2(new_n864), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n866), .A2(new_n869), .A3(KEYINPUT101), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT101), .ZN(new_n871));
  OAI211_X1 g446(.A(new_n871), .B(new_n862), .C1(new_n868), .C2(new_n864), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n600), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n800), .A2(G868), .ZN(new_n874));
  OR3_X1    g449(.A1(new_n873), .A2(KEYINPUT102), .A3(new_n874), .ZN(new_n875));
  OAI21_X1  g450(.A(KEYINPUT102), .B1(new_n873), .B2(new_n874), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(G295));
  INV_X1    g452(.A(KEYINPUT103), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n870), .A2(new_n872), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n879), .A2(G868), .ZN(new_n880));
  INV_X1    g455(.A(new_n874), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n878), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NOR3_X1   g457(.A1(new_n873), .A2(KEYINPUT103), .A3(new_n874), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n882), .A2(new_n883), .ZN(G331));
  INV_X1    g459(.A(KEYINPUT44), .ZN(new_n885));
  XNOR2_X1  g460(.A(KEYINPUT104), .B(KEYINPUT43), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  XOR2_X1   g462(.A(G168), .B(KEYINPUT105), .Z(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n812), .A2(G171), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n812), .A2(G171), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n889), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  OR2_X1    g468(.A1(new_n812), .A2(G171), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n894), .A2(new_n888), .A3(new_n890), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n896), .A2(new_n848), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n843), .B1(new_n893), .B2(new_n895), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n855), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  AND2_X1   g474(.A1(new_n899), .A2(new_n837), .ZN(new_n900));
  OR3_X1    g475(.A1(new_n897), .A2(new_n855), .A3(new_n898), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n887), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n899), .A2(new_n837), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n896), .A2(new_n841), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(new_n848), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n840), .A2(KEYINPUT41), .ZN(new_n906));
  XOR2_X1   g481(.A(new_n906), .B(KEYINPUT106), .Z(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(new_n896), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n855), .B1(new_n905), .B2(new_n908), .ZN(new_n909));
  NOR3_X1   g484(.A1(new_n903), .A2(new_n909), .A3(new_n886), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n885), .B1(new_n902), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(KEYINPUT43), .B1(new_n903), .B2(new_n909), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(KEYINPUT107), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT107), .ZN(new_n914));
  OAI211_X1 g489(.A(new_n914), .B(KEYINPUT43), .C1(new_n903), .C2(new_n909), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n913), .A2(KEYINPUT44), .A3(new_n915), .ZN(new_n916));
  AND3_X1   g491(.A1(new_n900), .A2(new_n887), .A3(new_n901), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n911), .B1(new_n916), .B2(new_n917), .ZN(G397));
  INV_X1    g493(.A(KEYINPUT45), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n919), .B1(new_n822), .B2(G1384), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n474), .A2(G2105), .ZN(new_n921));
  INV_X1    g496(.A(new_n470), .ZN(new_n922));
  AOI21_X1  g497(.A(KEYINPUT66), .B1(new_n464), .B2(new_n466), .ZN(new_n923));
  OAI211_X1 g498(.A(G40), .B(new_n921), .C1(new_n922), .C2(new_n923), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n920), .A2(new_n924), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n788), .B(new_n790), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n926), .B(KEYINPUT109), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n925), .B1(new_n927), .B2(new_n739), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT46), .ZN(new_n929));
  INV_X1    g504(.A(new_n925), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n929), .B1(new_n930), .B2(G1996), .ZN(new_n931));
  INV_X1    g506(.A(G1996), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n925), .A2(KEYINPUT46), .A3(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n928), .A2(new_n931), .A3(new_n933), .ZN(new_n934));
  XOR2_X1   g509(.A(new_n934), .B(KEYINPUT47), .Z(new_n935));
  XNOR2_X1  g510(.A(new_n739), .B(G1996), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n927), .A2(new_n936), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n679), .A2(new_n681), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  OR2_X1    g514(.A1(new_n788), .A2(G2067), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n930), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n941), .B(KEYINPUT127), .ZN(new_n942));
  XOR2_X1   g517(.A(new_n679), .B(new_n681), .Z(new_n943));
  NAND2_X1  g518(.A1(new_n937), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(new_n925), .ZN(new_n945));
  NOR2_X1   g520(.A1(G290), .A2(G1986), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n925), .A2(new_n946), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n947), .B(KEYINPUT48), .ZN(new_n948));
  AOI211_X1 g523(.A(new_n935), .B(new_n942), .C1(new_n945), .C2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT126), .ZN(new_n950));
  INV_X1    g525(.A(new_n946), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT108), .ZN(new_n952));
  NAND2_X1  g527(.A1(G290), .A2(G1986), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n951), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  OAI211_X1 g529(.A(new_n954), .B(new_n925), .C1(new_n952), .C2(new_n953), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n945), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(KEYINPUT111), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT55), .ZN(new_n959));
  INV_X1    g534(.A(G8), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n959), .B1(G166), .B2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT111), .ZN(new_n962));
  NAND4_X1  g537(.A1(G303), .A2(new_n962), .A3(KEYINPUT55), .A4(G8), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n958), .A2(new_n961), .A3(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT110), .ZN(new_n965));
  INV_X1    g540(.A(G1384), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n496), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n924), .B1(new_n967), .B2(KEYINPUT50), .ZN(new_n968));
  AOI21_X1  g543(.A(G1384), .B1(new_n490), .B2(new_n495), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT50), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n968), .A2(new_n971), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n965), .B1(new_n972), .B2(G2090), .ZN(new_n973));
  INV_X1    g548(.A(G2090), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n968), .A2(KEYINPUT110), .A3(new_n974), .A4(new_n971), .ZN(new_n975));
  OAI211_X1 g550(.A(KEYINPUT45), .B(new_n966), .C1(new_n820), .C2(new_n821), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n924), .B1(new_n967), .B2(new_n919), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(G1971), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n973), .A2(new_n975), .A3(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n964), .A2(G8), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(G305), .A2(G1981), .ZN(new_n983));
  OR3_X1    g558(.A1(new_n574), .A2(G1981), .A3(new_n578), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT49), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(new_n924), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(new_n969), .ZN(new_n989));
  INV_X1    g564(.A(new_n989), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n990), .A2(new_n960), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n983), .A2(KEYINPUT49), .A3(new_n984), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n987), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n569), .A2(new_n570), .A3(KEYINPUT112), .A4(G1976), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n989), .A2(G8), .A3(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(KEYINPUT52), .B1(G288), .B2(new_n688), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT114), .ZN(new_n998));
  OR2_X1    g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT112), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n1000), .B1(G288), .B2(new_n688), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n997), .A2(new_n998), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n996), .A2(new_n999), .A3(new_n1001), .A4(new_n1002), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n1001), .A2(new_n989), .A3(G8), .A4(new_n994), .ZN(new_n1004));
  AND3_X1   g579(.A1(new_n1004), .A2(KEYINPUT113), .A3(KEYINPUT52), .ZN(new_n1005));
  AOI21_X1  g580(.A(KEYINPUT113), .B1(new_n1004), .B2(KEYINPUT52), .ZN(new_n1006));
  OAI211_X1 g581(.A(new_n993), .B(new_n1003), .C1(new_n1005), .C2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n982), .A2(new_n1007), .ZN(new_n1008));
  AND3_X1   g583(.A1(new_n958), .A2(new_n961), .A3(new_n963), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT115), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n971), .A2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n969), .A2(KEYINPUT115), .A3(new_n970), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1013), .A2(new_n974), .A3(new_n968), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1014), .A2(new_n980), .A3(KEYINPUT116), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(G8), .ZN(new_n1016));
  AOI21_X1  g591(.A(KEYINPUT116), .B1(new_n1014), .B2(new_n980), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1009), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1007), .ZN(new_n1019));
  INV_X1    g594(.A(G1966), .ZN(new_n1020));
  OAI211_X1 g595(.A(G40), .B(G160), .C1(new_n969), .C2(KEYINPUT45), .ZN(new_n1021));
  AOI211_X1 g596(.A(new_n919), .B(G1384), .C1(new_n490), .C2(new_n495), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1020), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(KEYINPUT117), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n968), .A2(new_n730), .A3(new_n971), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT117), .ZN(new_n1026));
  OAI211_X1 g601(.A(new_n1026), .B(new_n1020), .C1(new_n1021), .C2(new_n1022), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1024), .A2(new_n1025), .A3(new_n1027), .ZN(new_n1028));
  AND3_X1   g603(.A1(new_n1028), .A2(G8), .A3(G168), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1018), .A2(new_n982), .A3(new_n1019), .A4(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT63), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n981), .A2(G8), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1031), .B1(new_n1009), .B2(new_n1033), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1034), .A2(new_n982), .A3(new_n1019), .A4(new_n1029), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1032), .A2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n993), .A2(new_n688), .A3(new_n685), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(new_n984), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(new_n991), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1036), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT61), .ZN(new_n1041));
  OR2_X1    g616(.A1(new_n1041), .A2(KEYINPUT121), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(KEYINPUT121), .ZN(new_n1043));
  AOI21_X1  g618(.A(G1956), .B1(new_n1013), .B2(new_n968), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT118), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT57), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n560), .A2(new_n562), .A3(new_n563), .A4(new_n1047), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1049));
  XNOR2_X1  g624(.A(new_n1048), .B(new_n1049), .ZN(new_n1050));
  XNOR2_X1  g625(.A(KEYINPUT56), .B(G2072), .ZN(new_n1051));
  AND3_X1   g626(.A1(new_n976), .A2(new_n977), .A3(new_n1051), .ZN(new_n1052));
  NOR3_X1   g627(.A1(new_n1044), .A2(new_n1050), .A3(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1049), .ZN(new_n1054));
  XNOR2_X1  g629(.A(new_n1048), .B(new_n1054), .ZN(new_n1055));
  AND3_X1   g630(.A1(new_n969), .A2(KEYINPUT115), .A3(new_n970), .ZN(new_n1056));
  AOI21_X1  g631(.A(KEYINPUT115), .B1(new_n969), .B2(new_n970), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n968), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(new_n778), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n976), .A2(new_n977), .A3(new_n1051), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1055), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n1042), .B(new_n1043), .C1(new_n1053), .C2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1050), .B1(new_n1044), .B2(new_n1052), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1059), .A2(new_n1055), .A3(new_n1060), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1063), .A2(KEYINPUT121), .A3(new_n1064), .A4(new_n1041), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1062), .A2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n976), .A2(new_n977), .A3(new_n932), .ZN(new_n1067));
  XOR2_X1   g642(.A(KEYINPUT58), .B(G1341), .Z(new_n1068));
  NAND2_X1  g643(.A1(new_n989), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1070), .A2(KEYINPUT120), .A3(new_n545), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(KEYINPUT59), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1070), .A2(new_n545), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT120), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1072), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1073), .A2(new_n1074), .A3(KEYINPUT59), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT119), .ZN(new_n1079));
  AOI21_X1  g654(.A(G1348), .B1(new_n968), .B2(new_n971), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n989), .A2(G2067), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1079), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  NOR3_X1   g658(.A1(new_n1080), .A2(new_n1081), .A3(new_n1079), .ZN(new_n1084));
  OAI21_X1  g659(.A(KEYINPUT60), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1084), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT60), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1086), .A2(new_n1087), .A3(new_n1082), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1085), .A2(new_n1088), .A3(new_n597), .ZN(new_n1089));
  OAI211_X1 g664(.A(KEYINPUT60), .B(new_n596), .C1(new_n1083), .C2(new_n1084), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1066), .A2(new_n1078), .A3(new_n1089), .A4(new_n1090), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1086), .A2(new_n1064), .A3(new_n597), .A4(new_n1082), .ZN(new_n1092));
  AND3_X1   g667(.A1(new_n1091), .A2(new_n1092), .A3(new_n1063), .ZN(new_n1093));
  AND3_X1   g668(.A1(new_n1018), .A2(new_n982), .A3(new_n1019), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT54), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT53), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1096), .B1(new_n978), .B2(G2078), .ZN(new_n1097));
  INV_X1    g672(.A(G1961), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n972), .A2(new_n1098), .ZN(new_n1099));
  AND2_X1   g674(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1096), .A2(G2078), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n977), .B(new_n1101), .C1(new_n919), .C2(new_n967), .ZN(new_n1102));
  AOI21_X1  g677(.A(G301), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n920), .A2(new_n988), .A3(new_n976), .A4(new_n1101), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1097), .A2(new_n1104), .A3(new_n1099), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1105), .A2(G171), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1095), .B1(new_n1103), .B2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1100), .A2(G301), .A3(new_n1102), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1095), .B1(new_n1105), .B2(G171), .ZN(new_n1109));
  AOI21_X1  g684(.A(KEYINPUT125), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  AND3_X1   g685(.A1(new_n1108), .A2(new_n1109), .A3(KEYINPUT125), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n1094), .B(new_n1107), .C1(new_n1110), .C2(new_n1111), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1093), .A2(new_n1112), .ZN(new_n1113));
  NOR2_X1   g688(.A1(G168), .A2(new_n960), .ZN(new_n1114));
  AOI211_X1 g689(.A(KEYINPUT51), .B(new_n1114), .C1(new_n1028), .C2(G8), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT122), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1028), .A2(new_n1117), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1024), .A2(KEYINPUT122), .A3(new_n1025), .A4(new_n1027), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1118), .A2(G8), .A3(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT123), .ZN(new_n1121));
  XNOR2_X1  g696(.A(new_n1114), .B(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(KEYINPUT124), .B1(new_n1123), .B2(KEYINPUT51), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT51), .ZN(new_n1126));
  AOI211_X1 g701(.A(new_n1125), .B(new_n1126), .C1(new_n1120), .C2(new_n1122), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1116), .B1(new_n1124), .B2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1118), .A2(new_n1114), .A3(new_n1119), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  AOI211_X1 g705(.A(new_n1008), .B(new_n1040), .C1(new_n1113), .C2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1123), .A2(KEYINPUT51), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1132), .A2(new_n1125), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1123), .A2(KEYINPUT124), .A3(KEYINPUT51), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1115), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1129), .ZN(new_n1136));
  OAI21_X1  g711(.A(KEYINPUT62), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT62), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1128), .A2(new_n1138), .A3(new_n1129), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1137), .A2(new_n1094), .A3(new_n1139), .A4(new_n1103), .ZN(new_n1140));
  AOI211_X1 g715(.A(new_n950), .B(new_n956), .C1(new_n1131), .C2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1008), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1040), .B1(new_n1113), .B2(new_n1130), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1140), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(new_n956), .ZN(new_n1145));
  AOI21_X1  g720(.A(KEYINPUT126), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n949), .B1(new_n1141), .B2(new_n1146), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g722(.A1(G229), .A2(new_n459), .ZN(new_n1149));
  OAI21_X1  g723(.A(new_n1149), .B1(new_n902), .B2(new_n910), .ZN(new_n1150));
  INV_X1    g724(.A(G227), .ZN(new_n1151));
  NAND3_X1  g725(.A1(new_n838), .A2(new_n637), .A3(new_n1151), .ZN(new_n1152));
  NOR2_X1   g726(.A1(new_n1150), .A2(new_n1152), .ZN(G308));
  OR2_X1    g727(.A1(new_n1150), .A2(new_n1152), .ZN(G225));
endmodule


