//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 0 1 0 0 1 1 0 1 0 0 1 0 0 0 0 1 1 0 0 0 0 0 0 1 1 1 0 0 0 0 1 1 0 0 0 0 1 0 0 1 1 0 1 1 0 0 1 1 1 1 1 1 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:26 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n577, new_n578,
    new_n579, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n595, new_n596, new_n597,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n629, new_n632,
    new_n634, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT64), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NOR4_X1   g029(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT65), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(new_n454), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G2106), .ZN(new_n460));
  INV_X1    g035(.A(G567), .ZN(new_n461));
  OR2_X1    g036(.A1(new_n455), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G101), .ZN(new_n468));
  XNOR2_X1  g043(.A(KEYINPUT3), .B(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(new_n465), .ZN(new_n470));
  INV_X1    g045(.A(G137), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n468), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT66), .ZN(new_n473));
  AND2_X1   g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  NOR2_X1   g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(G125), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n473), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n469), .A2(KEYINPUT66), .A3(G125), .ZN(new_n479));
  NAND2_X1  g054(.A1(G113), .A2(G2104), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n472), .B1(new_n481), .B2(G2105), .ZN(G160));
  OAI21_X1  g057(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(G112), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n483), .B1(new_n484), .B2(G2105), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT67), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n470), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n469), .A2(KEYINPUT67), .A3(new_n465), .ZN(new_n488));
  AND2_X1   g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AND2_X1   g064(.A1(new_n489), .A2(G136), .ZN(new_n490));
  OR2_X1    g065(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n491));
  NAND2_X1  g066(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n465), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  AOI211_X1 g068(.A(new_n485), .B(new_n490), .C1(G124), .C2(new_n493), .ZN(G162));
  NOR2_X1   g069(.A1(new_n465), .A2(G114), .ZN(new_n495));
  OAI21_X1  g070(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n496));
  OAI21_X1  g071(.A(KEYINPUT68), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  OR2_X1    g072(.A1(G102), .A2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(G114), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(G2105), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT68), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n498), .A2(new_n500), .A3(new_n501), .A4(G2104), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n497), .A2(new_n502), .ZN(new_n503));
  OAI211_X1 g078(.A(G138), .B(new_n465), .C1(new_n474), .C2(new_n475), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT4), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n469), .A2(KEYINPUT4), .A3(G138), .A4(new_n465), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n469), .A2(G126), .A3(G2105), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n503), .A2(new_n506), .A3(new_n507), .A4(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(G164));
  NAND2_X1  g085(.A1(G75), .A2(G543), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT69), .ZN(new_n512));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n512), .B1(new_n513), .B2(KEYINPUT5), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT5), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n515), .A2(KEYINPUT69), .A3(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n513), .A2(KEYINPUT5), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G62), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n511), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G651), .ZN(new_n522));
  XNOR2_X1  g097(.A(KEYINPUT6), .B(G651), .ZN(new_n523));
  XNOR2_X1  g098(.A(KEYINPUT70), .B(G88), .ZN(new_n524));
  NAND4_X1  g099(.A1(new_n517), .A2(new_n518), .A3(new_n523), .A4(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT71), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n523), .A2(G50), .A3(G543), .ZN(new_n527));
  AND3_X1   g102(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n526), .B1(new_n525), .B2(new_n527), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n522), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(KEYINPUT72), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT72), .ZN(new_n532));
  OAI211_X1 g107(.A(new_n522), .B(new_n532), .C1(new_n528), .C2(new_n529), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n531), .A2(new_n533), .ZN(G166));
  INV_X1    g109(.A(KEYINPUT74), .ZN(new_n535));
  AND2_X1   g110(.A1(new_n517), .A2(new_n518), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n536), .A2(G89), .A3(new_n523), .ZN(new_n537));
  AND2_X1   g112(.A1(new_n523), .A2(G543), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G51), .ZN(new_n539));
  AND2_X1   g114(.A1(G63), .A2(G651), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n536), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n537), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  NAND3_X1  g117(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT73), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT7), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n544), .B(new_n545), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n535), .B1(new_n542), .B2(new_n546), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n544), .B(KEYINPUT7), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n536), .A2(new_n540), .B1(new_n538), .B2(G51), .ZN(new_n549));
  NAND4_X1  g124(.A1(new_n548), .A2(new_n549), .A3(KEYINPUT74), .A4(new_n537), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n547), .A2(new_n550), .ZN(G168));
  AND2_X1   g126(.A1(new_n536), .A2(new_n523), .ZN(new_n552));
  XNOR2_X1  g127(.A(KEYINPUT76), .B(G90), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n552), .A2(new_n553), .B1(G52), .B2(new_n538), .ZN(new_n554));
  NAND2_X1  g129(.A1(G77), .A2(G543), .ZN(new_n555));
  INV_X1    g130(.A(G64), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n519), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G651), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(KEYINPUT75), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT75), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n557), .A2(new_n560), .A3(G651), .ZN(new_n561));
  AND3_X1   g136(.A1(new_n554), .A2(new_n559), .A3(new_n561), .ZN(G171));
  NAND2_X1  g137(.A1(G68), .A2(G543), .ZN(new_n563));
  INV_X1    g138(.A(G56), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n519), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G651), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n538), .A2(G43), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n536), .A2(G81), .A3(new_n523), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT77), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n566), .A2(KEYINPUT77), .A3(new_n567), .A4(new_n568), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(G860), .ZN(G153));
  NAND4_X1  g150(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g151(.A1(G1), .A2(G3), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n577), .B(KEYINPUT8), .ZN(new_n578));
  NAND4_X1  g153(.A1(G319), .A2(G483), .A3(G661), .A4(new_n578), .ZN(new_n579));
  XOR2_X1   g154(.A(new_n579), .B(KEYINPUT78), .Z(G188));
  NAND3_X1  g155(.A1(new_n523), .A2(G53), .A3(G543), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n581), .B(KEYINPUT9), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n536), .A2(G91), .A3(new_n523), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(G651), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n536), .A2(G65), .ZN(new_n586));
  NAND2_X1  g161(.A1(G78), .A2(G543), .ZN(new_n587));
  XNOR2_X1  g162(.A(new_n587), .B(KEYINPUT79), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n585), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n584), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(G299));
  NAND3_X1  g166(.A1(new_n554), .A2(new_n559), .A3(new_n561), .ZN(G301));
  INV_X1    g167(.A(G168), .ZN(G286));
  INV_X1    g168(.A(G166), .ZN(G303));
  OAI21_X1  g169(.A(G651), .B1(new_n536), .B2(G74), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n536), .A2(G87), .A3(new_n523), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n538), .A2(G49), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(G288));
  NAND3_X1  g173(.A1(new_n536), .A2(G86), .A3(new_n523), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n538), .A2(G48), .ZN(new_n600));
  AND2_X1   g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(G73), .A2(G543), .ZN(new_n602));
  INV_X1    g177(.A(G61), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n519), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n604), .A2(G651), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n601), .A2(new_n605), .ZN(G305));
  AOI22_X1  g181(.A1(new_n552), .A2(G85), .B1(G47), .B2(new_n538), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n536), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n585), .B2(new_n608), .ZN(G290));
  NAND2_X1  g184(.A1(G301), .A2(G868), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n552), .A2(KEYINPUT10), .A3(G92), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT10), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n536), .A2(new_n523), .ZN(new_n613));
  INV_X1    g188(.A(G92), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n612), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  AOI22_X1  g190(.A1(new_n611), .A2(new_n615), .B1(G54), .B2(new_n538), .ZN(new_n616));
  NAND2_X1  g191(.A1(G79), .A2(G543), .ZN(new_n617));
  INV_X1    g192(.A(G66), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n519), .B2(new_n618), .ZN(new_n619));
  OR2_X1    g194(.A1(new_n619), .A2(KEYINPUT80), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n619), .A2(KEYINPUT80), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n620), .A2(G651), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n616), .A2(new_n622), .ZN(new_n623));
  INV_X1    g198(.A(KEYINPUT81), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n623), .B(new_n624), .ZN(new_n625));
  INV_X1    g200(.A(new_n625), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n610), .B1(new_n626), .B2(G868), .ZN(G321));
  XOR2_X1   g202(.A(G321), .B(KEYINPUT82), .Z(G284));
  NOR2_X1   g203(.A1(G299), .A2(G868), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n629), .B1(G868), .B2(G168), .ZN(G297));
  XOR2_X1   g205(.A(G297), .B(KEYINPUT83), .Z(G280));
  INV_X1    g206(.A(G559), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n626), .B1(new_n632), .B2(G860), .ZN(G148));
  OAI21_X1  g208(.A(G868), .B1(new_n625), .B2(G559), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(G868), .B2(new_n574), .ZN(G323));
  XNOR2_X1  g210(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g211(.A1(new_n469), .A2(new_n467), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT12), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT84), .B(KEYINPUT13), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(KEYINPUT85), .B(G2100), .Z(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n489), .A2(G135), .ZN(new_n643));
  OAI21_X1  g218(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n644));
  INV_X1    g219(.A(G111), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n644), .B1(new_n645), .B2(G2105), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n646), .B1(G123), .B2(new_n493), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n643), .A2(new_n647), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n648), .A2(G2096), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n640), .A2(new_n641), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n648), .A2(G2096), .ZN(new_n651));
  NAND4_X1  g226(.A1(new_n642), .A2(new_n649), .A3(new_n650), .A4(new_n651), .ZN(G156));
  XNOR2_X1  g227(.A(KEYINPUT86), .B(KEYINPUT16), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT15), .B(G2435), .ZN(new_n655));
  INV_X1    g230(.A(G2438), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2427), .B(G2430), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  OAI21_X1  g234(.A(KEYINPUT14), .B1(new_n657), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n660), .A2(KEYINPUT87), .ZN(new_n661));
  INV_X1    g236(.A(KEYINPUT87), .ZN(new_n662));
  OAI211_X1 g237(.A(new_n662), .B(KEYINPUT14), .C1(new_n657), .C2(new_n659), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n657), .A2(new_n659), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1341), .B(G1348), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G2451), .B(G2454), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2443), .B(G2446), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n669), .B(new_n670), .Z(new_n671));
  INV_X1    g246(.A(new_n667), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n664), .A2(new_n665), .A3(new_n672), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n668), .A2(new_n671), .A3(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n671), .B1(new_n668), .B2(new_n673), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n654), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(new_n676), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n678), .A2(new_n674), .A3(new_n653), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n677), .A2(new_n679), .A3(G14), .ZN(new_n680));
  INV_X1    g255(.A(KEYINPUT88), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g257(.A1(new_n677), .A2(new_n679), .A3(KEYINPUT88), .A4(G14), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(G401));
  XOR2_X1   g260(.A(G2084), .B(G2090), .Z(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(G2072), .B(G2078), .Z(new_n688));
  XNOR2_X1  g263(.A(G2067), .B(G2678), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  NOR3_X1   g265(.A1(new_n687), .A2(new_n688), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT18), .ZN(new_n692));
  OR2_X1    g267(.A1(new_n688), .A2(KEYINPUT89), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n688), .A2(KEYINPUT89), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n693), .A2(new_n694), .A3(new_n690), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n688), .B(KEYINPUT17), .ZN(new_n696));
  OAI211_X1 g271(.A(new_n695), .B(new_n687), .C1(new_n696), .C2(new_n690), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n696), .A2(new_n690), .A3(new_n686), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n692), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(G2096), .B(G2100), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(G227));
  XOR2_X1   g276(.A(G1991), .B(G1996), .Z(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(G1971), .B(G1976), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT90), .B(KEYINPUT19), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(G1956), .B(G2474), .ZN(new_n709));
  XNOR2_X1  g284(.A(G1961), .B(G1966), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT20), .ZN(new_n713));
  INV_X1    g288(.A(new_n711), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n709), .A2(new_n710), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  MUX2_X1   g291(.A(new_n716), .B(new_n715), .S(new_n708), .Z(new_n717));
  NAND3_X1  g292(.A1(new_n713), .A2(KEYINPUT91), .A3(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  AOI21_X1  g294(.A(KEYINPUT91), .B1(new_n713), .B2(new_n717), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n705), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(new_n720), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n722), .A2(new_n718), .A3(new_n704), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n703), .B1(new_n721), .B2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  XNOR2_X1  g300(.A(G1981), .B(G1986), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n721), .A2(new_n723), .A3(new_n703), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n725), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(new_n726), .ZN(new_n729));
  INV_X1    g304(.A(new_n727), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n729), .B1(new_n730), .B2(new_n724), .ZN(new_n731));
  AND2_X1   g306(.A1(new_n728), .A2(new_n731), .ZN(G229));
  NOR2_X1   g307(.A1(G6), .A2(G16), .ZN(new_n733));
  INV_X1    g308(.A(G305), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n733), .B1(new_n734), .B2(G16), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT32), .ZN(new_n736));
  INV_X1    g311(.A(G1981), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  NOR2_X1   g313(.A1(G16), .A2(G22), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(G166), .B2(G16), .ZN(new_n740));
  INV_X1    g315(.A(G1971), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n742), .A2(KEYINPUT96), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n742), .A2(KEYINPUT96), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT95), .ZN(new_n745));
  NAND2_X1  g320(.A1(G288), .A2(new_n745), .ZN(new_n746));
  NAND4_X1  g321(.A1(new_n595), .A2(new_n596), .A3(KEYINPUT95), .A4(new_n597), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  MUX2_X1   g323(.A(G23), .B(new_n748), .S(G16), .Z(new_n749));
  XOR2_X1   g324(.A(KEYINPUT33), .B(G1976), .Z(new_n750));
  XOR2_X1   g325(.A(new_n749), .B(new_n750), .Z(new_n751));
  NAND4_X1  g326(.A1(new_n738), .A2(new_n743), .A3(new_n744), .A4(new_n751), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n752), .A2(KEYINPUT34), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(KEYINPUT34), .ZN(new_n754));
  NOR2_X1   g329(.A1(G16), .A2(G24), .ZN(new_n755));
  XOR2_X1   g330(.A(G290), .B(KEYINPUT94), .Z(new_n756));
  AOI21_X1  g331(.A(new_n755), .B1(new_n756), .B2(G16), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(G1986), .ZN(new_n758));
  INV_X1    g333(.A(G29), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n759), .A2(G25), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT92), .Z(new_n761));
  NAND2_X1  g336(.A1(new_n489), .A2(G131), .ZN(new_n762));
  OAI21_X1  g337(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n763));
  INV_X1    g338(.A(G107), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n763), .B1(new_n764), .B2(G2105), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(G119), .B2(new_n493), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n762), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT93), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n761), .B1(new_n768), .B2(G29), .ZN(new_n769));
  XOR2_X1   g344(.A(KEYINPUT35), .B(G1991), .Z(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n758), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n753), .A2(new_n754), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n773), .A2(KEYINPUT36), .ZN(new_n774));
  INV_X1    g349(.A(KEYINPUT36), .ZN(new_n775));
  NAND4_X1  g350(.A1(new_n753), .A2(new_n775), .A3(new_n754), .A4(new_n772), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(G16), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n778), .A2(G21), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G168), .B2(new_n778), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n780), .A2(G1966), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(KEYINPUT100), .Z(new_n782));
  NOR2_X1   g357(.A1(G171), .A2(new_n778), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(G5), .B2(new_n778), .ZN(new_n784));
  INV_X1    g359(.A(G1961), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  AND2_X1   g361(.A1(new_n780), .A2(G1966), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT99), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(new_n648), .B2(new_n759), .ZN(new_n789));
  NAND4_X1  g364(.A1(new_n643), .A2(KEYINPUT99), .A3(G29), .A4(new_n647), .ZN(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT30), .B(G28), .ZN(new_n791));
  OR2_X1    g366(.A1(KEYINPUT31), .A2(G11), .ZN(new_n792));
  NAND2_X1  g367(.A1(KEYINPUT31), .A2(G11), .ZN(new_n793));
  AOI22_X1  g368(.A1(new_n791), .A2(new_n759), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n789), .A2(new_n790), .A3(new_n794), .ZN(new_n795));
  NOR3_X1   g370(.A1(new_n786), .A2(new_n787), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n782), .A2(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(KEYINPUT101), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n782), .A2(new_n796), .A3(KEYINPUT101), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n759), .A2(G32), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n493), .A2(G129), .ZN(new_n802));
  INV_X1    g377(.A(KEYINPUT98), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NAND3_X1  g379(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT26), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n805), .A2(new_n806), .ZN(new_n808));
  AOI22_X1  g383(.A1(new_n807), .A2(new_n808), .B1(G105), .B2(new_n467), .ZN(new_n809));
  AND2_X1   g384(.A1(new_n804), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n489), .A2(G141), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(new_n812), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n801), .B1(new_n813), .B2(new_n759), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT27), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(G1996), .ZN(new_n816));
  INV_X1    g391(.A(G34), .ZN(new_n817));
  OR2_X1    g392(.A1(new_n817), .A2(KEYINPUT24), .ZN(new_n818));
  AOI21_X1  g393(.A(G29), .B1(new_n817), .B2(KEYINPUT24), .ZN(new_n819));
  AOI22_X1  g394(.A1(G160), .A2(G29), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n820), .A2(G2084), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(KEYINPUT102), .Z(new_n822));
  NAND2_X1  g397(.A1(new_n759), .A2(G33), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(KEYINPUT25), .Z(new_n825));
  AOI22_X1  g400(.A1(new_n469), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n825), .B1(new_n826), .B2(new_n465), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n827), .B1(new_n489), .B2(G139), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n823), .B1(new_n828), .B2(new_n759), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(new_n442), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n820), .A2(G2084), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n759), .A2(G27), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(G164), .B2(new_n759), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(new_n443), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n830), .A2(new_n831), .A3(new_n834), .ZN(new_n835));
  AOI211_X1 g410(.A(new_n822), .B(new_n835), .C1(new_n785), .C2(new_n784), .ZN(new_n836));
  NAND4_X1  g411(.A1(new_n799), .A2(new_n800), .A3(new_n816), .A4(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT103), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n837), .A2(new_n838), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n759), .A2(G35), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n841), .B1(G162), .B2(new_n759), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT29), .ZN(new_n843));
  OR2_X1    g418(.A1(new_n843), .A2(G2090), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n778), .A2(G20), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT23), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n846), .B1(new_n590), .B2(new_n778), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(G1956), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n848), .B1(new_n843), .B2(G2090), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n759), .A2(G26), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n850), .B(KEYINPUT28), .Z(new_n851));
  NAND2_X1  g426(.A1(new_n493), .A2(G128), .ZN(new_n852));
  XOR2_X1   g427(.A(new_n852), .B(KEYINPUT97), .Z(new_n853));
  NAND2_X1  g428(.A1(new_n489), .A2(G140), .ZN(new_n854));
  OR2_X1    g429(.A1(G104), .A2(G2105), .ZN(new_n855));
  OAI211_X1 g430(.A(new_n855), .B(G2104), .C1(G116), .C2(new_n465), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n853), .A2(new_n854), .A3(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n851), .B1(new_n857), .B2(G29), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(G2067), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n778), .A2(G19), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n860), .B1(new_n574), .B2(new_n778), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n861), .B(G1341), .Z(new_n862));
  NAND4_X1  g437(.A1(new_n844), .A2(new_n849), .A3(new_n859), .A4(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n778), .A2(G4), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n864), .B1(new_n626), .B2(new_n778), .ZN(new_n865));
  AND2_X1   g440(.A1(new_n865), .A2(G1348), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n865), .A2(G1348), .ZN(new_n867));
  NOR3_X1   g442(.A1(new_n863), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  NAND4_X1  g443(.A1(new_n777), .A2(new_n839), .A3(new_n840), .A4(new_n868), .ZN(G150));
  INV_X1    g444(.A(G150), .ZN(G311));
  NAND2_X1  g445(.A1(G80), .A2(G543), .ZN(new_n871));
  INV_X1    g446(.A(G67), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n871), .B1(new_n519), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(G651), .ZN(new_n874));
  XNOR2_X1  g449(.A(KEYINPUT105), .B(G93), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n536), .A2(new_n523), .A3(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT106), .ZN(new_n877));
  XOR2_X1   g452(.A(KEYINPUT104), .B(G55), .Z(new_n878));
  NAND2_X1  g453(.A1(new_n538), .A2(new_n878), .ZN(new_n879));
  AND3_X1   g454(.A1(new_n876), .A2(new_n877), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n877), .B1(new_n876), .B2(new_n879), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n874), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n882), .A2(new_n571), .A3(new_n572), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT107), .ZN(new_n884));
  OAI211_X1 g459(.A(new_n569), .B(new_n874), .C1(new_n880), .C2(new_n881), .ZN(new_n885));
  AND3_X1   g460(.A1(new_n883), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n884), .B1(new_n883), .B2(new_n885), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(KEYINPUT38), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n625), .A2(new_n632), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n889), .B(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT39), .ZN(new_n892));
  AOI21_X1  g467(.A(G860), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n893), .B1(new_n892), .B2(new_n891), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n882), .A2(G860), .ZN(new_n895));
  XOR2_X1   g470(.A(new_n895), .B(KEYINPUT37), .Z(new_n896));
  NAND2_X1  g471(.A1(new_n894), .A2(new_n896), .ZN(G145));
  OAI21_X1  g472(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n898));
  INV_X1    g473(.A(G118), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n898), .B1(new_n899), .B2(G2105), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n900), .B1(G130), .B2(new_n493), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n487), .A2(new_n488), .ZN(new_n902));
  INV_X1    g477(.A(G142), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n901), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(new_n638), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(new_n767), .ZN(new_n906));
  XOR2_X1   g481(.A(new_n906), .B(KEYINPUT109), .Z(new_n907));
  INV_X1    g482(.A(KEYINPUT108), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n509), .A2(new_n908), .ZN(new_n909));
  AOI22_X1  g484(.A1(new_n497), .A2(new_n502), .B1(new_n493), .B2(G126), .ZN(new_n910));
  NAND4_X1  g485(.A1(new_n910), .A2(KEYINPUT108), .A3(new_n506), .A4(new_n507), .ZN(new_n911));
  AND2_X1   g486(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n857), .B(new_n912), .ZN(new_n913));
  OR2_X1    g488(.A1(new_n913), .A2(new_n828), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n828), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n914), .A2(new_n813), .A3(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n813), .B1(new_n914), .B2(new_n915), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n907), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n914), .A2(new_n915), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(new_n812), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n906), .B(KEYINPUT109), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n921), .A2(new_n922), .A3(new_n916), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n919), .A2(new_n923), .ZN(new_n924));
  XOR2_X1   g499(.A(new_n648), .B(G160), .Z(new_n925));
  XNOR2_X1  g500(.A(new_n925), .B(G162), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(G37), .B1(new_n924), .B2(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n921), .A2(new_n916), .A3(new_n906), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n919), .A2(new_n929), .A3(new_n926), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n931), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g507(.A(KEYINPUT42), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n888), .A2(new_n626), .A3(new_n632), .ZN(new_n934));
  AND2_X1   g509(.A1(new_n616), .A2(new_n622), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(new_n590), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n623), .A2(G299), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT41), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n936), .A2(KEYINPUT41), .A3(new_n937), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  OAI22_X1  g517(.A1(new_n625), .A2(G559), .B1(new_n886), .B2(new_n887), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n934), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  AND2_X1   g519(.A1(new_n934), .A2(new_n943), .ZN(new_n945));
  INV_X1    g520(.A(new_n938), .ZN(new_n946));
  OAI211_X1 g521(.A(new_n933), .B(new_n944), .C1(new_n945), .C2(new_n946), .ZN(new_n947));
  AND3_X1   g522(.A1(new_n934), .A2(new_n942), .A3(new_n943), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n946), .B1(new_n934), .B2(new_n943), .ZN(new_n949));
  OAI21_X1  g524(.A(KEYINPUT42), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  XNOR2_X1  g525(.A(G166), .B(G290), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n748), .B(new_n734), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n951), .B(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  AND3_X1   g529(.A1(new_n947), .A2(new_n950), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n954), .B1(new_n947), .B2(new_n950), .ZN(new_n956));
  OAI21_X1  g531(.A(G868), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT110), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n876), .A2(new_n879), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(KEYINPUT106), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n876), .A2(new_n877), .A3(new_n879), .ZN(new_n961));
  AOI22_X1  g536(.A1(new_n960), .A2(new_n961), .B1(G651), .B2(new_n873), .ZN(new_n962));
  OR2_X1    g537(.A1(new_n962), .A2(G868), .ZN(new_n963));
  AND3_X1   g538(.A1(new_n957), .A2(new_n958), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n958), .B1(new_n957), .B2(new_n963), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n964), .A2(new_n965), .ZN(G295));
  NAND2_X1  g541(.A1(new_n957), .A2(new_n963), .ZN(G331));
  XNOR2_X1  g542(.A(G168), .B(G171), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n968), .B1(new_n886), .B2(new_n887), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n885), .B1(new_n573), .B2(new_n962), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(KEYINPUT107), .ZN(new_n971));
  XNOR2_X1  g546(.A(G168), .B(G301), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n883), .A2(new_n884), .A3(new_n885), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n971), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n969), .A2(new_n974), .A3(new_n946), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n972), .B1(new_n971), .B2(new_n973), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n974), .A2(KEYINPUT111), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT111), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n971), .A2(new_n972), .A3(new_n978), .A4(new_n973), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n976), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n975), .B1(new_n980), .B2(new_n942), .ZN(new_n981));
  AOI21_X1  g556(.A(G37), .B1(new_n981), .B2(new_n954), .ZN(new_n982));
  OAI211_X1 g557(.A(new_n953), .B(new_n975), .C1(new_n980), .C2(new_n942), .ZN(new_n983));
  AOI21_X1  g558(.A(KEYINPUT43), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n969), .A2(new_n946), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n985), .B1(new_n977), .B2(new_n979), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n942), .B1(new_n969), .B2(new_n974), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n954), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(G37), .ZN(new_n989));
  AND4_X1   g564(.A1(KEYINPUT43), .A2(new_n988), .A3(new_n989), .A4(new_n983), .ZN(new_n990));
  OAI21_X1  g565(.A(KEYINPUT44), .B1(new_n984), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n981), .A2(new_n954), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n992), .A2(new_n989), .A3(new_n983), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(KEYINPUT43), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT43), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n988), .A2(new_n983), .A3(new_n995), .A4(new_n989), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n991), .B1(new_n998), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g574(.A(G1384), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n909), .A2(new_n911), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT45), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(G160), .A2(G40), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(G1996), .ZN(new_n1006));
  XNOR2_X1  g581(.A(new_n812), .B(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(G2067), .ZN(new_n1008));
  XNOR2_X1  g583(.A(new_n857), .B(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  XOR2_X1   g585(.A(new_n767), .B(new_n770), .Z(new_n1011));
  OAI21_X1  g586(.A(new_n1005), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g587(.A1(G290), .A2(G1986), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1005), .A2(new_n1013), .A3(KEYINPUT48), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1005), .A2(new_n1013), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT48), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  AND3_X1   g592(.A1(new_n1012), .A2(new_n1014), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1009), .A2(new_n813), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT46), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1021));
  AOI22_X1  g596(.A1(new_n1019), .A2(new_n1005), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1021), .A2(new_n1020), .ZN(new_n1023));
  AND2_X1   g598(.A1(new_n1023), .A2(KEYINPUT126), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1023), .A2(KEYINPUT126), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1022), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  XOR2_X1   g601(.A(new_n1026), .B(KEYINPUT47), .Z(new_n1027));
  INV_X1    g602(.A(new_n768), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(new_n770), .ZN(new_n1029));
  OAI22_X1  g604(.A1(new_n1010), .A2(new_n1029), .B1(G2067), .B2(new_n857), .ZN(new_n1030));
  AOI211_X1 g605(.A(new_n1018), .B(new_n1027), .C1(new_n1005), .C2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n746), .A2(G1976), .A3(new_n747), .ZN(new_n1032));
  INV_X1    g607(.A(G8), .ZN(new_n1033));
  INV_X1    g608(.A(G40), .ZN(new_n1034));
  AOI211_X1 g609(.A(new_n1034), .B(new_n472), .C1(new_n481), .C2(G2105), .ZN(new_n1035));
  AND2_X1   g610(.A1(new_n509), .A2(new_n1000), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1033), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1032), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(KEYINPUT52), .ZN(new_n1039));
  INV_X1    g614(.A(G1976), .ZN(new_n1040));
  AOI21_X1  g615(.A(KEYINPUT52), .B1(G288), .B2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1032), .A2(new_n1037), .A3(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT117), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n601), .A2(new_n737), .A3(new_n605), .ZN(new_n1044));
  AND2_X1   g619(.A1(new_n604), .A2(G651), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n599), .A2(new_n600), .ZN(new_n1046));
  OAI21_X1  g621(.A(G1981), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1043), .B1(new_n1044), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT49), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1037), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  AOI211_X1 g625(.A(new_n1043), .B(KEYINPUT49), .C1(new_n1044), .C2(new_n1047), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1039), .B(new_n1042), .C1(new_n1050), .C2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n531), .A2(G8), .A3(new_n533), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT114), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(KEYINPUT55), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT50), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n509), .A2(new_n1058), .A3(new_n1000), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT113), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n509), .A2(new_n1000), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(KEYINPUT50), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1004), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(G2090), .ZN(new_n1065));
  AOI211_X1 g640(.A(KEYINPUT113), .B(new_n1058), .C1(new_n509), .C2(new_n1000), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1064), .A2(new_n1065), .A3(new_n1067), .ZN(new_n1068));
  XOR2_X1   g643(.A(KEYINPUT114), .B(KEYINPUT55), .Z(new_n1069));
  NAND4_X1  g644(.A1(new_n531), .A2(G8), .A3(new_n533), .A4(new_n1069), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n909), .A2(new_n911), .A3(KEYINPUT45), .A4(new_n1000), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1062), .A2(new_n1002), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1035), .A2(new_n1073), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n741), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1057), .A2(new_n1068), .A3(new_n1070), .A4(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(G2084), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1064), .A2(new_n1077), .A3(new_n1067), .ZN(new_n1078));
  INV_X1    g653(.A(G1966), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1062), .A2(new_n1002), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1079), .B1(new_n1074), .B2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1033), .B1(new_n1078), .B2(new_n1081), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1053), .A2(G168), .A3(new_n1076), .A4(new_n1082), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1084));
  OR2_X1    g659(.A1(G288), .A2(G1976), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1044), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  AOI22_X1  g661(.A1(new_n1083), .A2(KEYINPUT63), .B1(new_n1037), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT63), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1082), .A2(new_n1088), .A3(G168), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1057), .A2(new_n1070), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1075), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1058), .B1(new_n509), .B2(new_n1000), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT118), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1059), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n509), .A2(KEYINPUT118), .A3(new_n1058), .A4(new_n1000), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1095), .A2(new_n1035), .A3(new_n1096), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1097), .A2(G2090), .ZN(new_n1098));
  OAI21_X1  g673(.A(G8), .B1(new_n1092), .B2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1089), .B1(new_n1091), .B2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1033), .B1(new_n1068), .B2(new_n1075), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT115), .ZN(new_n1102));
  AND3_X1   g677(.A1(new_n1057), .A2(new_n1102), .A3(new_n1070), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1102), .B1(new_n1057), .B2(new_n1070), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1101), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(KEYINPUT116), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT116), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1107), .B(new_n1101), .C1(new_n1103), .C2(new_n1104), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1100), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1087), .B1(new_n1109), .B2(new_n1052), .ZN(new_n1110));
  INV_X1    g685(.A(G1956), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1097), .A2(new_n1111), .ZN(new_n1112));
  XNOR2_X1  g687(.A(KEYINPUT56), .B(G2072), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1071), .A2(new_n1035), .A3(new_n1073), .A4(new_n1113), .ZN(new_n1114));
  AND2_X1   g689(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n581), .A2(KEYINPUT9), .ZN(new_n1116));
  OR2_X1    g691(.A1(new_n581), .A2(KEYINPUT9), .ZN(new_n1117));
  AOI22_X1  g692(.A1(new_n552), .A2(G91), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n586), .A2(new_n588), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(G651), .ZN(new_n1120));
  OR2_X1    g695(.A1(KEYINPUT119), .A2(KEYINPUT57), .ZN(new_n1121));
  NAND2_X1  g696(.A1(KEYINPUT119), .A2(KEYINPUT57), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1118), .A2(new_n1120), .A3(new_n1121), .A4(new_n1122), .ZN(new_n1123));
  OAI211_X1 g698(.A(KEYINPUT119), .B(KEYINPUT57), .C1(new_n584), .C2(new_n589), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT120), .ZN(new_n1125));
  AND3_X1   g700(.A1(new_n1123), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1125), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1115), .A2(new_n1128), .ZN(new_n1129));
  AND2_X1   g704(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1112), .A2(new_n1114), .A3(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(G1348), .B1(new_n1064), .B2(new_n1067), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1004), .A2(new_n1062), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(new_n1008), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1134), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1132), .A2(new_n1135), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1136), .A2(new_n623), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1129), .B1(new_n1131), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT61), .ZN(new_n1139));
  AND3_X1   g714(.A1(new_n1112), .A2(new_n1114), .A3(new_n1130), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1130), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1139), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1136), .A2(KEYINPUT60), .A3(new_n623), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1071), .A2(new_n1035), .A3(new_n1006), .A4(new_n1073), .ZN(new_n1144));
  XNOR2_X1  g719(.A(KEYINPUT58), .B(G1341), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1144), .B1(new_n1133), .B2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(new_n574), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1147), .A2(KEYINPUT59), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT59), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1146), .A2(new_n1149), .A3(new_n574), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1142), .A2(new_n1143), .A3(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT60), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1153), .B1(new_n1132), .B2(new_n1135), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1093), .B1(new_n1060), .B2(new_n1059), .ZN(new_n1155));
  NOR3_X1   g730(.A1(new_n1155), .A2(new_n1004), .A3(new_n1066), .ZN(new_n1156));
  OAI211_X1 g731(.A(KEYINPUT60), .B(new_n1134), .C1(new_n1156), .C2(G1348), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1154), .A2(new_n1157), .A3(new_n935), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1131), .A2(KEYINPUT61), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1158), .B1(new_n1129), .B2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1138), .B1(new_n1152), .B2(new_n1160), .ZN(new_n1161));
  OR2_X1    g736(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1162));
  AND2_X1   g737(.A1(new_n1039), .A2(new_n1042), .ZN(new_n1163));
  OR2_X1    g738(.A1(new_n1097), .A2(G2090), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1033), .B1(new_n1164), .B2(new_n1075), .ZN(new_n1165));
  OAI211_X1 g740(.A(new_n1162), .B(new_n1163), .C1(new_n1165), .C2(new_n1090), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1166), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1071), .A2(new_n1035), .A3(new_n443), .A4(new_n1073), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT53), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1169), .A2(G2078), .ZN(new_n1171));
  NAND4_X1  g746(.A1(new_n1003), .A2(new_n1035), .A3(new_n1071), .A4(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1170), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1173), .ZN(new_n1174));
  NOR3_X1   g749(.A1(new_n1156), .A2(KEYINPUT121), .A3(G1961), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT121), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1064), .A2(new_n1067), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1176), .B1(new_n1177), .B2(new_n785), .ZN(new_n1178));
  OAI211_X1 g753(.A(new_n1174), .B(G301), .C1(new_n1175), .C2(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(new_n1171), .ZN(new_n1180));
  OR3_X1    g755(.A1(new_n1074), .A2(new_n1080), .A3(new_n1180), .ZN(new_n1181));
  OAI211_X1 g756(.A(new_n1181), .B(new_n1170), .C1(G1961), .C2(new_n1156), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1182), .A2(G171), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1179), .A2(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT54), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1078), .A2(new_n1081), .ZN(new_n1186));
  OAI21_X1  g761(.A(G8), .B1(new_n1186), .B2(G286), .ZN(new_n1187));
  AOI21_X1  g762(.A(G168), .B1(new_n1078), .B2(new_n1081), .ZN(new_n1188));
  OAI21_X1  g763(.A(KEYINPUT51), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT51), .ZN(new_n1190));
  OAI211_X1 g765(.A(new_n1190), .B(G8), .C1(new_n1186), .C2(G286), .ZN(new_n1191));
  AOI22_X1  g766(.A1(new_n1184), .A2(new_n1185), .B1(new_n1189), .B2(new_n1191), .ZN(new_n1192));
  AND3_X1   g767(.A1(new_n1161), .A2(new_n1167), .A3(new_n1192), .ZN(new_n1193));
  NOR2_X1   g768(.A1(new_n1182), .A2(G171), .ZN(new_n1194));
  NOR2_X1   g769(.A1(new_n1194), .A2(new_n1185), .ZN(new_n1195));
  OAI21_X1  g770(.A(KEYINPUT121), .B1(new_n1156), .B2(G1961), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1177), .A2(new_n1176), .A3(new_n785), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n1173), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  INV_X1    g773(.A(KEYINPUT122), .ZN(new_n1199));
  OAI21_X1  g774(.A(G171), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  OAI211_X1 g775(.A(new_n1174), .B(new_n1199), .C1(new_n1175), .C2(new_n1178), .ZN(new_n1201));
  INV_X1    g776(.A(new_n1201), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n1195), .B1(new_n1200), .B2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1203), .A2(KEYINPUT123), .ZN(new_n1204));
  INV_X1    g779(.A(KEYINPUT123), .ZN(new_n1205));
  OAI211_X1 g780(.A(new_n1195), .B(new_n1205), .C1(new_n1200), .C2(new_n1202), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1204), .A2(new_n1206), .ZN(new_n1207));
  AOI21_X1  g782(.A(new_n1110), .B1(new_n1193), .B2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1209));
  INV_X1    g784(.A(KEYINPUT62), .ZN(new_n1210));
  NAND3_X1  g785(.A1(new_n1189), .A2(new_n1210), .A3(new_n1191), .ZN(new_n1211));
  INV_X1    g786(.A(new_n1166), .ZN(new_n1212));
  INV_X1    g787(.A(new_n1183), .ZN(new_n1213));
  NAND4_X1  g788(.A1(new_n1209), .A2(new_n1211), .A3(new_n1212), .A4(new_n1213), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1214), .A2(KEYINPUT124), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1189), .A2(new_n1191), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n1216), .A2(KEYINPUT62), .ZN(new_n1217));
  INV_X1    g792(.A(KEYINPUT124), .ZN(new_n1218));
  NAND4_X1  g793(.A1(new_n1167), .A2(new_n1218), .A3(new_n1211), .A4(new_n1213), .ZN(new_n1219));
  NAND3_X1  g794(.A1(new_n1215), .A2(new_n1217), .A3(new_n1219), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n1208), .A2(new_n1220), .ZN(new_n1221));
  NAND3_X1  g796(.A1(new_n1005), .A2(G1986), .A3(G290), .ZN(new_n1222));
  NAND2_X1  g797(.A1(new_n1222), .A2(new_n1015), .ZN(new_n1223));
  XOR2_X1   g798(.A(new_n1223), .B(KEYINPUT112), .Z(new_n1224));
  NAND2_X1  g799(.A1(new_n1224), .A2(new_n1012), .ZN(new_n1225));
  INV_X1    g800(.A(new_n1225), .ZN(new_n1226));
  AOI21_X1  g801(.A(KEYINPUT125), .B1(new_n1221), .B2(new_n1226), .ZN(new_n1227));
  INV_X1    g802(.A(KEYINPUT125), .ZN(new_n1228));
  AOI211_X1 g803(.A(new_n1228), .B(new_n1225), .C1(new_n1208), .C2(new_n1220), .ZN(new_n1229));
  OAI21_X1  g804(.A(new_n1031), .B1(new_n1227), .B2(new_n1229), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g805(.A(KEYINPUT127), .ZN(new_n1232));
  NAND2_X1  g806(.A1(new_n728), .A2(new_n731), .ZN(new_n1233));
  NOR2_X1   g807(.A1(G227), .A2(new_n463), .ZN(new_n1234));
  NAND3_X1  g808(.A1(new_n684), .A2(new_n1233), .A3(new_n1234), .ZN(new_n1235));
  AOI21_X1  g809(.A(new_n1235), .B1(new_n928), .B2(new_n930), .ZN(new_n1236));
  AOI21_X1  g810(.A(new_n1232), .B1(new_n997), .B2(new_n1236), .ZN(new_n1237));
  AOI21_X1  g811(.A(new_n995), .B1(new_n982), .B2(new_n983), .ZN(new_n1238));
  INV_X1    g812(.A(new_n996), .ZN(new_n1239));
  OAI211_X1 g813(.A(new_n1236), .B(new_n1232), .C1(new_n1238), .C2(new_n1239), .ZN(new_n1240));
  INV_X1    g814(.A(new_n1240), .ZN(new_n1241));
  NOR2_X1   g815(.A1(new_n1237), .A2(new_n1241), .ZN(G308));
  NAND2_X1  g816(.A1(new_n997), .A2(new_n1236), .ZN(G225));
endmodule


