//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 0 0 0 1 0 0 1 1 0 0 0 1 1 0 0 0 1 0 1 1 0 1 1 0 1 0 0 0 1 1 1 0 0 1 0 0 1 0 1 0 0 0 0 1 1 1 0 1 1 0 1 1 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n779,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n955, new_n956, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n971, new_n972, new_n973, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1007, new_n1008;
  XNOR2_X1  g000(.A(G197gat), .B(G204gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G211gat), .B(G218gat), .ZN(new_n203));
  INV_X1    g002(.A(G218gat), .ZN(new_n204));
  INV_X1    g003(.A(G211gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(KEYINPUT68), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT68), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(G211gat), .ZN(new_n208));
  AOI21_X1  g007(.A(new_n204), .B1(new_n206), .B2(new_n208), .ZN(new_n209));
  OAI211_X1 g008(.A(new_n202), .B(new_n203), .C1(new_n209), .C2(KEYINPUT22), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT22), .ZN(new_n212));
  XNOR2_X1  g011(.A(KEYINPUT68), .B(G211gat), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n212), .B1(new_n213), .B2(new_n204), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n203), .B1(new_n214), .B2(new_n202), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n211), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(G226gat), .ZN(new_n217));
  INV_X1    g016(.A(G233gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(G169gat), .ZN(new_n221));
  INV_X1    g020(.A(G176gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n221), .A2(new_n222), .A3(KEYINPUT26), .ZN(new_n223));
  NAND2_X1  g022(.A1(G183gat), .A2(G190gat), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT26), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n225), .B1(G169gat), .B2(G176gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(G169gat), .A2(G176gat), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  OAI211_X1 g027(.A(new_n223), .B(new_n224), .C1(new_n226), .C2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(G183gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(KEYINPUT27), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT27), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(G183gat), .ZN(new_n233));
  INV_X1    g032(.A(G190gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n231), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT28), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(KEYINPUT27), .B(G183gat), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n238), .A2(KEYINPUT28), .A3(new_n234), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n229), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT23), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n241), .B1(G169gat), .B2(G176gat), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n234), .A2(KEYINPUT24), .A3(G183gat), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n242), .A2(new_n243), .A3(new_n227), .ZN(new_n244));
  NAND2_X1  g043(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(G190gat), .ZN(new_n246));
  NOR2_X1   g045(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n244), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n221), .A2(new_n222), .A3(KEYINPUT23), .ZN(new_n250));
  OAI211_X1 g049(.A(new_n249), .B(new_n250), .C1(KEYINPUT64), .C2(KEYINPUT25), .ZN(new_n251));
  AND2_X1   g050(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n252));
  AOI22_X1  g051(.A1(new_n252), .A2(new_n234), .B1(G169gat), .B2(G176gat), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT24), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(new_n230), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n255), .A2(G190gat), .A3(new_n245), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n253), .A2(new_n256), .A3(KEYINPUT64), .A4(new_n242), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n253), .A2(new_n256), .A3(new_n242), .A4(new_n250), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT25), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n257), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n240), .B1(new_n251), .B2(new_n260), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n220), .B1(new_n261), .B2(KEYINPUT29), .ZN(new_n262));
  INV_X1    g061(.A(new_n240), .ZN(new_n263));
  AND3_X1   g062(.A1(new_n257), .A2(new_n258), .A3(new_n259), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n258), .B1(new_n259), .B2(new_n257), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n263), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(new_n219), .ZN(new_n267));
  AOI21_X1  g066(.A(KEYINPUT69), .B1(new_n262), .B2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT69), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT29), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n266), .A2(new_n270), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n269), .B1(new_n271), .B2(new_n220), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n216), .B1(new_n268), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(KEYINPUT70), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT70), .ZN(new_n276));
  OAI211_X1 g075(.A(new_n276), .B(new_n216), .C1(new_n268), .C2(new_n272), .ZN(new_n277));
  AND2_X1   g076(.A1(new_n262), .A2(new_n267), .ZN(new_n278));
  INV_X1    g077(.A(new_n203), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n206), .A2(new_n208), .ZN(new_n280));
  AOI21_X1  g079(.A(KEYINPUT22), .B1(new_n280), .B2(G218gat), .ZN(new_n281));
  INV_X1    g080(.A(new_n202), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n279), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(new_n210), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n278), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n277), .A2(new_n285), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n275), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT37), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(G8gat), .B(G36gat), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n290), .B(KEYINPUT71), .ZN(new_n291));
  XNOR2_X1  g090(.A(G64gat), .B(G92gat), .ZN(new_n292));
  XOR2_X1   g091(.A(new_n291), .B(new_n292), .Z(new_n293));
  NAND2_X1  g092(.A1(new_n289), .A2(new_n293), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n287), .A2(new_n288), .ZN(new_n295));
  OAI21_X1  g094(.A(KEYINPUT38), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  OR3_X1    g095(.A1(new_n268), .A2(new_n272), .A3(new_n216), .ZN(new_n297));
  OR2_X1    g096(.A1(new_n297), .A2(KEYINPUT82), .ZN(new_n298));
  OR2_X1    g097(.A1(new_n278), .A2(new_n284), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n297), .A2(KEYINPUT82), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(KEYINPUT37), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT38), .ZN(new_n303));
  NAND4_X1  g102(.A1(new_n302), .A2(new_n303), .A3(new_n293), .A4(new_n289), .ZN(new_n304));
  INV_X1    g103(.A(G120gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(G113gat), .ZN(new_n306));
  INV_X1    g105(.A(G113gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(G120gat), .ZN(new_n308));
  AND3_X1   g107(.A1(new_n306), .A2(new_n308), .A3(KEYINPUT65), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT65), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n310), .A2(new_n307), .A3(G120gat), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT1), .ZN(new_n312));
  INV_X1    g111(.A(G134gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(G127gat), .ZN(new_n314));
  INV_X1    g113(.A(G127gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(G134gat), .ZN(new_n316));
  NAND4_X1  g115(.A1(new_n311), .A2(new_n312), .A3(new_n314), .A4(new_n316), .ZN(new_n317));
  AOI21_X1  g116(.A(KEYINPUT1), .B1(new_n306), .B2(new_n308), .ZN(new_n318));
  AND2_X1   g117(.A1(new_n314), .A2(new_n316), .ZN(new_n319));
  OAI22_X1  g118(.A1(new_n309), .A2(new_n317), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  AND2_X1   g119(.A1(G155gat), .A2(G162gat), .ZN(new_n321));
  NOR2_X1   g120(.A1(G155gat), .A2(G162gat), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(G141gat), .B(G148gat), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT2), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n325), .B1(G155gat), .B2(G162gat), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n323), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(G141gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(G148gat), .ZN(new_n329));
  INV_X1    g128(.A(G148gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(G141gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(G155gat), .B(G162gat), .ZN(new_n333));
  INV_X1    g132(.A(G155gat), .ZN(new_n334));
  INV_X1    g133(.A(G162gat), .ZN(new_n335));
  OAI21_X1  g134(.A(KEYINPUT2), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n332), .A2(new_n333), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n327), .A2(new_n337), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n320), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT4), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n338), .A2(KEYINPUT3), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT3), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n327), .A2(new_n337), .A3(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n342), .A2(new_n344), .A3(new_n320), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n341), .A2(new_n345), .ZN(new_n346));
  NOR3_X1   g145(.A1(new_n320), .A2(new_n338), .A3(KEYINPUT4), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(G225gat), .A2(G233gat), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT5), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n351), .A2(KEYINPUT73), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n349), .A2(new_n350), .A3(new_n352), .ZN(new_n353));
  AND2_X1   g152(.A1(new_n327), .A2(new_n337), .ZN(new_n354));
  OR2_X1    g153(.A1(new_n318), .A2(new_n319), .ZN(new_n355));
  OR2_X1    g154(.A1(new_n309), .A2(new_n317), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n320), .A2(new_n338), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n350), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n351), .B1(new_n359), .B2(KEYINPUT74), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT74), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n354), .B(new_n320), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n361), .B1(new_n362), .B2(new_n350), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n360), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n352), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n347), .B1(new_n341), .B2(new_n345), .ZN(new_n366));
  INV_X1    g165(.A(new_n350), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n365), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  XNOR2_X1  g167(.A(G1gat), .B(G29gat), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n369), .B(KEYINPUT0), .ZN(new_n370));
  XNOR2_X1  g169(.A(G57gat), .B(G85gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n370), .B(new_n371), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n353), .A2(new_n364), .A3(new_n368), .A4(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(KEYINPUT81), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n353), .A2(new_n364), .A3(new_n368), .ZN(new_n376));
  INV_X1    g175(.A(new_n372), .ZN(new_n377));
  AOI21_X1  g176(.A(KEYINPUT6), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT81), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n373), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n375), .A2(new_n378), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n374), .A2(KEYINPUT6), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n293), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n383), .B1(new_n287), .B2(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n296), .A2(new_n304), .A3(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(KEYINPUT3), .B1(new_n284), .B2(new_n270), .ZN(new_n387));
  AND2_X1   g186(.A1(new_n344), .A2(new_n270), .ZN(new_n388));
  OAI22_X1  g187(.A1(new_n387), .A2(new_n354), .B1(new_n284), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n344), .A2(new_n270), .ZN(new_n390));
  AOI21_X1  g189(.A(KEYINPUT75), .B1(new_n216), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(G228gat), .A2(G233gat), .ZN(new_n392));
  NOR3_X1   g191(.A1(new_n391), .A2(G22gat), .A3(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(G22gat), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT75), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n395), .B1(new_n388), .B2(new_n284), .ZN(new_n396));
  INV_X1    g195(.A(new_n392), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n394), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n389), .B1(new_n393), .B2(new_n398), .ZN(new_n399));
  XNOR2_X1  g198(.A(G78gat), .B(G106gat), .ZN(new_n400));
  XNOR2_X1  g199(.A(KEYINPUT31), .B(G50gat), .ZN(new_n401));
  XOR2_X1   g200(.A(new_n400), .B(new_n401), .Z(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n343), .B1(new_n216), .B2(KEYINPUT29), .ZN(new_n404));
  AOI22_X1  g203(.A1(new_n404), .A2(new_n338), .B1(new_n216), .B2(new_n390), .ZN(new_n405));
  OAI21_X1  g204(.A(G22gat), .B1(new_n391), .B2(new_n392), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n396), .A2(new_n394), .A3(new_n397), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n405), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n399), .A2(new_n403), .A3(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT77), .ZN(new_n410));
  AND2_X1   g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n409), .A2(new_n410), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT76), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n399), .A2(new_n408), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n413), .B1(new_n414), .B2(new_n402), .ZN(new_n415));
  AOI211_X1 g214(.A(KEYINPUT76), .B(new_n403), .C1(new_n399), .C2(new_n408), .ZN(new_n416));
  OAI22_X1  g215(.A1(new_n411), .A2(new_n412), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(KEYINPUT79), .B1(new_n349), .B2(new_n350), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT79), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n366), .A2(new_n420), .A3(new_n367), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT39), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n372), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n423), .B1(new_n362), .B2(new_n350), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n424), .B1(new_n422), .B2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT40), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n427), .A2(KEYINPUT80), .A3(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT80), .ZN(new_n430));
  OAI221_X1 g229(.A(new_n424), .B1(new_n430), .B2(KEYINPUT40), .C1(new_n422), .C2(new_n426), .ZN(new_n431));
  AND2_X1   g230(.A1(new_n375), .A2(new_n380), .ZN(new_n432));
  AND3_X1   g231(.A1(new_n429), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n274), .A2(new_n285), .A3(new_n277), .A4(new_n384), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT30), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AND2_X1   g235(.A1(new_n277), .A2(new_n285), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n293), .B1(new_n437), .B2(new_n274), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n384), .A2(KEYINPUT30), .ZN(new_n439));
  AND4_X1   g238(.A1(new_n274), .A2(new_n285), .A3(new_n277), .A4(new_n439), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n436), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n418), .B1(new_n433), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n378), .A2(new_n373), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(new_n382), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n436), .A2(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(KEYINPUT72), .B1(new_n438), .B2(new_n440), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n384), .B1(new_n275), .B2(new_n286), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n437), .A2(new_n274), .A3(new_n439), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT72), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n445), .B1(new_n446), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  XNOR2_X1  g251(.A(new_n417), .B(KEYINPUT78), .ZN(new_n453));
  AOI22_X1  g252(.A1(new_n386), .A2(new_n442), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(G227gat), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n455), .A2(new_n218), .ZN(new_n456));
  INV_X1    g255(.A(new_n320), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n251), .A2(new_n260), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n457), .B1(new_n458), .B2(new_n263), .ZN(new_n459));
  AOI211_X1 g258(.A(new_n320), .B(new_n240), .C1(new_n251), .C2(new_n260), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n456), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT33), .ZN(new_n462));
  XNOR2_X1  g261(.A(G15gat), .B(G43gat), .ZN(new_n463));
  XNOR2_X1  g262(.A(G71gat), .B(G99gat), .ZN(new_n464));
  XNOR2_X1  g263(.A(new_n463), .B(new_n464), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n461), .B(KEYINPUT32), .C1(new_n462), .C2(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n465), .B1(new_n461), .B2(KEYINPUT32), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT66), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n461), .A2(new_n462), .ZN(new_n469));
  AND3_X1   g268(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n468), .B1(new_n467), .B2(new_n469), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n466), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT34), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n459), .A2(new_n460), .ZN(new_n474));
  INV_X1    g273(.A(new_n456), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NOR4_X1   g275(.A1(new_n459), .A2(new_n460), .A3(KEYINPUT34), .A4(new_n456), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n472), .A2(new_n479), .ZN(new_n480));
  OAI211_X1 g279(.A(new_n478), .B(new_n466), .C1(new_n470), .C2(new_n471), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n480), .A2(KEYINPUT36), .A3(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(new_n466), .ZN(new_n483));
  INV_X1    g282(.A(new_n471), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(KEYINPUT67), .B1(new_n486), .B2(new_n478), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n480), .A2(new_n481), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n487), .B1(new_n488), .B2(KEYINPUT67), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n482), .B1(new_n489), .B2(KEYINPUT36), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n417), .A2(new_n480), .A3(new_n481), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT83), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n417), .A2(new_n480), .A3(KEYINPUT83), .A4(new_n481), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n451), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(KEYINPUT35), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT35), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n383), .A2(new_n417), .A3(new_n497), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n498), .A2(new_n441), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(new_n489), .ZN(new_n500));
  AOI22_X1  g299(.A1(new_n454), .A2(new_n490), .B1(new_n496), .B2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(G50gat), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(G43gat), .ZN(new_n503));
  INV_X1    g302(.A(G43gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(G50gat), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT85), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n503), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(KEYINPUT15), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n506), .B1(new_n503), .B2(new_n505), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(G29gat), .ZN(new_n511));
  INV_X1    g310(.A(G36gat), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n511), .A2(new_n512), .A3(KEYINPUT14), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT14), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n515), .B1(G29gat), .B2(G36gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n510), .B1(new_n513), .B2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT15), .ZN(new_n519));
  OR2_X1    g318(.A1(KEYINPUT88), .A2(G50gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(KEYINPUT88), .A2(G50gat), .ZN(new_n521));
  AOI21_X1  g320(.A(G43gat), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT87), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n523), .B1(new_n504), .B2(G50gat), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n502), .A2(KEYINPUT87), .A3(G43gat), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n519), .B1(new_n522), .B2(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(KEYINPUT89), .B1(new_n514), .B2(new_n516), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n528), .A2(new_n513), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT89), .ZN(new_n530));
  OAI211_X1 g329(.A(new_n527), .B(new_n529), .C1(new_n530), .C2(new_n517), .ZN(new_n531));
  OAI21_X1  g330(.A(KEYINPUT86), .B1(new_n508), .B2(new_n509), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n503), .A2(new_n505), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(KEYINPUT85), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT86), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n534), .A2(new_n535), .A3(KEYINPUT15), .A4(new_n507), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n532), .A2(new_n536), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n518), .B1(new_n531), .B2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(G8gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(G15gat), .B(G22gat), .ZN(new_n540));
  INV_X1    g339(.A(G1gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(KEYINPUT16), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT90), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n539), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n543), .B1(G1gat), .B2(new_n540), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  OAI221_X1 g346(.A(new_n543), .B1(new_n544), .B2(new_n539), .C1(G1gat), .C2(new_n540), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n538), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n549), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n517), .A2(new_n530), .ZN(new_n552));
  NOR3_X1   g351(.A1(new_n552), .A2(new_n513), .A3(new_n528), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n553), .A2(new_n527), .A3(new_n536), .A4(new_n532), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n551), .A2(new_n518), .A3(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n550), .A2(new_n555), .A3(KEYINPUT91), .ZN(new_n556));
  NAND2_X1  g355(.A1(G229gat), .A2(G233gat), .ZN(new_n557));
  XOR2_X1   g356(.A(new_n557), .B(KEYINPUT13), .Z(new_n558));
  INV_X1    g357(.A(KEYINPUT91), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n538), .A2(new_n559), .A3(new_n549), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n556), .A2(new_n558), .A3(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT92), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n556), .A2(KEYINPUT92), .A3(new_n558), .A4(new_n560), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT17), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n538), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n554), .A2(KEYINPUT17), .A3(new_n518), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n567), .A2(new_n551), .A3(new_n568), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n569), .A2(new_n557), .A3(new_n550), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT18), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT93), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n569), .A2(KEYINPUT18), .A3(new_n557), .A4(new_n550), .ZN(new_n575));
  XNOR2_X1  g374(.A(G113gat), .B(G141gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(G169gat), .B(G197gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n580), .B(KEYINPUT12), .ZN(new_n581));
  AND2_X1   g380(.A1(new_n575), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n570), .A2(KEYINPUT93), .A3(new_n571), .ZN(new_n583));
  AND4_X1   g382(.A1(new_n565), .A2(new_n574), .A3(new_n582), .A4(new_n583), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n549), .B1(new_n538), .B2(new_n566), .ZN(new_n585));
  AOI22_X1  g384(.A1(new_n585), .A2(new_n568), .B1(new_n549), .B2(new_n538), .ZN(new_n586));
  AOI21_X1  g385(.A(KEYINPUT18), .B1(new_n586), .B2(new_n557), .ZN(new_n587));
  INV_X1    g386(.A(new_n575), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n581), .B1(new_n589), .B2(new_n565), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n584), .A2(new_n590), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n501), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(G134gat), .B(G162gat), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(G99gat), .A2(G106gat), .ZN(new_n595));
  INV_X1    g394(.A(G85gat), .ZN(new_n596));
  INV_X1    g395(.A(G92gat), .ZN(new_n597));
  AOI22_X1  g396(.A1(KEYINPUT8), .A2(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(G85gat), .A2(G92gat), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT7), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g400(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n598), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G99gat), .B(G106gat), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  AND2_X1   g405(.A1(new_n601), .A2(new_n602), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n607), .A2(new_n604), .A3(new_n598), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n567), .A2(new_n568), .A3(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n609), .ZN(new_n611));
  AND2_X1   g410(.A1(G232gat), .A2(G233gat), .ZN(new_n612));
  AOI22_X1  g411(.A1(new_n538), .A2(new_n611), .B1(KEYINPUT41), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(G190gat), .B(G218gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(KEYINPUT96), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n617), .A2(KEYINPUT97), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n594), .B1(new_n614), .B2(new_n619), .ZN(new_n620));
  AOI211_X1 g419(.A(new_n618), .B(new_n593), .C1(new_n610), .C2(new_n613), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n617), .A2(KEYINPUT97), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n612), .A2(KEYINPUT41), .ZN(new_n623));
  XOR2_X1   g422(.A(new_n622), .B(new_n623), .Z(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  OR3_X1    g424(.A1(new_n620), .A2(new_n621), .A3(new_n625), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n625), .B1(new_n620), .B2(new_n621), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g427(.A(G57gat), .B(G64gat), .Z(new_n629));
  INV_X1    g428(.A(G71gat), .ZN(new_n630));
  INV_X1    g429(.A(G78gat), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(G71gat), .A2(G78gat), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT9), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n629), .A2(new_n634), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(G57gat), .B(G64gat), .ZN(new_n638));
  OAI211_X1 g437(.A(new_n633), .B(new_n632), .C1(new_n638), .C2(new_n635), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT21), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(G127gat), .B(G155gat), .ZN(new_n643));
  XOR2_X1   g442(.A(new_n642), .B(new_n643), .Z(new_n644));
  OAI21_X1  g443(.A(new_n551), .B1(new_n641), .B2(new_n640), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(KEYINPUT95), .ZN(new_n648));
  NAND2_X1  g447(.A1(G231gat), .A2(G233gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(KEYINPUT94), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n648), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(G183gat), .B(G211gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n646), .B(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n628), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(G230gat), .A2(G233gat), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n603), .A2(new_n605), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n604), .B1(new_n607), .B2(new_n598), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n640), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND4_X1  g458(.A1(new_n606), .A2(new_n608), .A3(new_n639), .A4(new_n637), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n659), .A2(KEYINPUT98), .A3(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT98), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n609), .A2(new_n662), .A3(new_n640), .ZN(new_n663));
  AOI21_X1  g462(.A(KEYINPUT10), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT10), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n660), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n656), .B1(new_n664), .B2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n656), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n661), .A2(new_n663), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g469(.A(G120gat), .B(G148gat), .Z(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(KEYINPUT99), .ZN(new_n672));
  XNOR2_X1  g471(.A(G176gat), .B(G204gat), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n672), .B(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n670), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n667), .A2(new_n669), .A3(new_n674), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n655), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n592), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n680), .A2(new_n444), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(new_n541), .ZN(G1324gat));
  INV_X1    g481(.A(new_n441), .ZN(new_n683));
  OR3_X1    g482(.A1(new_n680), .A2(KEYINPUT100), .A3(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(KEYINPUT100), .B1(new_n680), .B2(new_n683), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n684), .A2(G8gat), .A3(new_n685), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n680), .A2(new_n683), .ZN(new_n687));
  XOR2_X1   g486(.A(KEYINPUT16), .B(G8gat), .Z(new_n688));
  NAND3_X1  g487(.A1(new_n687), .A2(KEYINPUT42), .A3(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n688), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n690), .B1(new_n684), .B2(new_n685), .ZN(new_n691));
  OAI211_X1 g490(.A(new_n686), .B(new_n689), .C1(new_n691), .C2(KEYINPUT42), .ZN(G1325gat));
  OAI21_X1  g491(.A(G15gat), .B1(new_n680), .B2(new_n490), .ZN(new_n693));
  INV_X1    g492(.A(new_n489), .ZN(new_n694));
  OR2_X1    g493(.A1(new_n694), .A2(G15gat), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n693), .B1(new_n680), .B2(new_n695), .ZN(G1326gat));
  INV_X1    g495(.A(new_n453), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n680), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(KEYINPUT101), .ZN(new_n699));
  XNOR2_X1  g498(.A(KEYINPUT43), .B(G22gat), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n699), .B(new_n700), .ZN(G1327gat));
  NOR3_X1   g500(.A1(new_n628), .A2(new_n654), .A3(new_n678), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n592), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n444), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n704), .A2(new_n511), .A3(new_n705), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(KEYINPUT45), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n454), .A2(new_n490), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT103), .ZN(new_n709));
  AOI221_X4 g508(.A(new_n709), .B1(new_n499), .B2(new_n489), .C1(new_n495), .C2(KEYINPUT35), .ZN(new_n710));
  AOI21_X1  g509(.A(KEYINPUT103), .B1(new_n496), .B2(new_n500), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n708), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  XOR2_X1   g511(.A(KEYINPUT104), .B(KEYINPUT44), .Z(new_n713));
  NOR2_X1   g512(.A1(new_n628), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(KEYINPUT44), .B1(new_n501), .B2(new_n628), .ZN(new_n716));
  AND2_X1   g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT102), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n718), .B1(new_n584), .B2(new_n590), .ZN(new_n719));
  INV_X1    g518(.A(new_n581), .ZN(new_n720));
  INV_X1    g519(.A(new_n565), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n572), .A2(new_n575), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n720), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n565), .A2(new_n574), .A3(new_n582), .A4(new_n583), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n723), .A2(KEYINPUT102), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n719), .A2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(new_n654), .ZN(new_n728));
  INV_X1    g527(.A(new_n678), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n727), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  NOR3_X1   g529(.A1(new_n717), .A2(new_n444), .A3(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n707), .B1(new_n731), .B2(new_n511), .ZN(G1328gat));
  AND2_X1   g531(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n733));
  NOR2_X1   g532(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NOR3_X1   g534(.A1(new_n703), .A2(G36gat), .A3(new_n683), .ZN(new_n736));
  MUX2_X1   g535(.A(new_n735), .B(new_n733), .S(new_n736), .Z(new_n737));
  NOR3_X1   g536(.A1(new_n717), .A2(new_n683), .A3(new_n730), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n737), .B1(new_n512), .B2(new_n738), .ZN(G1329gat));
  NOR4_X1   g538(.A1(new_n717), .A2(new_n504), .A3(new_n490), .A4(new_n730), .ZN(new_n740));
  AOI21_X1  g539(.A(G43gat), .B1(new_n704), .B2(new_n489), .ZN(new_n741));
  OR3_X1    g540(.A1(new_n740), .A2(KEYINPUT47), .A3(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(KEYINPUT47), .B1(new_n740), .B2(new_n741), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(G1330gat));
  NOR2_X1   g543(.A1(new_n704), .A2(KEYINPUT106), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n520), .A2(new_n521), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT106), .ZN(new_n748));
  OAI211_X1 g547(.A(new_n453), .B(new_n747), .C1(new_n703), .C2(new_n748), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n745), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n717), .A2(new_n730), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(new_n453), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n750), .B1(new_n752), .B2(new_n746), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n747), .B1(new_n751), .B2(new_n418), .ZN(new_n754));
  OAI21_X1  g553(.A(KEYINPUT48), .B1(new_n745), .B2(new_n749), .ZN(new_n755));
  OAI22_X1  g554(.A1(new_n753), .A2(KEYINPUT48), .B1(new_n754), .B2(new_n755), .ZN(G1331gat));
  NOR3_X1   g555(.A1(new_n727), .A2(new_n655), .A3(new_n729), .ZN(new_n757));
  AND2_X1   g556(.A1(new_n712), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(new_n705), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g559(.A1(new_n712), .A2(new_n757), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n761), .A2(new_n683), .ZN(new_n762));
  NOR2_X1   g561(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n763));
  AND2_X1   g562(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n762), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n765), .B1(new_n762), .B2(new_n763), .ZN(G1333gat));
  NAND3_X1  g565(.A1(new_n758), .A2(new_n630), .A3(new_n489), .ZN(new_n767));
  OAI21_X1  g566(.A(G71gat), .B1(new_n761), .B2(new_n490), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT108), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n767), .A2(KEYINPUT108), .A3(new_n768), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g572(.A(KEYINPUT107), .B(KEYINPUT50), .ZN(new_n774));
  INV_X1    g573(.A(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n771), .A2(new_n772), .A3(new_n774), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(G1334gat));
  NOR2_X1   g577(.A1(new_n761), .A2(new_n697), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(new_n631), .ZN(G1335gat));
  NAND3_X1  g579(.A1(new_n726), .A2(new_n728), .A3(new_n678), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n781), .B1(new_n715), .B2(new_n716), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(G85gat), .B1(new_n783), .B2(new_n444), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n727), .A2(new_n654), .A3(new_n628), .ZN(new_n785));
  AND3_X1   g584(.A1(new_n712), .A2(KEYINPUT51), .A3(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(KEYINPUT51), .B1(new_n712), .B2(new_n785), .ZN(new_n787));
  OR2_X1    g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n729), .B1(new_n788), .B2(KEYINPUT109), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n789), .B1(KEYINPUT109), .B2(new_n788), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n705), .A2(new_n596), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n784), .B1(new_n790), .B2(new_n791), .ZN(G1336gat));
  NOR3_X1   g591(.A1(new_n683), .A2(G92gat), .A3(new_n729), .ZN(new_n793));
  XOR2_X1   g592(.A(KEYINPUT111), .B(KEYINPUT51), .Z(new_n794));
  AOI21_X1  g593(.A(new_n794), .B1(new_n712), .B2(new_n785), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n793), .B1(new_n786), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n597), .B1(new_n782), .B2(new_n441), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT110), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n796), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  AOI211_X1 g598(.A(KEYINPUT110), .B(new_n597), .C1(new_n782), .C2(new_n441), .ZN(new_n800));
  OAI21_X1  g599(.A(KEYINPUT52), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(KEYINPUT52), .B1(new_n788), .B2(new_n793), .ZN(new_n802));
  OAI21_X1  g601(.A(G92gat), .B1(new_n783), .B2(new_n683), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n801), .A2(new_n804), .ZN(G1337gat));
  OAI21_X1  g604(.A(G99gat), .B1(new_n783), .B2(new_n490), .ZN(new_n806));
  OR2_X1    g605(.A1(new_n694), .A2(G99gat), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n806), .B1(new_n790), .B2(new_n807), .ZN(G1338gat));
  NAND2_X1  g607(.A1(new_n782), .A2(new_n453), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(G106gat), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n417), .A2(G106gat), .A3(new_n729), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n811), .B1(new_n786), .B2(new_n795), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT112), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OAI211_X1 g613(.A(KEYINPUT112), .B(new_n811), .C1(new_n786), .C2(new_n795), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n810), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(KEYINPUT53), .ZN(new_n817));
  AOI21_X1  g616(.A(KEYINPUT53), .B1(new_n788), .B2(new_n811), .ZN(new_n818));
  OAI21_X1  g617(.A(G106gat), .B1(new_n783), .B2(new_n417), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n817), .A2(new_n820), .ZN(G1339gat));
  INV_X1    g620(.A(new_n628), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT55), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n661), .A2(new_n663), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(new_n665), .ZN(new_n825));
  INV_X1    g624(.A(new_n666), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n825), .A2(new_n826), .A3(new_n668), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n827), .A2(new_n667), .A3(KEYINPUT54), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n675), .B1(new_n667), .B2(KEYINPUT54), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n823), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT113), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n668), .B1(new_n825), .B2(new_n826), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n826), .A2(new_n668), .ZN(new_n834));
  OAI21_X1  g633(.A(KEYINPUT54), .B1(new_n664), .B2(new_n834), .ZN(new_n835));
  OAI21_X1  g634(.A(KEYINPUT55), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n832), .B1(new_n836), .B2(new_n830), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT54), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n674), .B1(new_n833), .B2(new_n838), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n839), .A2(KEYINPUT113), .A3(KEYINPUT55), .A4(new_n828), .ZN(new_n840));
  AND4_X1   g639(.A1(new_n677), .A2(new_n831), .A3(new_n837), .A4(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n719), .A2(new_n725), .A3(new_n841), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n586), .A2(new_n557), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n558), .B1(new_n556), .B2(new_n560), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n580), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n724), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n678), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n822), .B1(new_n842), .B2(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n822), .A2(new_n841), .A3(new_n846), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n728), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n679), .A2(new_n726), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n453), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n853), .A2(new_n705), .A3(new_n489), .A4(new_n683), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n854), .A2(new_n307), .A3(new_n591), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n851), .A2(new_n852), .ZN(new_n856));
  AND2_X1   g655(.A1(new_n493), .A2(new_n494), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n856), .A2(new_n705), .A3(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT114), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n444), .B1(new_n851), .B2(new_n852), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n861), .A2(KEYINPUT114), .A3(new_n857), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n441), .B1(new_n860), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(new_n727), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n855), .B1(new_n864), .B2(new_n307), .ZN(G1340gat));
  NOR3_X1   g664(.A1(new_n854), .A2(new_n305), .A3(new_n729), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n863), .A2(new_n678), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n866), .B1(new_n867), .B2(new_n305), .ZN(G1341gat));
  NOR3_X1   g667(.A1(new_n854), .A2(new_n315), .A3(new_n728), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n863), .A2(new_n654), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT115), .ZN(new_n871));
  OR2_X1    g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(G127gat), .B1(new_n870), .B2(new_n871), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n869), .B1(new_n872), .B2(new_n873), .ZN(G1342gat));
  INV_X1    g673(.A(KEYINPUT118), .ZN(new_n875));
  OAI21_X1  g674(.A(G134gat), .B1(new_n854), .B2(new_n628), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT116), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n441), .A2(G134gat), .A3(new_n628), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n879), .B1(new_n860), .B2(new_n862), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT56), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n877), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  AND4_X1   g681(.A1(KEYINPUT114), .A2(new_n856), .A3(new_n705), .A4(new_n857), .ZN(new_n883));
  AOI21_X1  g682(.A(KEYINPUT114), .B1(new_n861), .B2(new_n857), .ZN(new_n884));
  OAI211_X1 g683(.A(new_n881), .B(new_n878), .C1(new_n883), .C2(new_n884), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n885), .A2(KEYINPUT116), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n876), .B1(new_n882), .B2(new_n886), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n880), .A2(KEYINPUT117), .A3(new_n881), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT117), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n878), .B1(new_n883), .B2(new_n884), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n889), .B1(new_n890), .B2(KEYINPUT56), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n875), .B1(new_n887), .B2(new_n892), .ZN(new_n893));
  XNOR2_X1  g692(.A(new_n885), .B(KEYINPUT116), .ZN(new_n894));
  OAI21_X1  g693(.A(KEYINPUT117), .B1(new_n880), .B2(new_n881), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n890), .A2(new_n889), .A3(KEYINPUT56), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND4_X1  g696(.A1(new_n894), .A2(KEYINPUT118), .A3(new_n897), .A4(new_n876), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n893), .A2(new_n898), .ZN(G1343gat));
  INV_X1    g698(.A(new_n490), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n900), .A2(new_n417), .A3(new_n441), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n861), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n591), .A2(G141gat), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT58), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NOR3_X1   g705(.A1(new_n900), .A2(new_n444), .A3(new_n441), .ZN(new_n907));
  INV_X1    g706(.A(new_n907), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n417), .B1(new_n851), .B2(new_n852), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT57), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n908), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  AND3_X1   g710(.A1(new_n837), .A2(new_n840), .A3(new_n677), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT119), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n913), .B1(new_n829), .B2(new_n830), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n839), .A2(KEYINPUT119), .A3(new_n828), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n914), .A2(new_n823), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n912), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n591), .B1(new_n917), .B2(KEYINPUT120), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT120), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n912), .A2(new_n919), .A3(new_n916), .ZN(new_n920));
  AOI22_X1  g719(.A1(new_n918), .A2(new_n920), .B1(new_n678), .B2(new_n846), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n849), .B1(new_n921), .B2(new_n822), .ZN(new_n922));
  AOI22_X1  g721(.A1(new_n922), .A2(new_n728), .B1(new_n679), .B2(new_n726), .ZN(new_n923));
  OAI21_X1  g722(.A(KEYINPUT57), .B1(new_n923), .B2(new_n697), .ZN(new_n924));
  OAI211_X1 g723(.A(new_n911), .B(new_n924), .C1(new_n590), .C2(new_n584), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n906), .B1(new_n925), .B2(G141gat), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n926), .A2(KEYINPUT121), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n926), .A2(KEYINPUT121), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n911), .A2(new_n924), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n929), .A2(new_n727), .ZN(new_n930));
  AOI22_X1  g729(.A1(new_n930), .A2(G141gat), .B1(new_n902), .B2(new_n903), .ZN(new_n931));
  OAI22_X1  g730(.A1(new_n927), .A2(new_n928), .B1(new_n905), .B2(new_n931), .ZN(G1344gat));
  NAND3_X1  g731(.A1(new_n902), .A2(new_n330), .A3(new_n678), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT59), .ZN(new_n934));
  INV_X1    g733(.A(new_n909), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(KEYINPUT57), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n908), .A2(new_n729), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n654), .B1(new_n922), .B2(KEYINPUT122), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT122), .ZN(new_n939));
  OAI211_X1 g738(.A(new_n939), .B(new_n849), .C1(new_n921), .C2(new_n822), .ZN(new_n940));
  AOI22_X1  g739(.A1(new_n938), .A2(new_n940), .B1(new_n591), .B2(new_n679), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n453), .A2(new_n910), .ZN(new_n942));
  OAI211_X1 g741(.A(new_n936), .B(new_n937), .C1(new_n941), .C2(new_n942), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n934), .B1(new_n943), .B2(G148gat), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n934), .A2(G148gat), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n945), .B1(new_n929), .B2(new_n678), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n933), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT123), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  OAI211_X1 g748(.A(KEYINPUT123), .B(new_n933), .C1(new_n944), .C2(new_n946), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(G1345gat));
  AOI21_X1  g750(.A(new_n334), .B1(new_n929), .B2(new_n654), .ZN(new_n952));
  AND3_X1   g751(.A1(new_n902), .A2(new_n334), .A3(new_n654), .ZN(new_n953));
  OR2_X1    g752(.A1(new_n952), .A2(new_n953), .ZN(G1346gat));
  AOI21_X1  g753(.A(G162gat), .B1(new_n902), .B2(new_n822), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n628), .A2(new_n335), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n955), .B1(new_n929), .B2(new_n956), .ZN(G1347gat));
  NOR2_X1   g756(.A1(new_n683), .A2(new_n705), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n856), .A2(new_n857), .A3(new_n958), .ZN(new_n959));
  INV_X1    g758(.A(new_n959), .ZN(new_n960));
  AOI21_X1  g759(.A(G169gat), .B1(new_n960), .B2(new_n727), .ZN(new_n961));
  AND3_X1   g760(.A1(new_n853), .A2(new_n489), .A3(new_n958), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n591), .A2(new_n221), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n961), .B1(new_n962), .B2(new_n963), .ZN(G1348gat));
  NAND3_X1  g763(.A1(new_n962), .A2(G176gat), .A3(new_n678), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT124), .ZN(new_n966));
  AND2_X1   g765(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n965), .A2(new_n966), .ZN(new_n968));
  AOI21_X1  g767(.A(G176gat), .B1(new_n960), .B2(new_n678), .ZN(new_n969));
  NOR3_X1   g768(.A1(new_n967), .A2(new_n968), .A3(new_n969), .ZN(G1349gat));
  AOI21_X1  g769(.A(new_n230), .B1(new_n962), .B2(new_n654), .ZN(new_n971));
  AND2_X1   g770(.A1(new_n654), .A2(new_n238), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n971), .B1(new_n960), .B2(new_n972), .ZN(new_n973));
  XOR2_X1   g772(.A(new_n973), .B(KEYINPUT60), .Z(G1350gat));
  NAND3_X1  g773(.A1(new_n960), .A2(new_n234), .A3(new_n822), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n962), .A2(new_n822), .ZN(new_n976));
  NOR2_X1   g775(.A1(KEYINPUT125), .A2(KEYINPUT61), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n234), .B1(KEYINPUT125), .B2(KEYINPUT61), .ZN(new_n978));
  AND3_X1   g777(.A1(new_n976), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n977), .B1(new_n976), .B2(new_n978), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n975), .B1(new_n979), .B2(new_n980), .ZN(G1351gat));
  OR2_X1    g780(.A1(new_n941), .A2(new_n942), .ZN(new_n982));
  AND2_X1   g781(.A1(new_n490), .A2(new_n958), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n982), .A2(new_n936), .A3(new_n983), .ZN(new_n984));
  INV_X1    g783(.A(G197gat), .ZN(new_n985));
  NOR3_X1   g784(.A1(new_n984), .A2(new_n985), .A3(new_n591), .ZN(new_n986));
  AND2_X1   g785(.A1(new_n909), .A2(new_n983), .ZN(new_n987));
  AOI21_X1  g786(.A(G197gat), .B1(new_n987), .B2(new_n727), .ZN(new_n988));
  NOR2_X1   g787(.A1(new_n986), .A2(new_n988), .ZN(G1352gat));
  INV_X1    g788(.A(G204gat), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n987), .A2(new_n990), .A3(new_n678), .ZN(new_n991));
  AND2_X1   g790(.A1(new_n991), .A2(KEYINPUT126), .ZN(new_n992));
  NOR2_X1   g791(.A1(new_n991), .A2(KEYINPUT126), .ZN(new_n993));
  INV_X1    g792(.A(KEYINPUT62), .ZN(new_n994));
  OR3_X1    g793(.A1(new_n992), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  OAI21_X1  g794(.A(G204gat), .B1(new_n984), .B2(new_n729), .ZN(new_n996));
  OAI21_X1  g795(.A(new_n994), .B1(new_n992), .B2(new_n993), .ZN(new_n997));
  NAND3_X1  g796(.A1(new_n995), .A2(new_n996), .A3(new_n997), .ZN(G1353gat));
  NAND3_X1  g797(.A1(new_n987), .A2(new_n213), .A3(new_n654), .ZN(new_n999));
  INV_X1    g798(.A(KEYINPUT127), .ZN(new_n1000));
  NAND4_X1  g799(.A1(new_n982), .A2(new_n654), .A3(new_n936), .A4(new_n983), .ZN(new_n1001));
  AND4_X1   g800(.A1(new_n1000), .A2(new_n1001), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n1002));
  INV_X1    g801(.A(KEYINPUT63), .ZN(new_n1003));
  AOI21_X1  g802(.A(new_n205), .B1(KEYINPUT127), .B2(new_n1003), .ZN(new_n1004));
  AOI22_X1  g803(.A1(new_n1001), .A2(new_n1004), .B1(new_n1000), .B2(KEYINPUT63), .ZN(new_n1005));
  OAI21_X1  g804(.A(new_n999), .B1(new_n1002), .B2(new_n1005), .ZN(G1354gat));
  OAI21_X1  g805(.A(G218gat), .B1(new_n984), .B2(new_n628), .ZN(new_n1007));
  NAND3_X1  g806(.A1(new_n987), .A2(new_n204), .A3(new_n822), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n1007), .A2(new_n1008), .ZN(G1355gat));
endmodule


