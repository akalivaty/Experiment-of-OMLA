//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 1 1 0 0 0 0 0 1 1 0 0 1 0 1 1 1 0 0 0 0 0 0 1 0 0 0 1 0 0 1 0 0 1 0 0 0 1 0 1 0 0 0 1 0 0 0 1 1 0 0 0 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:09 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1128, new_n1129, new_n1130, new_n1131, new_n1132, new_n1133,
    new_n1134, new_n1135, new_n1136, new_n1137, new_n1138, new_n1139,
    new_n1140, new_n1141, new_n1142, new_n1143, new_n1144, new_n1145,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1168, new_n1169, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1222, new_n1223, new_n1224, new_n1225;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XOR2_X1   g0003(.A(new_n203), .B(KEYINPUT64), .Z(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  AND2_X1   g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(G20), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT65), .ZN(new_n212));
  OAI21_X1  g0012(.A(G50), .B1(G58), .B2(G68), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n214));
  INV_X1    g0014(.A(G244), .ZN(new_n215));
  INV_X1    g0015(.A(G87), .ZN(new_n216));
  INV_X1    g0016(.A(G250), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n214), .B1(new_n202), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n219));
  INV_X1    g0019(.A(G58), .ZN(new_n220));
  INV_X1    g0020(.A(G232), .ZN(new_n221));
  INV_X1    g0021(.A(G68), .ZN(new_n222));
  INV_X1    g0022(.A(G238), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n206), .B1(new_n218), .B2(new_n224), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n209), .B1(new_n212), .B2(new_n213), .C1(KEYINPUT1), .C2(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT2), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(G226), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(new_n221), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G264), .B(G270), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n231), .B(new_n234), .ZN(G358));
  XOR2_X1   g0035(.A(G68), .B(G77), .Z(new_n236));
  XOR2_X1   g0036(.A(G50), .B(G58), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G351));
  NAND2_X1  g0042(.A1(G33), .A2(G41), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n210), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(KEYINPUT3), .B(G33), .ZN(new_n245));
  INV_X1    g0045(.A(G1698), .ZN(new_n246));
  AND2_X1   g0046(.A1(new_n246), .A2(G222), .ZN(new_n247));
  INV_X1    g0047(.A(G223), .ZN(new_n248));
  NOR2_X1   g0048(.A1(new_n248), .A2(new_n246), .ZN(new_n249));
  OAI21_X1  g0049(.A(new_n245), .B1(new_n247), .B2(new_n249), .ZN(new_n250));
  OAI21_X1  g0050(.A(new_n250), .B1(new_n202), .B2(new_n245), .ZN(new_n251));
  AOI21_X1  g0051(.A(new_n244), .B1(new_n251), .B2(KEYINPUT66), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n252), .B1(KEYINPUT66), .B2(new_n251), .ZN(new_n253));
  INV_X1    g0053(.A(G274), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n254), .B1(new_n210), .B2(new_n243), .ZN(new_n255));
  INV_X1    g0055(.A(G1), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n256), .B1(G41), .B2(G45), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n255), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n244), .A2(new_n257), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G226), .ZN(new_n262));
  AND3_X1   g0062(.A1(new_n253), .A2(new_n259), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G190), .ZN(new_n264));
  XNOR2_X1  g0064(.A(KEYINPUT71), .B(G200), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  OAI211_X1 g0066(.A(new_n264), .B(KEYINPUT73), .C1(new_n266), .C2(new_n263), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT10), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n263), .A2(new_n266), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n270), .B1(G190), .B2(new_n263), .ZN(new_n271));
  NOR2_X1   g0071(.A1(KEYINPUT72), .A2(KEYINPUT9), .ZN(new_n272));
  NOR2_X1   g0072(.A1(G20), .A2(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G150), .ZN(new_n274));
  INV_X1    g0074(.A(G20), .ZN(new_n275));
  XNOR2_X1  g0075(.A(KEYINPUT8), .B(G58), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(G33), .ZN(new_n277));
  OAI221_X1 g0077(.A(new_n274), .B1(new_n201), .B2(new_n275), .C1(new_n276), .C2(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(G1), .A2(G13), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n256), .A2(G13), .A3(G20), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT67), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND4_X1  g0084(.A1(new_n256), .A2(KEYINPUT67), .A3(G13), .A4(G20), .ZN(new_n285));
  AND2_X1   g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G50), .ZN(new_n287));
  AOI22_X1  g0087(.A1(new_n278), .A2(new_n281), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n284), .A2(new_n285), .ZN(new_n289));
  INV_X1    g0089(.A(new_n281), .ZN(new_n290));
  OAI211_X1 g0090(.A(new_n289), .B(new_n290), .C1(G1), .C2(new_n275), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n288), .B1(new_n287), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(KEYINPUT72), .A2(KEYINPUT9), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n272), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n292), .A2(new_n272), .ZN(new_n296));
  NAND4_X1  g0096(.A1(new_n269), .A2(new_n271), .A3(new_n295), .A4(new_n296), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n271), .A2(new_n295), .A3(new_n296), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n298), .A2(new_n268), .A3(new_n267), .ZN(new_n299));
  INV_X1    g0099(.A(G179), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n263), .A2(new_n300), .ZN(new_n301));
  OAI211_X1 g0101(.A(new_n301), .B(new_n292), .C1(G169), .C2(new_n263), .ZN(new_n302));
  NAND2_X1  g0102(.A1(G238), .A2(G1698), .ZN(new_n303));
  OAI211_X1 g0103(.A(new_n245), .B(new_n303), .C1(new_n221), .C2(G1698), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n280), .B1(G33), .B2(G41), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n304), .B(new_n305), .C1(G107), .C2(new_n245), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n261), .A2(G244), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n306), .A2(new_n259), .A3(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT68), .ZN(new_n309));
  OR2_X1    g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n308), .A2(new_n309), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(G190), .ZN(new_n313));
  XNOR2_X1  g0113(.A(KEYINPUT15), .B(G87), .ZN(new_n314));
  OAI22_X1  g0114(.A1(new_n314), .A2(new_n277), .B1(new_n275), .B2(new_n202), .ZN(new_n315));
  XNOR2_X1  g0115(.A(new_n276), .B(KEYINPUT69), .ZN(new_n316));
  XNOR2_X1  g0116(.A(new_n273), .B(KEYINPUT70), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n315), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n318), .A2(new_n290), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n291), .A2(new_n202), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n289), .A2(G77), .ZN(new_n321));
  NOR3_X1   g0121(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  OAI211_X1 g0122(.A(new_n313), .B(new_n322), .C1(new_n266), .C2(new_n312), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n312), .A2(new_n300), .ZN(new_n324));
  INV_X1    g0124(.A(new_n322), .ZN(new_n325));
  INV_X1    g0125(.A(G169), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n310), .A2(new_n326), .A3(new_n311), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n324), .A2(new_n325), .A3(new_n327), .ZN(new_n328));
  AND2_X1   g0128(.A1(new_n323), .A2(new_n328), .ZN(new_n329));
  AND4_X1   g0129(.A1(new_n297), .A2(new_n299), .A3(new_n302), .A4(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT18), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT7), .ZN(new_n332));
  NOR3_X1   g0132(.A1(new_n245), .A2(new_n332), .A3(G20), .ZN(new_n333));
  AND2_X1   g0133(.A1(KEYINPUT3), .A2(G33), .ZN(new_n334));
  NOR2_X1   g0134(.A1(KEYINPUT3), .A2(G33), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(KEYINPUT7), .B1(new_n336), .B2(new_n275), .ZN(new_n337));
  OAI21_X1  g0137(.A(G68), .B1(new_n333), .B2(new_n337), .ZN(new_n338));
  XNOR2_X1  g0138(.A(G58), .B(G68), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n339), .A2(G20), .B1(G159), .B2(new_n273), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT16), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n290), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n338), .A2(KEYINPUT16), .A3(new_n340), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n286), .A2(new_n276), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n346), .B1(new_n291), .B2(new_n276), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n248), .A2(new_n246), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n245), .B(new_n350), .C1(G226), .C2(new_n246), .ZN(new_n351));
  NAND2_X1  g0151(.A1(G33), .A2(G87), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n244), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n259), .B1(new_n221), .B2(new_n260), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(new_n300), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n356), .B1(G169), .B2(new_n355), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n331), .B1(new_n349), .B2(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n347), .B1(new_n343), .B2(new_n344), .ZN(new_n360));
  NOR3_X1   g0160(.A1(new_n360), .A2(KEYINPUT18), .A3(new_n357), .ZN(new_n361));
  OAI21_X1  g0161(.A(KEYINPUT76), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n349), .A2(new_n358), .A3(new_n331), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT76), .ZN(new_n364));
  OAI21_X1  g0164(.A(KEYINPUT18), .B1(new_n360), .B2(new_n357), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(G200), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n355), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n368), .B1(G190), .B2(new_n355), .ZN(new_n369));
  XNOR2_X1  g0169(.A(KEYINPUT77), .B(KEYINPUT17), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n369), .A2(new_n360), .A3(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT78), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n369), .A2(new_n360), .ZN(new_n374));
  AOI22_X1  g0174(.A1(new_n372), .A2(new_n373), .B1(new_n374), .B2(KEYINPUT17), .ZN(new_n375));
  OR2_X1    g0175(.A1(new_n372), .A2(new_n373), .ZN(new_n376));
  AOI22_X1  g0176(.A1(new_n362), .A2(new_n366), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n286), .A2(KEYINPUT12), .A3(new_n222), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT12), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n379), .B1(new_n289), .B2(G68), .ZN(new_n380));
  OAI211_X1 g0180(.A(new_n378), .B(new_n380), .C1(new_n291), .C2(new_n222), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT75), .ZN(new_n382));
  OR2_X1    g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n381), .A2(new_n382), .ZN(new_n384));
  AOI22_X1  g0184(.A1(new_n273), .A2(G50), .B1(G20), .B2(new_n222), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n385), .B1(new_n202), .B2(new_n277), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(new_n281), .ZN(new_n387));
  XNOR2_X1  g0187(.A(new_n387), .B(KEYINPUT11), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n383), .A2(new_n384), .A3(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n259), .B1(new_n223), .B2(new_n260), .ZN(new_n390));
  NAND2_X1  g0190(.A1(G33), .A2(G97), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n221), .A2(G1698), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n392), .B1(G226), .B2(G1698), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n391), .B1(new_n393), .B2(new_n336), .ZN(new_n394));
  OR2_X1    g0194(.A1(new_n394), .A2(KEYINPUT74), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n244), .B1(new_n394), .B2(KEYINPUT74), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n390), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT13), .ZN(new_n398));
  XNOR2_X1  g0198(.A(new_n397), .B(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT14), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n399), .A2(new_n400), .A3(G169), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n401), .B1(new_n300), .B2(new_n399), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n400), .B1(new_n399), .B2(G169), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n389), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n389), .B1(G200), .B2(new_n399), .ZN(new_n405));
  INV_X1    g0205(.A(G190), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n405), .B1(new_n406), .B2(new_n399), .ZN(new_n407));
  AND2_X1   g0207(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  AND3_X1   g0208(.A1(new_n330), .A2(new_n377), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(KEYINPUT85), .A2(KEYINPUT25), .ZN(new_n410));
  INV_X1    g0210(.A(G107), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n411), .B1(KEYINPUT85), .B2(KEYINPUT25), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n410), .B1(new_n289), .B2(new_n412), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n286), .A2(KEYINPUT85), .A3(KEYINPUT25), .A4(new_n411), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT79), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n415), .B1(new_n256), .B2(G33), .ZN(new_n416));
  INV_X1    g0216(.A(G33), .ZN(new_n417));
  NOR3_X1   g0217(.A1(new_n417), .A2(KEYINPUT79), .A3(G1), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  AND3_X1   g0219(.A1(new_n289), .A2(new_n419), .A3(new_n290), .ZN(new_n420));
  AOI22_X1  g0220(.A1(new_n413), .A2(new_n414), .B1(new_n420), .B2(G107), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n245), .A2(new_n275), .A3(G87), .ZN(new_n422));
  AND2_X1   g0222(.A1(KEYINPUT83), .A2(KEYINPUT22), .ZN(new_n423));
  NOR2_X1   g0223(.A1(KEYINPUT83), .A2(KEYINPUT22), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n422), .A2(new_n425), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n245), .A2(new_n275), .A3(G87), .A4(new_n423), .ZN(new_n427));
  NAND2_X1  g0227(.A1(G33), .A2(G116), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n428), .A2(G20), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT23), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n430), .B1(new_n275), .B2(G107), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n411), .A2(KEYINPUT23), .A3(G20), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n429), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n426), .A2(new_n427), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(KEYINPUT84), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT84), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n426), .A2(new_n436), .A3(new_n427), .A4(new_n433), .ZN(new_n437));
  AND3_X1   g0237(.A1(new_n435), .A2(KEYINPUT24), .A3(new_n437), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n281), .B1(new_n435), .B2(KEYINPUT24), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n421), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(G41), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n256), .B(G45), .C1(new_n441), .C2(KEYINPUT5), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT5), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n444), .A2(G41), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n443), .A2(new_n255), .A3(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT88), .ZN(new_n448));
  OAI211_X1 g0248(.A(G250), .B(new_n246), .C1(new_n334), .C2(new_n335), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(KEYINPUT86), .ZN(new_n450));
  INV_X1    g0250(.A(G294), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n417), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(G257), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n453), .A2(new_n246), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n452), .B1(new_n245), .B2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT86), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n245), .A2(new_n456), .A3(G250), .A4(new_n246), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n450), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n305), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n244), .B(G264), .C1(new_n442), .C2(new_n445), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n448), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n460), .ZN(new_n462));
  AOI211_X1 g0262(.A(KEYINPUT88), .B(new_n462), .C1(new_n458), .C2(new_n305), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n447), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(new_n367), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n462), .B1(new_n458), .B2(new_n305), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n447), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT87), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n466), .A2(KEYINPUT87), .A3(new_n447), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n469), .A2(new_n406), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n440), .B1(new_n465), .B2(new_n471), .ZN(new_n472));
  OAI211_X1 g0272(.A(G179), .B(new_n447), .C1(new_n461), .C2(new_n463), .ZN(new_n473));
  AND4_X1   g0273(.A1(KEYINPUT87), .A2(new_n459), .A3(new_n447), .A4(new_n460), .ZN(new_n474));
  AOI21_X1  g0274(.A(KEYINPUT87), .B1(new_n466), .B2(new_n447), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n473), .B1(new_n476), .B2(new_n326), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n472), .B1(new_n477), .B2(new_n440), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT4), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n479), .A2(G1698), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n480), .B(G244), .C1(new_n335), .C2(new_n334), .ZN(new_n481));
  NAND2_X1  g0281(.A1(G33), .A2(G283), .ZN(new_n482));
  OR2_X1    g0282(.A1(KEYINPUT3), .A2(G33), .ZN(new_n483));
  NAND2_X1  g0283(.A1(KEYINPUT3), .A2(G33), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n215), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n481), .B(new_n482), .C1(new_n485), .C2(KEYINPUT4), .ZN(new_n486));
  OAI21_X1  g0286(.A(G250), .B1(new_n334), .B2(new_n335), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n246), .B1(new_n487), .B2(KEYINPUT4), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n305), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n244), .B(G257), .C1(new_n442), .C2(new_n445), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n447), .A2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n273), .A2(G77), .ZN(new_n494));
  AND3_X1   g0294(.A1(new_n411), .A2(KEYINPUT6), .A3(G97), .ZN(new_n495));
  XNOR2_X1  g0295(.A(G97), .B(G107), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT6), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n494), .B1(new_n498), .B2(new_n275), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n332), .B1(new_n245), .B2(G20), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n336), .A2(KEYINPUT7), .A3(new_n275), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n411), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n281), .B1(new_n499), .B2(new_n502), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n289), .A2(G97), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n504), .B1(new_n420), .B2(G97), .ZN(new_n505));
  AOI22_X1  g0305(.A1(new_n493), .A2(new_n326), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n489), .A2(KEYINPUT80), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT80), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n508), .B(new_n305), .C1(new_n486), .C2(new_n488), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n507), .A2(new_n300), .A3(new_n509), .A4(new_n492), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(G97), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n216), .A2(new_n512), .A3(new_n411), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n391), .A2(new_n275), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n513), .A2(new_n514), .A3(KEYINPUT19), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n275), .B(G68), .C1(new_n334), .C2(new_n335), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT19), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n517), .B1(new_n277), .B2(new_n512), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n515), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(new_n281), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n286), .A2(new_n314), .ZN(new_n521));
  INV_X1    g0321(.A(new_n314), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n289), .A2(new_n419), .A3(new_n290), .A4(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n520), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n223), .A2(new_n246), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n215), .A2(G1698), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n525), .B(new_n526), .C1(new_n334), .C2(new_n335), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n244), .B1(new_n527), .B2(new_n428), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n256), .A2(new_n254), .A3(G45), .ZN(new_n529));
  INV_X1    g0329(.A(G45), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n217), .B1(new_n530), .B2(G1), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n244), .A2(new_n529), .A3(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n326), .B1(new_n528), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g0334(.A1(G238), .A2(G1698), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n535), .B1(new_n215), .B2(G1698), .ZN(new_n536));
  AOI22_X1  g0336(.A1(new_n536), .A2(new_n245), .B1(G33), .B2(G116), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n300), .B(new_n532), .C1(new_n537), .C2(new_n244), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n524), .A2(new_n534), .A3(new_n538), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n519), .A2(new_n281), .B1(new_n286), .B2(new_n314), .ZN(new_n540));
  OAI211_X1 g0340(.A(G190), .B(new_n532), .C1(new_n537), .C2(new_n244), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n265), .B1(new_n528), .B2(new_n533), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n289), .A2(new_n419), .A3(new_n290), .A4(G87), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n540), .A2(new_n541), .A3(new_n542), .A4(new_n543), .ZN(new_n544));
  AND2_X1   g0344(.A1(new_n539), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n491), .B1(new_n489), .B2(KEYINPUT80), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n367), .B1(new_n546), .B2(new_n509), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n503), .B(new_n505), .C1(new_n493), .C2(new_n406), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n511), .B(new_n545), .C1(new_n547), .C2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n420), .A2(G116), .ZN(new_n550));
  INV_X1    g0350(.A(G116), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n279), .A2(new_n280), .B1(G20), .B2(new_n551), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n482), .B(new_n275), .C1(G33), .C2(new_n512), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n552), .A2(KEYINPUT20), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(KEYINPUT82), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT82), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n552), .A2(new_n556), .A3(new_n553), .A4(KEYINPUT20), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n552), .A2(new_n553), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT20), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n555), .A2(new_n557), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n286), .A2(new_n551), .ZN(new_n562));
  AND3_X1   g0362(.A1(new_n550), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(G303), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n483), .A2(new_n564), .A3(new_n484), .ZN(new_n565));
  NAND2_X1  g0365(.A1(G264), .A2(G1698), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n566), .B1(new_n453), .B2(G1698), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n565), .B(new_n305), .C1(new_n336), .C2(new_n567), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n244), .B(G270), .C1(new_n442), .C2(new_n445), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n568), .A2(new_n447), .A3(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT81), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n568), .A2(new_n447), .A3(KEYINPUT81), .A4(new_n569), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n572), .A2(G200), .A3(new_n573), .ZN(new_n574));
  AND2_X1   g0374(.A1(new_n572), .A2(new_n573), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n563), .B(new_n574), .C1(new_n575), .C2(new_n406), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n550), .A2(new_n561), .A3(new_n562), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n575), .A2(KEYINPUT21), .A3(G169), .A4(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT21), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n572), .A2(G169), .A3(new_n573), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n579), .B1(new_n563), .B2(new_n580), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n570), .A2(new_n300), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n577), .A2(new_n582), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n576), .A2(new_n578), .A3(new_n581), .A4(new_n583), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n549), .A2(new_n584), .ZN(new_n585));
  AND3_X1   g0385(.A1(new_n409), .A2(new_n478), .A3(new_n585), .ZN(G372));
  NAND2_X1  g0386(.A1(new_n546), .A2(new_n509), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(G200), .ZN(new_n588));
  AND3_X1   g0388(.A1(new_n489), .A2(G190), .A3(new_n492), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n503), .A2(new_n505), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n588), .A2(new_n591), .B1(new_n506), .B2(new_n510), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n476), .A2(new_n406), .B1(new_n464), .B2(new_n367), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n592), .B(new_n545), .C1(new_n593), .C2(new_n440), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n578), .A2(new_n581), .A3(new_n583), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n595), .B1(new_n477), .B2(new_n440), .ZN(new_n596));
  OAI21_X1  g0396(.A(KEYINPUT89), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n539), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT26), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n539), .A2(new_n544), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n599), .B1(new_n511), .B2(new_n600), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n545), .A2(KEYINPUT26), .A3(new_n510), .A4(new_n506), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n598), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n472), .A2(new_n549), .ZN(new_n604));
  INV_X1    g0404(.A(new_n473), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n326), .B1(new_n469), .B2(new_n470), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n440), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(new_n595), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT89), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n604), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n597), .A2(new_n603), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n409), .A2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n302), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n359), .A2(new_n361), .ZN(new_n615));
  INV_X1    g0415(.A(new_n404), .ZN(new_n616));
  INV_X1    g0416(.A(new_n328), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n616), .B1(new_n407), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n375), .A2(new_n376), .ZN(new_n619));
  INV_X1    g0419(.A(new_n619), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n615), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  AND2_X1   g0421(.A1(new_n299), .A2(new_n297), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n614), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n613), .A2(new_n623), .ZN(G369));
  NAND3_X1  g0424(.A1(new_n256), .A2(new_n275), .A3(G13), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n625), .A2(KEYINPUT27), .ZN(new_n626));
  XOR2_X1   g0426(.A(new_n626), .B(KEYINPUT90), .Z(new_n627));
  INV_X1    g0427(.A(G213), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n625), .A2(KEYINPUT27), .ZN(new_n630));
  XOR2_X1   g0430(.A(new_n630), .B(KEYINPUT91), .Z(new_n631));
  NAND2_X1  g0431(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(G343), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n607), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n608), .A2(new_n634), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n635), .B1(new_n478), .B2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n634), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n607), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n440), .A2(new_n634), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n639), .B1(new_n478), .B2(new_n640), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n638), .A2(new_n563), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n595), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n643), .B1(new_n584), .B2(new_n642), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(G330), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n637), .B1(new_n641), .B2(new_n645), .ZN(G399));
  INV_X1    g0446(.A(new_n207), .ZN(new_n647));
  OAI21_X1  g0447(.A(KEYINPUT92), .B1(new_n647), .B2(G41), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  NOR3_X1   g0449(.A1(new_n647), .A2(KEYINPUT92), .A3(G41), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NOR4_X1   g0451(.A1(new_n651), .A2(new_n256), .A3(G116), .A4(new_n513), .ZN(new_n652));
  INV_X1    g0452(.A(new_n213), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n652), .B1(new_n653), .B2(new_n651), .ZN(new_n654));
  XOR2_X1   g0454(.A(new_n654), .B(KEYINPUT28), .Z(new_n655));
  INV_X1    g0455(.A(G330), .ZN(new_n656));
  XOR2_X1   g0456(.A(KEYINPUT93), .B(KEYINPUT31), .Z(new_n657));
  NOR2_X1   g0457(.A1(new_n528), .A2(new_n533), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n658), .A2(G179), .ZN(new_n659));
  AND4_X1   g0459(.A1(new_n464), .A2(new_n575), .A3(new_n587), .A4(new_n659), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n658), .B1(new_n461), .B2(new_n463), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT94), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  OAI211_X1 g0463(.A(KEYINPUT94), .B(new_n658), .C1(new_n461), .C2(new_n463), .ZN(new_n664));
  NOR3_X1   g0464(.A1(new_n493), .A2(new_n300), .A3(new_n570), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n663), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g0466(.A(KEYINPUT95), .B(KEYINPUT30), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n660), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT96), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n663), .A2(KEYINPUT30), .A3(new_n664), .A4(new_n665), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n671), .B1(new_n668), .B2(new_n669), .ZN(new_n672));
  OAI211_X1 g0472(.A(new_n634), .B(new_n657), .C1(new_n670), .C2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n472), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n585), .A2(new_n607), .A3(new_n674), .A4(new_n638), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(KEYINPUT31), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n638), .B1(new_n668), .B2(new_n671), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n656), .B1(new_n673), .B2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(KEYINPUT98), .B1(new_n594), .B2(new_n596), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT97), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n602), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(new_n601), .ZN(new_n684));
  OAI211_X1 g0484(.A(new_n682), .B(new_n599), .C1(new_n511), .C2(new_n600), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n598), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT98), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n604), .A2(new_n609), .A3(new_n687), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n681), .A2(new_n686), .A3(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n689), .A2(KEYINPUT99), .A3(new_n638), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  AOI21_X1  g0491(.A(KEYINPUT99), .B1(new_n689), .B2(new_n638), .ZN(new_n692));
  OAI21_X1  g0492(.A(KEYINPUT29), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n612), .A2(new_n638), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT29), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n680), .B1(new_n693), .B2(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n655), .B1(new_n697), .B2(G1), .ZN(G364));
  NAND2_X1  g0498(.A1(new_n275), .A2(G13), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n256), .B1(new_n700), .B2(G45), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n651), .A2(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n703), .B1(new_n644), .B2(G330), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(G330), .B2(new_n644), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n245), .A2(new_n207), .ZN(new_n706));
  INV_X1    g0506(.A(G355), .ZN(new_n707));
  OAI22_X1  g0507(.A1(new_n706), .A2(new_n707), .B1(G116), .B2(new_n207), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n238), .A2(G45), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n647), .A2(new_n245), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n711), .B1(new_n530), .B2(new_n653), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n708), .B1(new_n709), .B2(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(G13), .A2(G33), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(G20), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n280), .B1(G20), .B2(new_n326), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n703), .B1(new_n713), .B2(new_n719), .ZN(new_n720));
  NOR3_X1   g0520(.A1(new_n275), .A2(new_n300), .A3(new_n367), .ZN(new_n721));
  OR2_X1    g0521(.A1(new_n721), .A2(KEYINPUT101), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(KEYINPUT101), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(new_n406), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n722), .A2(new_n406), .A3(new_n723), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  XNOR2_X1  g0527(.A(KEYINPUT33), .B(G317), .ZN(new_n728));
  AOI22_X1  g0528(.A1(G326), .A2(new_n725), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n300), .A2(G200), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n275), .A2(G190), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(G311), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n336), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n730), .A2(G20), .A3(G190), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n734), .B1(G322), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n731), .A2(new_n300), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n266), .A2(new_n738), .ZN(new_n739));
  NOR3_X1   g0539(.A1(new_n406), .A2(G179), .A3(G200), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(new_n275), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  AOI22_X1  g0542(.A1(new_n739), .A2(G283), .B1(new_n742), .B2(G294), .ZN(new_n743));
  NOR3_X1   g0543(.A1(new_n275), .A2(new_n406), .A3(G179), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n265), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n738), .A2(G200), .ZN(new_n747));
  AOI22_X1  g0547(.A1(new_n746), .A2(G303), .B1(new_n747), .B2(G329), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n729), .A2(new_n737), .A3(new_n743), .A4(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n741), .A2(new_n512), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n245), .B1(new_n745), .B2(new_n216), .ZN(new_n751));
  AOI211_X1 g0551(.A(new_n750), .B(new_n751), .C1(G107), .C2(new_n739), .ZN(new_n752));
  INV_X1    g0552(.A(new_n725), .ZN(new_n753));
  OAI221_X1 g0553(.A(new_n752), .B1(new_n222), .B2(new_n726), .C1(new_n287), .C2(new_n753), .ZN(new_n754));
  OAI22_X1  g0554(.A1(new_n735), .A2(new_n220), .B1(new_n732), .B2(new_n202), .ZN(new_n755));
  XNOR2_X1  g0555(.A(new_n755), .B(KEYINPUT100), .ZN(new_n756));
  INV_X1    g0556(.A(new_n747), .ZN(new_n757));
  INV_X1    g0557(.A(G159), .ZN(new_n758));
  OAI21_X1  g0558(.A(KEYINPUT32), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  OR3_X1    g0559(.A1(new_n757), .A2(KEYINPUT32), .A3(new_n758), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n756), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n749), .B1(new_n754), .B2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(KEYINPUT102), .ZN(new_n763));
  OR2_X1    g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n717), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n765), .B1(new_n762), .B2(new_n763), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n720), .B1(new_n764), .B2(new_n766), .ZN(new_n767));
  XNOR2_X1  g0567(.A(new_n716), .B(KEYINPUT103), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n767), .B1(new_n644), .B2(new_n768), .ZN(new_n769));
  AND2_X1   g0569(.A1(new_n705), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(G396));
  OAI21_X1  g0571(.A(KEYINPUT104), .B1(new_n638), .B2(new_n322), .ZN(new_n772));
  INV_X1    g0572(.A(KEYINPUT104), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n325), .A2(new_n773), .A3(new_n634), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n323), .A2(new_n772), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(new_n328), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n617), .A2(new_n638), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n694), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n778), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n780), .A2(new_n612), .A3(new_n638), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n680), .B1(new_n779), .B2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(new_n703), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n680), .A2(new_n779), .A3(new_n781), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n703), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n717), .A2(new_n714), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n786), .B1(new_n202), .B2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n739), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n216), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(new_n750), .ZN(new_n791));
  OAI221_X1 g0591(.A(new_n791), .B1(new_n411), .B2(new_n745), .C1(new_n733), .C2(new_n757), .ZN(new_n792));
  OAI221_X1 g0592(.A(new_n336), .B1(new_n732), .B2(new_n551), .C1(new_n451), .C2(new_n735), .ZN(new_n793));
  INV_X1    g0593(.A(G283), .ZN(new_n794));
  OAI22_X1  g0594(.A1(new_n753), .A2(new_n564), .B1(new_n794), .B2(new_n726), .ZN(new_n795));
  NOR3_X1   g0595(.A1(new_n792), .A2(new_n793), .A3(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n732), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n736), .A2(G143), .B1(new_n797), .B2(G159), .ZN(new_n798));
  INV_X1    g0598(.A(G150), .ZN(new_n799));
  INV_X1    g0599(.A(G137), .ZN(new_n800));
  OAI221_X1 g0600(.A(new_n798), .B1(new_n799), .B2(new_n726), .C1(new_n753), .C2(new_n800), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n801), .B(KEYINPUT34), .ZN(new_n802));
  INV_X1    g0602(.A(G132), .ZN(new_n803));
  OAI22_X1  g0603(.A1(new_n757), .A2(new_n803), .B1(new_n287), .B2(new_n745), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n245), .B1(new_n789), .B2(new_n222), .ZN(new_n805));
  AOI211_X1 g0605(.A(new_n804), .B(new_n805), .C1(G58), .C2(new_n742), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n796), .B1(new_n802), .B2(new_n806), .ZN(new_n807));
  OAI221_X1 g0607(.A(new_n788), .B1(new_n765), .B2(new_n807), .C1(new_n780), .C2(new_n715), .ZN(new_n808));
  AND2_X1   g0608(.A1(new_n785), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(G384));
  INV_X1    g0610(.A(new_n498), .ZN(new_n811));
  AND2_X1   g0611(.A1(new_n811), .A2(KEYINPUT35), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n811), .A2(KEYINPUT35), .ZN(new_n813));
  NOR4_X1   g0613(.A1(new_n812), .A2(new_n813), .A3(new_n551), .A4(new_n212), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n814), .B(KEYINPUT36), .ZN(new_n815));
  OAI211_X1 g0615(.A(new_n653), .B(G77), .C1(new_n220), .C2(new_n222), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n287), .A2(G68), .ZN(new_n817));
  AOI211_X1 g0617(.A(new_n256), .B(G13), .C1(new_n816), .C2(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT40), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT38), .ZN(new_n821));
  INV_X1    g0621(.A(new_n632), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n349), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n362), .A2(new_n366), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n823), .B1(new_n824), .B2(new_n619), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n349), .A2(new_n358), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT105), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n826), .B(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT37), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n823), .A2(new_n829), .A3(new_n374), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n826), .A2(new_n823), .A3(new_n374), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n828), .A2(new_n831), .B1(KEYINPUT37), .B2(new_n832), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n821), .B1(new_n825), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n832), .A2(KEYINPUT37), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n826), .B(KEYINPUT105), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n835), .B1(new_n836), .B2(new_n830), .ZN(new_n837));
  OAI211_X1 g0637(.A(new_n837), .B(KEYINPUT38), .C1(new_n377), .C2(new_n823), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n834), .A2(KEYINPUT106), .A3(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n825), .A2(new_n833), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT106), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n840), .A2(new_n841), .A3(KEYINPUT38), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  AND2_X1   g0643(.A1(new_n677), .A2(KEYINPUT31), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n675), .B1(new_n677), .B2(new_n657), .ZN(new_n845));
  OR2_X1    g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n389), .A2(new_n634), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n404), .A2(new_n407), .A3(new_n847), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n389), .B(new_n634), .C1(new_n402), .C2(new_n403), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n778), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n846), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n820), .B1(new_n843), .B2(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n823), .B1(new_n619), .B2(new_n615), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n821), .B1(new_n853), .B2(new_n833), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n820), .B1(new_n854), .B2(new_n838), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n855), .A2(new_n846), .A3(new_n850), .ZN(new_n856));
  AND2_X1   g0656(.A1(new_n852), .A2(new_n856), .ZN(new_n857));
  AND2_X1   g0657(.A1(new_n409), .A2(new_n846), .ZN(new_n858));
  AND2_X1   g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n857), .A2(new_n858), .ZN(new_n860));
  NOR3_X1   g0660(.A1(new_n859), .A2(new_n860), .A3(new_n656), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n781), .A2(new_n777), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n848), .A2(new_n849), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  OAI22_X1  g0664(.A1(new_n864), .A2(new_n843), .B1(new_n615), .B2(new_n822), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n616), .A2(new_n638), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT39), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n854), .A2(new_n838), .A3(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n869), .B1(new_n843), .B2(new_n868), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n865), .B1(new_n867), .B2(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n693), .A2(new_n409), .A3(new_n696), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n623), .ZN(new_n873));
  XNOR2_X1  g0673(.A(new_n871), .B(new_n873), .ZN(new_n874));
  OAI22_X1  g0674(.A1(new_n861), .A2(new_n874), .B1(new_n256), .B2(new_n700), .ZN(new_n875));
  AND2_X1   g0675(.A1(new_n861), .A2(new_n874), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n819), .B1(new_n875), .B2(new_n876), .ZN(G367));
  NAND2_X1  g0677(.A1(new_n234), .A2(new_n710), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n719), .B1(new_n647), .B2(new_n522), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n786), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n540), .A2(new_n543), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n634), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(new_n545), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n883), .B1(new_n539), .B2(new_n882), .ZN(new_n884));
  AOI22_X1  g0684(.A1(G143), .A2(new_n725), .B1(new_n727), .B2(G159), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n245), .B1(new_n732), .B2(new_n287), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n886), .B1(G150), .B2(new_n736), .ZN(new_n887));
  AOI22_X1  g0687(.A1(G68), .A2(new_n742), .B1(new_n747), .B2(G137), .ZN(new_n888));
  AOI22_X1  g0688(.A1(G77), .A2(new_n739), .B1(new_n746), .B2(G58), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n885), .A2(new_n887), .A3(new_n888), .A4(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n739), .A2(G97), .ZN(new_n891));
  INV_X1    g0691(.A(G317), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n891), .B1(new_n892), .B2(new_n757), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n893), .B1(G107), .B2(new_n742), .ZN(new_n894));
  OAI221_X1 g0694(.A(new_n894), .B1(new_n451), .B2(new_n726), .C1(new_n753), .C2(new_n733), .ZN(new_n895));
  OAI221_X1 g0695(.A(new_n336), .B1(new_n732), .B2(new_n794), .C1(new_n564), .C2(new_n735), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT46), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n746), .A2(G116), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n899), .B1(new_n897), .B2(new_n898), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n890), .B1(new_n895), .B2(new_n900), .ZN(new_n901));
  XOR2_X1   g0701(.A(new_n901), .B(KEYINPUT47), .Z(new_n902));
  OAI221_X1 g0702(.A(new_n880), .B1(new_n768), .B2(new_n884), .C1(new_n902), .C2(new_n765), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n634), .A2(new_n590), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n592), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n634), .A2(new_n510), .A3(new_n506), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n637), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n908), .B(KEYINPUT107), .ZN(new_n909));
  OR2_X1    g0709(.A1(new_n909), .A2(KEYINPUT44), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(KEYINPUT44), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n637), .A2(new_n907), .ZN(new_n912));
  XOR2_X1   g0712(.A(new_n912), .B(KEYINPUT45), .Z(new_n913));
  NAND3_X1  g0713(.A1(new_n910), .A2(new_n911), .A3(new_n913), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n641), .A2(new_n645), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n914), .A2(KEYINPUT108), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(KEYINPUT108), .ZN(new_n917));
  NAND4_X1  g0717(.A1(new_n910), .A2(new_n917), .A3(new_n911), .A4(new_n913), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  MUX2_X1   g0719(.A(new_n641), .B(new_n478), .S(new_n636), .Z(new_n920));
  XNOR2_X1  g0720(.A(new_n920), .B(new_n645), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n697), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  XOR2_X1   g0722(.A(new_n651), .B(KEYINPUT41), .Z(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n702), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n478), .A2(new_n907), .A3(new_n636), .ZN(new_n926));
  OR2_X1    g0726(.A1(new_n926), .A2(KEYINPUT42), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n511), .B1(new_n905), .B2(new_n607), .ZN(new_n928));
  AOI22_X1  g0728(.A1(new_n926), .A2(KEYINPUT42), .B1(new_n638), .B2(new_n928), .ZN(new_n929));
  AOI22_X1  g0729(.A1(new_n927), .A2(new_n929), .B1(KEYINPUT43), .B2(new_n884), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n884), .A2(KEYINPUT43), .ZN(new_n931));
  XOR2_X1   g0731(.A(new_n930), .B(new_n931), .Z(new_n932));
  NAND2_X1  g0732(.A1(new_n915), .A2(new_n907), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n932), .B(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n903), .B1(new_n925), .B2(new_n934), .ZN(G387));
  AOI22_X1  g0735(.A1(new_n736), .A2(G317), .B1(new_n797), .B2(G303), .ZN(new_n936));
  INV_X1    g0736(.A(G322), .ZN(new_n937));
  OAI221_X1 g0737(.A(new_n936), .B1(new_n733), .B2(new_n726), .C1(new_n753), .C2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT48), .ZN(new_n939));
  OR2_X1    g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n938), .A2(new_n939), .ZN(new_n941));
  AOI22_X1  g0741(.A1(new_n746), .A2(G294), .B1(new_n742), .B2(G283), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT49), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n336), .B1(new_n789), .B2(new_n551), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n946), .B1(G326), .B2(new_n747), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n948), .B1(new_n944), .B2(new_n943), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n725), .A2(G159), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n950), .B(KEYINPUT109), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n726), .A2(new_n276), .ZN(new_n952));
  OAI221_X1 g0752(.A(new_n245), .B1(new_n732), .B2(new_n222), .C1(new_n287), .C2(new_n735), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n746), .A2(G77), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n747), .A2(G150), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n742), .A2(new_n522), .ZN(new_n956));
  NAND4_X1  g0756(.A1(new_n891), .A2(new_n954), .A3(new_n955), .A4(new_n956), .ZN(new_n957));
  NOR4_X1   g0757(.A1(new_n951), .A2(new_n952), .A3(new_n953), .A4(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n717), .B1(new_n949), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n231), .A2(G45), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n316), .A2(new_n287), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT50), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n513), .A2(G116), .ZN(new_n963));
  OAI211_X1 g0763(.A(new_n963), .B(new_n530), .C1(new_n222), .C2(new_n202), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n960), .B(new_n710), .C1(new_n962), .C2(new_n964), .ZN(new_n965));
  OAI221_X1 g0765(.A(new_n965), .B1(G107), .B2(new_n207), .C1(new_n963), .C2(new_n706), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n786), .B1(new_n966), .B2(new_n718), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n959), .A2(new_n967), .ZN(new_n968));
  XOR2_X1   g0768(.A(new_n968), .B(KEYINPUT110), .Z(new_n969));
  INV_X1    g0769(.A(new_n768), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n969), .B1(new_n641), .B2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n921), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n971), .B1(new_n972), .B2(new_n702), .ZN(new_n973));
  INV_X1    g0773(.A(new_n651), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n974), .B1(new_n697), .B2(new_n972), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n697), .B2(new_n972), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n973), .A2(new_n976), .ZN(G393));
  OR2_X1    g0777(.A1(new_n914), .A2(new_n915), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n914), .A2(new_n915), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n978), .A2(new_n979), .A3(new_n702), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n905), .A2(new_n716), .A3(new_n906), .ZN(new_n981));
  XOR2_X1   g0781(.A(new_n981), .B(KEYINPUT111), .Z(new_n982));
  OAI22_X1  g0782(.A1(new_n757), .A2(new_n937), .B1(new_n794), .B2(new_n745), .ZN(new_n983));
  OAI221_X1 g0783(.A(new_n336), .B1(new_n732), .B2(new_n451), .C1(new_n789), .C2(new_n411), .ZN(new_n984));
  AOI211_X1 g0784(.A(new_n983), .B(new_n984), .C1(G116), .C2(new_n742), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n564), .B2(new_n726), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n725), .A2(G317), .B1(G311), .B2(new_n736), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT52), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n725), .A2(G150), .B1(G159), .B2(new_n736), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT51), .ZN(new_n990));
  AOI211_X1 g0790(.A(new_n336), .B(new_n790), .C1(new_n316), .C2(new_n797), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n745), .A2(new_n222), .B1(new_n741), .B2(new_n202), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n992), .B1(G143), .B2(new_n747), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n991), .B(new_n993), .C1(new_n287), .C2(new_n726), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n986), .A2(new_n988), .B1(new_n990), .B2(new_n994), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT112), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(new_n717), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n718), .B1(new_n512), .B2(new_n207), .C1(new_n241), .C2(new_n711), .ZN(new_n998));
  NAND4_X1  g0798(.A1(new_n982), .A2(new_n997), .A3(new_n703), .A4(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n980), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n697), .A2(new_n972), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n919), .A2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n1002), .A2(new_n974), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n978), .A2(new_n979), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1004), .A2(new_n1001), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1000), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(G390));
  AOI21_X1  g0807(.A(new_n867), .B1(new_n862), .B2(new_n863), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n870), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n689), .A2(new_n638), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT99), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1012), .A2(new_n690), .A3(new_n777), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1013), .A2(new_n776), .A3(new_n863), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n867), .B1(new_n854), .B2(new_n838), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT113), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1014), .A2(KEYINPUT113), .A3(new_n1015), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1009), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n850), .B(G330), .C1(new_n844), .C2(new_n845), .ZN(new_n1021));
  OAI21_X1  g0821(.A(KEYINPUT114), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT114), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1021), .ZN(new_n1024));
  AND3_X1   g0824(.A1(new_n1014), .A2(KEYINPUT113), .A3(new_n1015), .ZN(new_n1025));
  AOI21_X1  g0825(.A(KEYINPUT113), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n1023), .B(new_n1024), .C1(new_n1027), .C2(new_n1009), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n680), .A2(new_n780), .A3(new_n863), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1020), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1022), .A2(new_n1028), .A3(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT115), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n409), .A2(G330), .A3(new_n846), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1032), .B1(new_n873), .B2(new_n1034), .ZN(new_n1035));
  NAND4_X1  g0835(.A1(new_n872), .A2(new_n1033), .A3(KEYINPUT115), .A4(new_n623), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n863), .B1(new_n680), .B2(new_n780), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n862), .B1(new_n1024), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1013), .A2(new_n776), .ZN(new_n1039));
  OAI211_X1 g0839(.A(G330), .B(new_n780), .C1(new_n844), .C2(new_n845), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1040), .A2(new_n848), .A3(new_n849), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1039), .A2(new_n1029), .A3(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1038), .A2(new_n1042), .ZN(new_n1043));
  AND3_X1   g0843(.A1(new_n1035), .A2(new_n1036), .A3(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1031), .A2(new_n1045), .ZN(new_n1046));
  NAND4_X1  g0846(.A1(new_n1022), .A2(new_n1028), .A3(new_n1030), .A4(new_n1044), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1046), .A2(new_n651), .A3(new_n1047), .ZN(new_n1048));
  OR2_X1    g0848(.A1(new_n870), .A2(new_n715), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n741), .A2(new_n758), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(KEYINPUT54), .B(G143), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n735), .A2(new_n803), .B1(new_n732), .B2(new_n1051), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n1050), .B(new_n1052), .C1(new_n727), .C2(G137), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n745), .A2(new_n799), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT53), .ZN(new_n1055));
  INV_X1    g0855(.A(G128), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1053), .B(new_n1055), .C1(new_n1056), .C2(new_n753), .ZN(new_n1057));
  INV_X1    g0857(.A(G125), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n245), .B1(new_n757), .B2(new_n1058), .C1(new_n789), .C2(new_n287), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT116), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n1057), .A2(new_n1060), .ZN(new_n1061));
  OR2_X1    g0861(.A1(new_n1061), .A2(KEYINPUT117), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1061), .A2(KEYINPUT117), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n789), .A2(new_n222), .B1(new_n216), .B2(new_n745), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n336), .B1(new_n732), .B2(new_n512), .C1(new_n551), .C2(new_n735), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n757), .A2(new_n451), .B1(new_n202), .B2(new_n741), .ZN(new_n1066));
  NOR3_X1   g0866(.A1(new_n1064), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n1067), .B1(new_n411), .B2(new_n726), .C1(new_n794), .C2(new_n753), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1062), .A2(new_n1063), .A3(new_n1068), .ZN(new_n1069));
  AND2_X1   g0869(.A1(new_n1069), .A2(new_n717), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n786), .B(new_n1070), .C1(new_n276), .C2(new_n787), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1049), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1072), .ZN(new_n1073));
  AND3_X1   g0873(.A1(new_n1022), .A2(new_n1028), .A3(new_n1030), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1073), .B1(new_n1074), .B2(new_n702), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1048), .A2(new_n1075), .ZN(G378));
  NAND3_X1  g0876(.A1(new_n852), .A2(G330), .A3(new_n856), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n622), .A2(new_n302), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1079), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n622), .A2(new_n302), .A3(new_n1081), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n1080), .A2(new_n292), .A3(new_n822), .A4(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n822), .A2(new_n292), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1077), .A2(new_n1083), .A3(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1086), .A2(new_n1083), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n1088), .A2(G330), .A3(new_n852), .A4(new_n856), .ZN(new_n1089));
  AND3_X1   g0889(.A1(new_n1087), .A2(new_n1089), .A3(new_n871), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n871), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n1088), .A2(new_n715), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n245), .A2(G41), .ZN(new_n1094));
  AOI211_X1 g0894(.A(G50), .B(new_n1094), .C1(new_n417), .C2(new_n441), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n739), .A2(G58), .ZN(new_n1096));
  XOR2_X1   g0896(.A(new_n1096), .B(KEYINPUT118), .Z(new_n1097));
  OAI221_X1 g0897(.A(new_n1097), .B1(new_n512), .B2(new_n726), .C1(new_n551), .C2(new_n753), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n1094), .B1(new_n314), .B2(new_n732), .C1(new_n411), .C2(new_n735), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n954), .B1(new_n222), .B2(new_n741), .C1(new_n794), .C2(new_n757), .ZN(new_n1100));
  NOR3_X1   g0900(.A1(new_n1098), .A2(new_n1099), .A3(new_n1100), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(KEYINPUT119), .B(KEYINPUT58), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1095), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n735), .A2(new_n1056), .B1(new_n732), .B2(new_n800), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n745), .A2(new_n1051), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n1105), .B(new_n1106), .C1(G150), .C2(new_n742), .ZN(new_n1107));
  OAI221_X1 g0907(.A(new_n1107), .B1(new_n803), .B2(new_n726), .C1(new_n1058), .C2(new_n753), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n1108), .A2(KEYINPUT59), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1108), .A2(KEYINPUT59), .ZN(new_n1110));
  AOI211_X1 g0910(.A(G33), .B(G41), .C1(new_n747), .C2(G124), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1111), .B1(new_n758), .B2(new_n789), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT120), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1110), .A2(new_n1113), .ZN(new_n1114));
  OAI221_X1 g0914(.A(new_n1104), .B1(new_n1109), .B2(new_n1114), .C1(new_n1103), .C2(new_n1101), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(new_n717), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n787), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1116), .B(new_n703), .C1(G50), .C2(new_n1117), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n1092), .A2(new_n701), .B1(new_n1093), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1092), .B1(new_n1047), .B2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n651), .B1(new_n1123), .B2(KEYINPUT57), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT57), .ZN(new_n1125));
  AOI211_X1 g0925(.A(new_n1125), .B(new_n1092), .C1(new_n1047), .C2(new_n1122), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1120), .B1(new_n1124), .B2(new_n1126), .ZN(G375));
  INV_X1    g0927(.A(new_n1043), .ZN(new_n1128));
  AOI21_X1  g0928(.A(KEYINPUT122), .B1(new_n1121), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT122), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n1130), .B(new_n1043), .C1(new_n1035), .C2(new_n1036), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n923), .B(KEYINPUT121), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1044), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1043), .A2(new_n702), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT123), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(new_n1136), .B(new_n1137), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n703), .B1(G68), .B2(new_n1117), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n956), .B1(new_n789), .B2(new_n202), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n757), .A2(new_n564), .B1(new_n512), .B2(new_n745), .ZN(new_n1141));
  OAI221_X1 g0941(.A(new_n336), .B1(new_n732), .B2(new_n411), .C1(new_n794), .C2(new_n735), .ZN(new_n1142));
  NOR3_X1   g0942(.A1(new_n1140), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  OAI221_X1 g0943(.A(new_n1143), .B1(new_n551), .B2(new_n726), .C1(new_n451), .C2(new_n753), .ZN(new_n1144));
  OAI221_X1 g0944(.A(new_n1097), .B1(new_n803), .B2(new_n753), .C1(new_n726), .C2(new_n1051), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n746), .A2(G159), .B1(new_n742), .B2(G50), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n245), .B1(new_n732), .B2(new_n799), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1147), .B1(G137), .B2(new_n736), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1146), .B(new_n1148), .C1(new_n1056), .C2(new_n757), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1144), .B1(new_n1145), .B2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1139), .B1(new_n1150), .B2(new_n717), .ZN(new_n1151));
  XOR2_X1   g0951(.A(new_n1151), .B(KEYINPUT124), .Z(new_n1152));
  OAI21_X1  g0952(.A(new_n1152), .B1(new_n863), .B2(new_n715), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1138), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1135), .A2(new_n1155), .ZN(G381));
  NOR2_X1   g0956(.A1(G393), .A2(G396), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(new_n809), .ZN(new_n1158));
  XOR2_X1   g0958(.A(new_n1158), .B(KEYINPUT125), .Z(new_n1159));
  OR2_X1    g0959(.A1(new_n925), .A2(new_n934), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1160), .A2(new_n903), .A3(new_n1006), .ZN(new_n1161));
  NOR3_X1   g0961(.A1(new_n1159), .A2(G381), .A3(new_n1161), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1072), .B1(new_n1031), .B2(new_n701), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n974), .B1(new_n1031), .B2(new_n1045), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1163), .B1(new_n1047), .B2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(G375), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1162), .A2(new_n1165), .A3(new_n1166), .ZN(G407));
  NOR2_X1   g0967(.A1(new_n628), .A2(G343), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1166), .A2(new_n1165), .A3(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(G407), .A2(new_n1169), .A3(G213), .ZN(G409));
  XOR2_X1   g0970(.A(KEYINPUT127), .B(KEYINPUT61), .Z(new_n1171));
  AOI21_X1  g0971(.A(new_n770), .B1(new_n973), .B2(new_n976), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1157), .A2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1006), .B1(new_n1160), .B2(new_n903), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(G390), .A2(G387), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1173), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(G390), .A2(G387), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n1161), .B(new_n1177), .C1(new_n1157), .C2(new_n1172), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1171), .B1(new_n1176), .B2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1168), .A2(G2897), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1121), .A2(new_n1128), .A3(KEYINPUT60), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(new_n651), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1045), .A2(KEYINPUT60), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1182), .B1(new_n1132), .B2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n809), .B1(new_n1184), .B2(new_n1154), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT60), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1044), .A2(new_n1186), .ZN(new_n1187));
  NOR3_X1   g0987(.A1(new_n1187), .A2(new_n1129), .A3(new_n1131), .ZN(new_n1188));
  OAI211_X1 g0988(.A(G384), .B(new_n1155), .C1(new_n1188), .C2(new_n1182), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1180), .B1(new_n1185), .B2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1185), .A2(new_n1189), .A3(new_n1180), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  OAI211_X1 g0993(.A(G378), .B(new_n1120), .C1(new_n1124), .C2(new_n1126), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n1133), .B(new_n1092), .C1(new_n1047), .C2(new_n1122), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1165), .B1(new_n1119), .B2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1168), .B1(new_n1194), .B2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1179), .B1(new_n1193), .B2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1185), .A2(new_n1189), .ZN(new_n1199));
  AOI211_X1 g0999(.A(new_n1168), .B(new_n1199), .C1(new_n1194), .C2(new_n1196), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1200), .A2(KEYINPUT62), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1199), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1168), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1202), .A2(new_n1203), .A3(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(KEYINPUT62), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1198), .B1(new_n1201), .B2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT126), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n1200), .B2(KEYINPUT63), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT63), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1205), .A2(KEYINPUT126), .A3(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1200), .A2(KEYINPUT63), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1202), .A2(new_n1204), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1192), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1215), .A2(new_n1190), .ZN(new_n1216));
  AOI21_X1  g1016(.A(KEYINPUT61), .B1(new_n1214), .B2(new_n1216), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n1210), .A2(new_n1212), .A3(new_n1213), .A4(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1176), .A2(new_n1178), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1208), .B1(new_n1218), .B2(new_n1220), .ZN(G405));
  NAND2_X1  g1021(.A1(G375), .A2(new_n1165), .ZN(new_n1222));
  AND3_X1   g1022(.A1(new_n1222), .A2(new_n1194), .A3(new_n1199), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1199), .B1(new_n1222), .B2(new_n1194), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  XNOR2_X1  g1025(.A(new_n1225), .B(new_n1220), .ZN(G402));
endmodule


