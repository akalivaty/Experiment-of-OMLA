//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 1 0 0 1 1 1 1 0 1 0 1 1 1 0 1 0 1 0 0 1 0 0 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 1 1 1 0 0 1 0 0 0 0 0 0 1 0 0 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:58 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n449, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n491, new_n492, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n508, new_n509, new_n510, new_n511, new_n512,
    new_n513, new_n514, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n522, new_n523, new_n524, new_n525, new_n526, new_n527, new_n530,
    new_n531, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n546, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n590, new_n591, new_n594, new_n596, new_n597, new_n598,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  INV_X1    g022(.A(G567), .ZN(new_n448));
  NOR2_X1   g023(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT64), .Z(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G2106), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n453), .A2(new_n457), .B1(new_n448), .B2(new_n454), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT65), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G125), .ZN(new_n462));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(new_n460), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  AND3_X1   g039(.A1(KEYINPUT66), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(KEYINPUT3), .B1(KEYINPUT66), .B2(G2104), .ZN(new_n466));
  OAI21_X1  g041(.A(G137), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(G101), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(G2105), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n464), .A2(new_n469), .ZN(G160));
  NOR2_X1   g045(.A1(new_n465), .A2(new_n466), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G136), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n471), .A2(new_n460), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G124), .ZN(new_n475));
  NOR2_X1   g050(.A1(G100), .A2(G2105), .ZN(new_n476));
  OAI21_X1  g051(.A(G2104), .B1(new_n460), .B2(G112), .ZN(new_n477));
  OAI211_X1 g052(.A(new_n473), .B(new_n475), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  XOR2_X1   g053(.A(new_n478), .B(KEYINPUT67), .Z(G162));
  NAND2_X1  g054(.A1(KEYINPUT4), .A2(G138), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n481), .B1(new_n465), .B2(new_n466), .ZN(new_n482));
  NAND2_X1  g057(.A1(G102), .A2(G2104), .ZN(new_n483));
  AOI21_X1  g058(.A(G2105), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  OAI21_X1  g059(.A(G126), .B1(new_n465), .B2(new_n466), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT4), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n486), .B1(G114), .B2(G2104), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n460), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  AOI21_X1  g063(.A(KEYINPUT4), .B1(new_n461), .B2(G138), .ZN(new_n489));
  NOR3_X1   g064(.A1(new_n484), .A2(new_n488), .A3(new_n489), .ZN(G164));
  INV_X1    g065(.A(G651), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT6), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT6), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G651), .ZN(new_n494));
  AND2_X1   g069(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G543), .ZN(new_n496));
  INV_X1    g071(.A(G50), .ZN(new_n497));
  OR2_X1    g072(.A1(KEYINPUT5), .A2(G543), .ZN(new_n498));
  NAND2_X1  g073(.A1(KEYINPUT5), .A2(G543), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n500), .A2(new_n492), .A3(new_n494), .ZN(new_n501));
  INV_X1    g076(.A(G88), .ZN(new_n502));
  OAI22_X1  g077(.A1(new_n496), .A2(new_n497), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n500), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n504), .A2(new_n491), .ZN(new_n505));
  OR2_X1    g080(.A1(new_n503), .A2(new_n505), .ZN(G303));
  INV_X1    g081(.A(G303), .ZN(G166));
  NAND3_X1  g082(.A1(new_n500), .A2(G63), .A3(G651), .ZN(new_n508));
  INV_X1    g083(.A(G51), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n508), .B1(new_n496), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g085(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n511));
  XNOR2_X1  g086(.A(new_n511), .B(KEYINPUT7), .ZN(new_n512));
  INV_X1    g087(.A(G89), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n512), .B1(new_n501), .B2(new_n513), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n510), .A2(new_n514), .ZN(G168));
  INV_X1    g090(.A(G52), .ZN(new_n516));
  INV_X1    g091(.A(G90), .ZN(new_n517));
  OAI22_X1  g092(.A1(new_n496), .A2(new_n516), .B1(new_n501), .B2(new_n517), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n500), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n519), .A2(new_n491), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n518), .A2(new_n520), .ZN(G171));
  INV_X1    g096(.A(G43), .ZN(new_n522));
  INV_X1    g097(.A(G81), .ZN(new_n523));
  OAI22_X1  g098(.A1(new_n496), .A2(new_n522), .B1(new_n501), .B2(new_n523), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n500), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n525), .A2(new_n491), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G860), .ZN(G153));
  NAND4_X1  g103(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g104(.A1(G1), .A2(G3), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT8), .ZN(new_n531));
  NAND4_X1  g106(.A1(G319), .A2(G483), .A3(G661), .A4(new_n531), .ZN(G188));
  INV_X1    g107(.A(new_n496), .ZN(new_n533));
  INV_X1    g108(.A(G53), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n534), .B1(KEYINPUT68), .B2(KEYINPUT9), .ZN(new_n535));
  OAI211_X1 g110(.A(new_n533), .B(new_n535), .C1(KEYINPUT68), .C2(KEYINPUT9), .ZN(new_n536));
  XNOR2_X1  g111(.A(KEYINPUT69), .B(G65), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n500), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(G78), .A2(G543), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G651), .ZN(new_n541));
  INV_X1    g116(.A(new_n501), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G91), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT68), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT9), .ZN(new_n545));
  OAI211_X1 g120(.A(new_n544), .B(new_n545), .C1(new_n496), .C2(new_n534), .ZN(new_n546));
  NAND4_X1  g121(.A1(new_n536), .A2(new_n541), .A3(new_n543), .A4(new_n546), .ZN(G299));
  OR2_X1    g122(.A1(new_n518), .A2(new_n520), .ZN(G301));
  INV_X1    g123(.A(G168), .ZN(G286));
  NAND3_X1  g124(.A1(new_n495), .A2(G49), .A3(G543), .ZN(new_n550));
  OAI21_X1  g125(.A(G651), .B1(new_n500), .B2(G74), .ZN(new_n551));
  AND2_X1   g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT70), .ZN(new_n553));
  AND3_X1   g128(.A1(new_n495), .A2(G87), .A3(new_n500), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n552), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n550), .A2(new_n551), .ZN(new_n557));
  OAI21_X1  g132(.A(KEYINPUT70), .B1(new_n557), .B2(new_n554), .ZN(new_n558));
  AND2_X1   g133(.A1(new_n556), .A2(new_n558), .ZN(G288));
  INV_X1    g134(.A(G61), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n560), .B1(new_n498), .B2(new_n499), .ZN(new_n561));
  NAND2_X1  g136(.A1(G73), .A2(G543), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(new_n563));
  OAI21_X1  g138(.A(G651), .B1(new_n561), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n495), .A2(G86), .A3(new_n500), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n495), .A2(G48), .A3(G543), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(G305));
  INV_X1    g142(.A(G47), .ZN(new_n568));
  INV_X1    g143(.A(G85), .ZN(new_n569));
  OAI22_X1  g144(.A1(new_n496), .A2(new_n568), .B1(new_n501), .B2(new_n569), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n500), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n571), .A2(new_n491), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(G290));
  INV_X1    g149(.A(G868), .ZN(new_n575));
  NOR2_X1   g150(.A1(G301), .A2(new_n575), .ZN(new_n576));
  AND3_X1   g151(.A1(new_n495), .A2(G92), .A3(new_n500), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n577), .B(KEYINPUT10), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n500), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n579));
  OR2_X1    g154(.A1(new_n579), .A2(new_n491), .ZN(new_n580));
  INV_X1    g155(.A(G54), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT71), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n581), .B1(new_n496), .B2(new_n582), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n583), .B1(new_n582), .B2(new_n496), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n578), .A2(new_n580), .A3(new_n584), .ZN(new_n585));
  XNOR2_X1  g160(.A(new_n585), .B(KEYINPUT72), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n576), .B1(new_n587), .B2(new_n575), .ZN(G284));
  AOI21_X1  g163(.A(new_n576), .B1(new_n587), .B2(new_n575), .ZN(G321));
  NAND2_X1  g164(.A1(G286), .A2(G868), .ZN(new_n590));
  INV_X1    g165(.A(G299), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n591), .B2(G868), .ZN(G297));
  XNOR2_X1  g167(.A(G297), .B(KEYINPUT73), .ZN(G280));
  INV_X1    g168(.A(G559), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n587), .B1(new_n594), .B2(G860), .ZN(G148));
  INV_X1    g170(.A(new_n527), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n596), .A2(new_n575), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n586), .A2(G559), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n598), .B2(new_n575), .ZN(G323));
  XNOR2_X1  g174(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g175(.A1(new_n472), .A2(G135), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n601), .B(KEYINPUT74), .ZN(new_n602));
  OR2_X1    g177(.A1(G99), .A2(G2105), .ZN(new_n603));
  INV_X1    g178(.A(G2104), .ZN(new_n604));
  INV_X1    g179(.A(G111), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n604), .B1(new_n605), .B2(G2105), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n474), .A2(G123), .B1(new_n603), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n602), .A2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(G2096), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n608), .B(new_n609), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n460), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT12), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT13), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(G2100), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n610), .A2(new_n614), .ZN(G156));
  XNOR2_X1  g190(.A(G2443), .B(G2446), .ZN(new_n616));
  XNOR2_X1  g191(.A(G2451), .B(G2454), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n616), .B(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(new_n618), .ZN(new_n619));
  XNOR2_X1  g194(.A(G2427), .B(G2438), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(G2430), .ZN(new_n621));
  XNOR2_X1  g196(.A(KEYINPUT15), .B(G2435), .ZN(new_n622));
  OR2_X1    g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n621), .A2(new_n622), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n623), .A2(KEYINPUT14), .A3(new_n624), .ZN(new_n625));
  XNOR2_X1  g200(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g202(.A(new_n627), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n625), .A2(new_n626), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n619), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n625), .A2(new_n626), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n631), .A2(new_n618), .A3(new_n627), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(G1341), .B(G1348), .ZN(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(new_n635));
  OAI21_X1  g210(.A(G14), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  NOR3_X1   g211(.A1(new_n628), .A2(new_n629), .A3(new_n619), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n618), .B1(new_n631), .B2(new_n627), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n635), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  INV_X1    g214(.A(KEYINPUT76), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n633), .A2(KEYINPUT76), .A3(new_n635), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n636), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT77), .ZN(G401));
  XNOR2_X1  g219(.A(G2072), .B(G2078), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2067), .B(G2678), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g222(.A(KEYINPUT78), .ZN(new_n648));
  XOR2_X1   g223(.A(G2084), .B(G2090), .Z(new_n649));
  OR3_X1    g224(.A1(new_n647), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n648), .B1(new_n647), .B2(new_n649), .ZN(new_n651));
  INV_X1    g226(.A(new_n646), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n645), .B(KEYINPUT17), .Z(new_n653));
  OAI211_X1 g228(.A(new_n650), .B(new_n651), .C1(new_n652), .C2(new_n653), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n649), .A2(new_n645), .A3(new_n646), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n655), .B(KEYINPUT18), .Z(new_n656));
  NAND3_X1  g231(.A1(new_n653), .A2(new_n649), .A3(new_n652), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n654), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(new_n609), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n659), .A2(G2100), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(G2100), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(G227));
  XOR2_X1   g237(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n663));
  XNOR2_X1  g238(.A(G1971), .B(G1976), .ZN(new_n664));
  INV_X1    g239(.A(KEYINPUT79), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT19), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1956), .B(G2474), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1961), .B(G1966), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(KEYINPUT20), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n668), .B(new_n669), .ZN(new_n674));
  OR2_X1    g249(.A1(new_n667), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NOR3_X1   g252(.A1(new_n673), .A2(G1986), .A3(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(G1986), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n671), .B(KEYINPUT20), .ZN(new_n680));
  INV_X1    g255(.A(new_n677), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n679), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n663), .B1(new_n678), .B2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1991), .B(G1996), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT80), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(G1981), .ZN(new_n686));
  OAI21_X1  g261(.A(G1986), .B1(new_n673), .B2(new_n677), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n680), .A2(new_n681), .A3(new_n679), .ZN(new_n688));
  INV_X1    g263(.A(new_n663), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n687), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  AND3_X1   g265(.A1(new_n683), .A2(new_n686), .A3(new_n690), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n686), .B1(new_n683), .B2(new_n690), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(G229));
  INV_X1    g269(.A(G29), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(G25), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n474), .A2(G119), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT81), .ZN(new_n698));
  OR2_X1    g273(.A1(G95), .A2(G2105), .ZN(new_n699));
  INV_X1    g274(.A(G107), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n604), .B1(new_n700), .B2(G2105), .ZN(new_n701));
  AOI22_X1  g276(.A1(new_n472), .A2(G131), .B1(new_n699), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n698), .A2(new_n702), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT82), .Z(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n696), .B1(new_n705), .B2(new_n695), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT83), .ZN(new_n707));
  XOR2_X1   g282(.A(KEYINPUT35), .B(G1991), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  MUX2_X1   g284(.A(G6), .B(G305), .S(G16), .Z(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT32), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n711), .A2(G1981), .ZN(new_n712));
  INV_X1    g287(.A(G16), .ZN(new_n713));
  AND2_X1   g288(.A1(new_n713), .A2(G23), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n552), .A2(new_n555), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n714), .B1(new_n715), .B2(G16), .ZN(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT33), .B(G1976), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(G303), .A2(G16), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n713), .A2(G22), .ZN(new_n720));
  AND2_X1   g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n718), .B1(new_n722), .B2(G1971), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n711), .A2(G1981), .ZN(new_n724));
  INV_X1    g299(.A(G1971), .ZN(new_n725));
  AOI22_X1  g300(.A1(new_n721), .A2(new_n725), .B1(new_n716), .B2(new_n717), .ZN(new_n726));
  NAND4_X1  g301(.A1(new_n712), .A2(new_n723), .A3(new_n724), .A4(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(KEYINPUT34), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n727), .A2(KEYINPUT34), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n713), .A2(G24), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(new_n573), .B2(new_n713), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(G1986), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n729), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n709), .A2(new_n728), .A3(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT36), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n735), .A2(KEYINPUT84), .ZN(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n735), .A2(KEYINPUT84), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n734), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  NAND4_X1  g314(.A1(new_n709), .A2(new_n728), .A3(new_n733), .A4(new_n736), .ZN(new_n740));
  NOR2_X1   g315(.A1(G4), .A2(G16), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(new_n587), .B2(G16), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(G1348), .Z(new_n743));
  OAI21_X1  g318(.A(new_n695), .B1(KEYINPUT24), .B2(G34), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(KEYINPUT24), .B2(G34), .ZN(new_n745));
  INV_X1    g320(.A(G160), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n745), .B1(new_n746), .B2(G29), .ZN(new_n747));
  INV_X1    g322(.A(G2084), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT87), .Z(new_n750));
  NAND2_X1  g325(.A1(new_n695), .A2(G33), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n472), .A2(G139), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT25), .Z(new_n754));
  AOI22_X1  g329(.A1(new_n461), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n755));
  OAI211_X1 g330(.A(new_n752), .B(new_n754), .C1(new_n460), .C2(new_n755), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT86), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n751), .B1(new_n757), .B2(new_n695), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n750), .B1(new_n758), .B2(G2072), .ZN(new_n759));
  OAI211_X1 g334(.A(new_n743), .B(new_n759), .C1(G2072), .C2(new_n758), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n713), .A2(G20), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT23), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(new_n591), .B2(new_n713), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(G1956), .ZN(new_n764));
  NOR2_X1   g339(.A1(G27), .A2(G29), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(G164), .B2(G29), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n764), .B1(G2078), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n472), .A2(G140), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n474), .A2(G128), .ZN(new_n769));
  NOR2_X1   g344(.A1(G104), .A2(G2105), .ZN(new_n770));
  OAI21_X1  g345(.A(G2104), .B1(new_n460), .B2(G116), .ZN(new_n771));
  OAI211_X1 g346(.A(new_n768), .B(new_n769), .C1(new_n770), .C2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n772), .A2(G29), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n695), .A2(G26), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT28), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  XOR2_X1   g351(.A(KEYINPUT85), .B(G2067), .Z(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n713), .A2(G21), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G168), .B2(new_n713), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n780), .A2(G1966), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT90), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n767), .A2(new_n778), .A3(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(new_n608), .ZN(new_n784));
  AOI22_X1  g359(.A1(new_n784), .A2(G29), .B1(G1966), .B2(new_n780), .ZN(new_n785));
  INV_X1    g360(.A(G1961), .ZN(new_n786));
  NOR2_X1   g361(.A1(G171), .A2(new_n713), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(G5), .B2(new_n713), .ZN(new_n788));
  OAI221_X1 g363(.A(new_n785), .B1(new_n786), .B2(new_n788), .C1(G2078), .C2(new_n766), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n713), .A2(G19), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(new_n527), .B2(new_n713), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(G1341), .Z(new_n792));
  INV_X1    g367(.A(KEYINPUT30), .ZN(new_n793));
  AND2_X1   g368(.A1(new_n793), .A2(G28), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n695), .B1(new_n793), .B2(G28), .ZN(new_n795));
  AND2_X1   g370(.A1(KEYINPUT31), .A2(G11), .ZN(new_n796));
  NOR2_X1   g371(.A1(KEYINPUT31), .A2(G11), .ZN(new_n797));
  OAI22_X1  g372(.A1(new_n794), .A2(new_n795), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(new_n788), .B2(new_n786), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n747), .A2(new_n748), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n792), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n789), .A2(new_n801), .ZN(new_n802));
  XOR2_X1   g377(.A(KEYINPUT88), .B(KEYINPUT26), .Z(new_n803));
  NAND3_X1  g378(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n472), .A2(G141), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n474), .A2(G129), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n460), .A2(G105), .A3(G2104), .ZN(new_n808));
  NAND4_X1  g383(.A1(new_n805), .A2(new_n806), .A3(new_n807), .A4(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT89), .ZN(new_n810));
  OR2_X1    g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n809), .A2(new_n810), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  MUX2_X1   g388(.A(G32), .B(new_n813), .S(G29), .Z(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT27), .B(G1996), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n695), .A2(G35), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(G162), .B2(new_n695), .ZN(new_n818));
  XOR2_X1   g393(.A(KEYINPUT29), .B(G2090), .Z(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n816), .A2(new_n820), .ZN(new_n821));
  NOR4_X1   g396(.A1(new_n760), .A2(new_n783), .A3(new_n802), .A4(new_n821), .ZN(new_n822));
  AND3_X1   g397(.A1(new_n739), .A2(new_n740), .A3(new_n822), .ZN(G311));
  NAND3_X1  g398(.A1(new_n739), .A2(new_n740), .A3(new_n822), .ZN(G150));
  NAND2_X1  g399(.A1(new_n587), .A2(G559), .ZN(new_n825));
  XNOR2_X1  g400(.A(KEYINPUT91), .B(KEYINPUT38), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n500), .A2(G67), .ZN(new_n828));
  NAND2_X1  g403(.A1(G80), .A2(G543), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT92), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n491), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(new_n831), .B2(new_n830), .ZN(new_n833));
  INV_X1    g408(.A(G55), .ZN(new_n834));
  XNOR2_X1  g409(.A(KEYINPUT93), .B(G93), .ZN(new_n835));
  OAI22_X1  g410(.A1(new_n496), .A2(new_n834), .B1(new_n501), .B2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n833), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(new_n596), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n833), .A2(new_n527), .A3(new_n837), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n827), .B(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT39), .ZN(new_n843));
  AOI21_X1  g418(.A(G860), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n844), .B1(new_n843), .B2(new_n842), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n838), .A2(G860), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n846), .B(KEYINPUT37), .Z(new_n847));
  NAND2_X1  g422(.A1(new_n845), .A2(new_n847), .ZN(G145));
  INV_X1    g423(.A(KEYINPUT96), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n472), .A2(G142), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n474), .A2(G130), .ZN(new_n851));
  OR2_X1    g426(.A1(G106), .A2(G2105), .ZN(new_n852));
  OAI211_X1 g427(.A(new_n852), .B(G2104), .C1(G118), .C2(new_n460), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n850), .A2(new_n851), .A3(new_n853), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n698), .A2(new_n612), .A3(new_n702), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n612), .B1(new_n698), .B2(new_n702), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n854), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n857), .ZN(new_n859));
  INV_X1    g434(.A(new_n854), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n859), .A2(new_n860), .A3(new_n855), .ZN(new_n861));
  AND3_X1   g436(.A1(new_n858), .A2(new_n861), .A3(KEYINPUT95), .ZN(new_n862));
  AOI21_X1  g437(.A(KEYINPUT95), .B1(new_n858), .B2(new_n861), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n772), .B(G164), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n813), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n485), .A2(new_n487), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n867), .A2(G2105), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n482), .A2(new_n483), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(new_n460), .ZN(new_n870));
  INV_X1    g445(.A(new_n489), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n868), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n772), .B(new_n872), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n873), .A2(new_n812), .A3(new_n811), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n866), .A2(new_n874), .A3(new_n756), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(KEYINPUT94), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT94), .ZN(new_n877));
  NAND4_X1  g452(.A1(new_n866), .A2(new_n874), .A3(new_n877), .A4(new_n756), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n866), .A2(new_n874), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n879), .A2(new_n757), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n876), .A2(new_n878), .A3(new_n880), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n849), .B1(new_n864), .B2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT95), .ZN(new_n883));
  INV_X1    g458(.A(new_n861), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n860), .B1(new_n859), .B2(new_n855), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n883), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n858), .A2(new_n861), .A3(KEYINPUT95), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AOI22_X1  g463(.A1(new_n875), .A2(KEYINPUT94), .B1(new_n879), .B2(new_n757), .ZN(new_n889));
  NAND4_X1  g464(.A1(new_n888), .A2(new_n889), .A3(KEYINPUT96), .A4(new_n878), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n882), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n864), .A2(new_n881), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n608), .B(G160), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(G162), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n884), .A2(new_n885), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n895), .B1(new_n881), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(G37), .B1(new_n891), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n896), .A2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g476(.A1(new_n838), .A2(new_n575), .ZN(new_n902));
  AND2_X1   g477(.A1(new_n839), .A2(new_n840), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n598), .B(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n591), .A2(new_n585), .ZN(new_n905));
  NAND4_X1  g480(.A1(G299), .A2(new_n578), .A3(new_n580), .A4(new_n584), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n904), .ZN(new_n909));
  XOR2_X1   g484(.A(KEYINPUT98), .B(KEYINPUT41), .Z(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n905), .A2(new_n906), .A3(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n907), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n912), .B1(new_n913), .B2(KEYINPUT41), .ZN(new_n914));
  AOI22_X1  g489(.A1(new_n908), .A2(KEYINPUT97), .B1(new_n909), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n915), .B1(KEYINPUT97), .B2(new_n908), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n573), .B(new_n715), .ZN(new_n917));
  AND2_X1   g492(.A1(new_n917), .A2(KEYINPUT99), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n917), .A2(KEYINPUT99), .ZN(new_n919));
  XNOR2_X1  g494(.A(G303), .B(G305), .ZN(new_n920));
  OR3_X1    g495(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n920), .A2(KEYINPUT99), .A3(new_n917), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n923), .B(KEYINPUT42), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n916), .B(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n902), .B1(new_n925), .B2(new_n575), .ZN(G295));
  OAI21_X1  g501(.A(new_n902), .B1(new_n925), .B2(new_n575), .ZN(G331));
  INV_X1    g502(.A(KEYINPUT100), .ZN(new_n928));
  NAND2_X1  g503(.A1(G301), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(G171), .A2(KEYINPUT100), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n929), .A2(G286), .A3(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(G171), .A2(G168), .A3(KEYINPUT100), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n931), .A2(new_n839), .A3(new_n840), .A4(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  AOI22_X1  g509(.A1(new_n931), .A2(new_n932), .B1(new_n839), .B2(new_n840), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n905), .A2(new_n906), .A3(new_n911), .ZN(new_n936));
  AOI21_X1  g511(.A(KEYINPUT41), .B1(new_n905), .B2(new_n906), .ZN(new_n937));
  OAI22_X1  g512(.A1(new_n934), .A2(new_n935), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(KEYINPUT101), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n931), .A2(new_n932), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(new_n841), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(new_n933), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT101), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n914), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n933), .B(KEYINPUT102), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n913), .A2(new_n935), .ZN(new_n946));
  AOI22_X1  g521(.A1(new_n939), .A2(new_n944), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(G37), .B1(new_n947), .B2(new_n923), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT43), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n945), .A2(new_n946), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n938), .A2(KEYINPUT101), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n943), .B1(new_n914), .B2(new_n942), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n950), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n923), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n948), .A2(new_n949), .A3(new_n955), .ZN(new_n956));
  OR2_X1    g531(.A1(new_n956), .A2(KEYINPUT104), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n907), .A2(KEYINPUT41), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n958), .B1(new_n907), .B2(new_n911), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n903), .A2(KEYINPUT102), .A3(new_n932), .A4(new_n931), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT102), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n933), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n960), .A2(new_n941), .A3(new_n962), .ZN(new_n963));
  AOI22_X1  g538(.A1(new_n959), .A2(new_n963), .B1(new_n933), .B2(new_n946), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT103), .ZN(new_n965));
  OR3_X1    g540(.A1(new_n964), .A2(new_n965), .A3(new_n923), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n965), .B1(new_n964), .B2(new_n923), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n948), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(KEYINPUT43), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n956), .A2(KEYINPUT104), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n957), .A2(KEYINPUT44), .A3(new_n969), .A4(new_n970), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n948), .A2(new_n966), .A3(new_n949), .A4(new_n967), .ZN(new_n972));
  INV_X1    g547(.A(G37), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n973), .B1(new_n953), .B2(new_n954), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n947), .A2(new_n923), .ZN(new_n975));
  OAI21_X1  g550(.A(KEYINPUT43), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n972), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n971), .B1(new_n978), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g554(.A(KEYINPUT45), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n980), .B1(G164), .B2(G1384), .ZN(new_n981));
  XNOR2_X1  g556(.A(KEYINPUT105), .B(G40), .ZN(new_n982));
  NOR3_X1   g557(.A1(new_n464), .A2(new_n469), .A3(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n981), .A2(new_n984), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n772), .B(G2067), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  XOR2_X1   g562(.A(new_n987), .B(KEYINPUT106), .Z(new_n988));
  XNOR2_X1  g563(.A(new_n813), .B(G1996), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n988), .B1(new_n985), .B2(new_n989), .ZN(new_n990));
  XOR2_X1   g565(.A(new_n703), .B(new_n708), .Z(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(new_n985), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n573), .B(new_n679), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n993), .B1(new_n985), .B2(new_n994), .ZN(new_n995));
  XNOR2_X1  g570(.A(KEYINPUT110), .B(G8), .ZN(new_n996));
  NOR2_X1   g571(.A1(G168), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n489), .B1(new_n869), .B2(new_n460), .ZN(new_n999));
  AOI21_X1  g574(.A(G1384), .B1(new_n999), .B2(new_n868), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT50), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n983), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NOR3_X1   g577(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1000), .A2(KEYINPUT45), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1005), .A2(new_n981), .A3(new_n983), .ZN(new_n1006));
  INV_X1    g581(.A(G1966), .ZN(new_n1007));
  AOI22_X1  g582(.A1(new_n1004), .A2(new_n748), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(G8), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n998), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NOR3_X1   g585(.A1(G164), .A2(new_n980), .A3(G1384), .ZN(new_n1011));
  INV_X1    g586(.A(G1384), .ZN(new_n1012));
  AOI21_X1  g587(.A(KEYINPUT45), .B1(new_n872), .B2(new_n1012), .ZN(new_n1013));
  NOR3_X1   g588(.A1(new_n1011), .A2(new_n1013), .A3(new_n984), .ZN(new_n1014));
  OAI21_X1  g589(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n872), .A2(new_n1001), .A3(new_n1012), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1015), .A2(new_n983), .A3(new_n1016), .ZN(new_n1017));
  OAI22_X1  g592(.A1(new_n1014), .A2(G1966), .B1(G2084), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(new_n996), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n997), .A2(KEYINPUT51), .ZN(new_n1021));
  AOI22_X1  g596(.A1(new_n1010), .A2(KEYINPUT51), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT121), .ZN(new_n1023));
  NOR3_X1   g598(.A1(new_n1008), .A2(new_n1023), .A3(new_n998), .ZN(new_n1024));
  AOI21_X1  g599(.A(KEYINPUT121), .B1(new_n1018), .B2(new_n997), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(KEYINPUT62), .B1(new_n1022), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT108), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT107), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1029), .B1(new_n1005), .B2(new_n981), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n983), .B1(new_n1013), .B2(KEYINPUT107), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1028), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(KEYINPUT107), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n984), .B1(new_n981), .B2(new_n1029), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1033), .A2(new_n1034), .A3(KEYINPUT108), .ZN(new_n1035));
  AOI21_X1  g610(.A(G2078), .B1(new_n1032), .B2(new_n1035), .ZN(new_n1036));
  OR2_X1    g611(.A1(new_n1036), .A2(KEYINPUT53), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT119), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1017), .A2(new_n1038), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1015), .A2(KEYINPUT119), .A3(new_n1016), .A4(new_n983), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT53), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1042), .A2(G2078), .ZN(new_n1043));
  AOI22_X1  g618(.A1(new_n1041), .A2(new_n786), .B1(new_n1014), .B2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(G301), .B1(new_n1037), .B2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n997), .B1(new_n1018), .B2(G8), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT51), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1008), .A2(new_n996), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1021), .ZN(new_n1049));
  OAI22_X1  g624(.A1(new_n1046), .A2(new_n1047), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT62), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1023), .B1(new_n1008), .B2(new_n998), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1018), .A2(KEYINPUT121), .A3(new_n997), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1050), .A2(new_n1051), .A3(new_n1054), .ZN(new_n1055));
  AND3_X1   g630(.A1(new_n1027), .A2(new_n1045), .A3(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(G303), .A2(G8), .ZN(new_n1057));
  XOR2_X1   g632(.A(new_n1057), .B(KEYINPUT55), .Z(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  XNOR2_X1  g634(.A(KEYINPUT109), .B(G1971), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1032), .A2(new_n1035), .A3(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT114), .ZN(new_n1062));
  AOI21_X1  g637(.A(G2090), .B1(new_n1017), .B2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1063), .B1(new_n1062), .B2(new_n1017), .ZN(new_n1064));
  AND2_X1   g639(.A1(new_n1061), .A2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1059), .B1(new_n1065), .B2(new_n996), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1061), .B1(G2090), .B2(new_n1017), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1067), .A2(G8), .A3(new_n1058), .ZN(new_n1068));
  NAND2_X1  g643(.A1(G305), .A2(G1981), .ZN(new_n1069));
  INV_X1    g644(.A(G1981), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n564), .A2(new_n565), .A3(new_n566), .A4(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT49), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1000), .A2(new_n983), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1069), .A2(KEYINPUT49), .A3(new_n1071), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1074), .A2(new_n1019), .A3(new_n1075), .A4(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n552), .A2(G1976), .A3(new_n555), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT111), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n552), .A2(new_n555), .A3(KEYINPUT111), .A4(G1976), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1075), .A2(new_n1080), .A3(new_n1019), .A4(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT52), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n556), .A2(new_n558), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1083), .B1(new_n1084), .B2(G1976), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1077), .B1(new_n1082), .B2(new_n1085), .ZN(new_n1086));
  AND2_X1   g661(.A1(new_n1082), .A2(KEYINPUT52), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  AND3_X1   g663(.A1(new_n1066), .A2(new_n1068), .A3(new_n1088), .ZN(new_n1089));
  OAI21_X1  g664(.A(KEYINPUT112), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1090));
  OR2_X1    g665(.A1(new_n1082), .A2(new_n1085), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT112), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1082), .A2(KEYINPUT52), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1091), .A2(new_n1092), .A3(new_n1093), .A4(new_n1077), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1090), .A2(new_n1094), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1095), .A2(new_n1067), .A3(G8), .A4(new_n1058), .ZN(new_n1096));
  NOR2_X1   g671(.A1(G288), .A2(G1976), .ZN(new_n1097));
  AND2_X1   g672(.A1(new_n1077), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1071), .ZN(new_n1099));
  OAI211_X1 g674(.A(new_n1019), .B(new_n1075), .C1(new_n1098), .C2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1096), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(KEYINPUT113), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT113), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1096), .A2(new_n1100), .A3(new_n1103), .ZN(new_n1104));
  AOI22_X1  g679(.A1(new_n1056), .A2(new_n1089), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  XNOR2_X1  g680(.A(G299), .B(KEYINPUT57), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1106), .ZN(new_n1107));
  XNOR2_X1  g682(.A(KEYINPUT56), .B(G2072), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1033), .A2(new_n1034), .A3(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(G1956), .ZN(new_n1110));
  AND3_X1   g685(.A1(new_n1017), .A2(KEYINPUT117), .A3(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(KEYINPUT117), .B1(new_n1017), .B2(new_n1110), .ZN(new_n1112));
  OAI211_X1 g687(.A(new_n1107), .B(new_n1109), .C1(new_n1111), .C2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(G1348), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT118), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1075), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1000), .A2(KEYINPUT118), .A3(new_n983), .ZN(new_n1118));
  AOI21_X1  g693(.A(G2067), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n587), .B1(new_n1115), .B2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1109), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(new_n1106), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1114), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT60), .ZN(new_n1124));
  NOR4_X1   g699(.A1(new_n1115), .A2(new_n586), .A3(new_n1124), .A4(new_n1119), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1115), .A2(new_n1119), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n587), .B1(new_n1126), .B2(KEYINPUT60), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(KEYINPUT60), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1125), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT61), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1110), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT117), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1017), .A2(KEYINPUT117), .A3(new_n1110), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1107), .B1(new_n1135), .B2(new_n1109), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1130), .B1(new_n1114), .B2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1122), .A2(KEYINPUT61), .A3(new_n1113), .ZN(new_n1138));
  NOR3_X1   g713(.A1(new_n1030), .A2(new_n1031), .A3(G1996), .ZN(new_n1139));
  XOR2_X1   g714(.A(KEYINPUT58), .B(G1341), .Z(new_n1140));
  AND3_X1   g715(.A1(new_n1117), .A2(new_n1118), .A3(new_n1140), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n527), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(KEYINPUT59), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT59), .ZN(new_n1144));
  OAI211_X1 g719(.A(new_n1144), .B(new_n527), .C1(new_n1139), .C2(new_n1141), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1137), .A2(new_n1138), .A3(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT120), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1129), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1137), .A2(KEYINPUT120), .A3(new_n1146), .A4(new_n1138), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1123), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT54), .ZN(new_n1152));
  AND3_X1   g727(.A1(new_n1041), .A2(KEYINPUT122), .A3(new_n786), .ZN(new_n1153));
  AOI21_X1  g728(.A(KEYINPUT122), .B1(new_n1041), .B2(new_n786), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1156), .A2(G40), .A3(G160), .A4(new_n1043), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1157), .B1(new_n1036), .B2(KEYINPUT53), .ZN(new_n1158));
  NOR3_X1   g733(.A1(new_n1155), .A2(new_n1158), .A3(G171), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1152), .B1(new_n1159), .B2(new_n1045), .ZN(new_n1160));
  OAI21_X1  g735(.A(G171), .B1(new_n1155), .B2(new_n1158), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT123), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1037), .A2(new_n1162), .A3(G301), .A4(new_n1044), .ZN(new_n1163));
  OAI211_X1 g738(.A(new_n1044), .B(G301), .C1(new_n1036), .C2(KEYINPUT53), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(KEYINPUT123), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1161), .A2(new_n1163), .A3(KEYINPUT54), .A4(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1050), .A2(new_n1054), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1160), .A2(new_n1166), .A3(new_n1089), .A4(new_n1167), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1105), .B1(new_n1151), .B2(new_n1168), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1020), .A2(G286), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1066), .A2(new_n1068), .A3(new_n1088), .A4(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT115), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT63), .ZN(new_n1173));
  AND3_X1   g748(.A1(new_n1171), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  NAND4_X1  g749(.A1(new_n1018), .A2(KEYINPUT63), .A3(G168), .A4(new_n1019), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1175), .B1(new_n1090), .B2(new_n1094), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1068), .A2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1058), .B1(new_n1067), .B2(G8), .ZN(new_n1178));
  OAI21_X1  g753(.A(KEYINPUT116), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1067), .A2(G8), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1180), .A2(new_n1059), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT116), .ZN(new_n1182));
  NAND4_X1  g757(.A1(new_n1181), .A2(new_n1182), .A3(new_n1068), .A4(new_n1176), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1179), .A2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1172), .B1(new_n1171), .B2(new_n1173), .ZN(new_n1185));
  NOR3_X1   g760(.A1(new_n1174), .A2(new_n1184), .A3(new_n1185), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n995), .B1(new_n1169), .B2(new_n1186), .ZN(new_n1187));
  OR2_X1    g762(.A1(new_n813), .A2(new_n986), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT46), .ZN(new_n1189));
  INV_X1    g764(.A(G1996), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n985), .A2(new_n1190), .ZN(new_n1191));
  AOI22_X1  g766(.A1(new_n1188), .A2(new_n985), .B1(new_n1189), .B2(new_n1191), .ZN(new_n1192));
  NOR2_X1   g767(.A1(new_n1191), .A2(new_n1189), .ZN(new_n1193));
  INV_X1    g768(.A(new_n1193), .ZN(new_n1194));
  AND2_X1   g769(.A1(new_n1194), .A2(KEYINPUT124), .ZN(new_n1195));
  NOR2_X1   g770(.A1(new_n1194), .A2(KEYINPUT124), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n1192), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  XOR2_X1   g772(.A(new_n1197), .B(KEYINPUT47), .Z(new_n1198));
  INV_X1    g773(.A(KEYINPUT125), .ZN(new_n1199));
  NOR2_X1   g774(.A1(new_n993), .A2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g775(.A(KEYINPUT125), .B1(new_n990), .B2(new_n992), .ZN(new_n1201));
  NAND3_X1  g776(.A1(new_n985), .A2(new_n679), .A3(new_n573), .ZN(new_n1202));
  XOR2_X1   g777(.A(new_n1202), .B(KEYINPUT48), .Z(new_n1203));
  NOR3_X1   g778(.A1(new_n1200), .A2(new_n1201), .A3(new_n1203), .ZN(new_n1204));
  NAND3_X1  g779(.A1(new_n990), .A2(new_n705), .A3(new_n708), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1205), .B1(G2067), .B2(new_n772), .ZN(new_n1206));
  AOI211_X1 g781(.A(new_n1198), .B(new_n1204), .C1(new_n985), .C2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1187), .A2(new_n1207), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g783(.A(KEYINPUT126), .ZN(new_n1210));
  INV_X1    g784(.A(new_n458), .ZN(new_n1211));
  NAND3_X1  g785(.A1(new_n660), .A2(new_n1211), .A3(new_n661), .ZN(new_n1212));
  OAI21_X1  g786(.A(new_n1210), .B1(new_n643), .B2(new_n1212), .ZN(new_n1213));
  INV_X1    g787(.A(new_n1212), .ZN(new_n1214));
  AND2_X1   g788(.A1(new_n641), .A2(new_n642), .ZN(new_n1215));
  OAI211_X1 g789(.A(KEYINPUT126), .B(new_n1214), .C1(new_n1215), .C2(new_n636), .ZN(new_n1216));
  NAND3_X1  g790(.A1(new_n693), .A2(new_n1213), .A3(new_n1216), .ZN(new_n1217));
  AOI21_X1  g791(.A(new_n1217), .B1(new_n896), .B2(new_n899), .ZN(new_n1218));
  INV_X1    g792(.A(KEYINPUT127), .ZN(new_n1219));
  AND3_X1   g793(.A1(new_n1218), .A2(new_n977), .A3(new_n1219), .ZN(new_n1220));
  AOI21_X1  g794(.A(new_n1219), .B1(new_n1218), .B2(new_n977), .ZN(new_n1221));
  NOR2_X1   g795(.A1(new_n1220), .A2(new_n1221), .ZN(G308));
  NAND2_X1  g796(.A1(new_n1218), .A2(new_n977), .ZN(G225));
endmodule


