//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 1 0 1 1 0 1 1 1 0 0 1 0 0 1 0 1 1 1 1 0 1 0 0 1 0 0 1 1 1 0 0 1 0 0 1 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n739, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n835,
    new_n836, new_n838, new_n839, new_n840, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n887, new_n888, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n937,
    new_n938, new_n940, new_n941, new_n942, new_n943, new_n944, new_n946,
    new_n947, new_n948;
  INV_X1    g000(.A(KEYINPUT39), .ZN(new_n202));
  INV_X1    g001(.A(G141gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(G148gat), .ZN(new_n204));
  INV_X1    g003(.A(G148gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G141gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207));
  AOI22_X1  g006(.A1(new_n204), .A2(new_n206), .B1(KEYINPUT2), .B2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(new_n207), .ZN(new_n209));
  NOR2_X1   g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT78), .ZN(new_n211));
  NOR3_X1   g010(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G155gat), .ZN(new_n213));
  INV_X1    g012(.A(G162gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  AOI21_X1  g014(.A(KEYINPUT78), .B1(new_n215), .B2(new_n207), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n208), .B1(new_n212), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT77), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n210), .B1(new_n218), .B2(new_n207), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n209), .A2(KEYINPUT77), .ZN(new_n220));
  AND2_X1   g019(.A1(new_n207), .A2(KEYINPUT2), .ZN(new_n221));
  XNOR2_X1  g020(.A(G141gat), .B(G148gat), .ZN(new_n222));
  OAI211_X1 g021(.A(new_n219), .B(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  AND2_X1   g022(.A1(new_n217), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(G120gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(G113gat), .ZN(new_n226));
  INV_X1    g025(.A(G113gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(G120gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT1), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT67), .ZN(new_n232));
  INV_X1    g031(.A(G134gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(KEYINPUT67), .A2(G134gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n234), .A2(G127gat), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT68), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n233), .A2(G127gat), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  AND3_X1   g038(.A1(new_n236), .A2(new_n237), .A3(new_n239), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n237), .B1(new_n236), .B2(new_n239), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n231), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT4), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT69), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n244), .B1(new_n227), .B2(G120gat), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n225), .A2(KEYINPUT69), .A3(G113gat), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n245), .A2(new_n246), .A3(new_n228), .ZN(new_n247));
  INV_X1    g046(.A(G127gat), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n230), .B1(new_n248), .B2(G134gat), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n249), .A2(new_n238), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n247), .A2(new_n250), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n224), .A2(new_n242), .A3(new_n243), .A4(new_n251), .ZN(new_n252));
  AND2_X1   g051(.A1(KEYINPUT67), .A2(G134gat), .ZN(new_n253));
  NOR2_X1   g052(.A1(KEYINPUT67), .A2(G134gat), .ZN(new_n254));
  NOR3_X1   g053(.A1(new_n253), .A2(new_n254), .A3(new_n248), .ZN(new_n255));
  OAI21_X1  g054(.A(KEYINPUT68), .B1(new_n255), .B2(new_n238), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n236), .A2(new_n237), .A3(new_n239), .ZN(new_n257));
  AOI22_X1  g056(.A1(new_n256), .A2(new_n257), .B1(new_n230), .B2(new_n229), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n217), .A2(new_n251), .A3(new_n223), .ZN(new_n259));
  OAI21_X1  g058(.A(KEYINPUT4), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT81), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n252), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n242), .A2(new_n251), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n217), .A2(new_n223), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(KEYINPUT3), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT3), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n217), .A2(new_n266), .A3(new_n223), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n263), .A2(new_n265), .A3(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n224), .A2(new_n251), .A3(new_n242), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n269), .A2(KEYINPUT81), .A3(KEYINPUT4), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n262), .A2(new_n268), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(G225gat), .A2(G233gat), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  AND3_X1   g072(.A1(new_n271), .A2(KEYINPUT87), .A3(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(KEYINPUT87), .B1(new_n271), .B2(new_n273), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n202), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n271), .A2(new_n273), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT87), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n271), .A2(KEYINPUT87), .A3(new_n273), .ZN(new_n280));
  INV_X1    g079(.A(new_n251), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n258), .A2(new_n281), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n269), .B1(new_n282), .B2(new_n224), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n283), .A2(new_n273), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n284), .A2(new_n202), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n279), .A2(new_n280), .A3(new_n285), .ZN(new_n286));
  XOR2_X1   g085(.A(G1gat), .B(G29gat), .Z(new_n287));
  XNOR2_X1  g086(.A(G57gat), .B(G85gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n287), .B(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n289), .B(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n276), .A2(new_n286), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(KEYINPUT88), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(KEYINPUT40), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT82), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n262), .A2(new_n270), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT5), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n268), .A2(new_n297), .A3(new_n272), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n295), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  AND3_X1   g098(.A1(new_n268), .A2(new_n297), .A3(new_n272), .ZN(new_n300));
  NAND4_X1  g099(.A1(new_n300), .A2(KEYINPUT82), .A3(new_n270), .A4(new_n262), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  AND2_X1   g101(.A1(new_n252), .A2(new_n260), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n265), .A2(new_n267), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n272), .B1(new_n304), .B2(new_n282), .ZN(new_n305));
  OAI21_X1  g104(.A(KEYINPUT79), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n252), .A2(new_n260), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT79), .ZN(new_n308));
  NAND4_X1  g107(.A1(new_n307), .A2(new_n308), .A3(new_n272), .A4(new_n268), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n297), .B1(new_n283), .B2(new_n273), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n306), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n291), .B1(new_n302), .B2(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(G197gat), .B(G204gat), .ZN(new_n313));
  AND2_X1   g112(.A1(G211gat), .A2(G218gat), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n313), .B1(KEYINPUT22), .B2(new_n314), .ZN(new_n315));
  XOR2_X1   g114(.A(G211gat), .B(G218gat), .Z(new_n316));
  XNOR2_X1  g115(.A(new_n315), .B(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(G183gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(KEYINPUT27), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT27), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(G183gat), .ZN(new_n322));
  INV_X1    g121(.A(G190gat), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n320), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  AND2_X1   g123(.A1(KEYINPUT65), .A2(KEYINPUT28), .ZN(new_n325));
  NOR2_X1   g124(.A1(KEYINPUT65), .A2(KEYINPUT28), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n324), .A2(new_n327), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n320), .A2(new_n322), .A3(new_n323), .A4(new_n326), .ZN(new_n329));
  AOI21_X1  g128(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n330), .B1(G169gat), .B2(G176gat), .ZN(new_n331));
  NOR2_X1   g130(.A1(G169gat), .A2(G176gat), .ZN(new_n332));
  AOI22_X1  g131(.A1(new_n332), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n333));
  NAND4_X1  g132(.A1(new_n328), .A2(new_n329), .A3(new_n331), .A4(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT66), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AND2_X1   g135(.A1(new_n331), .A2(new_n333), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n337), .A2(KEYINPUT66), .A3(new_n329), .A4(new_n328), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(G169gat), .A2(G176gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(G183gat), .A2(G190gat), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n340), .B1(new_n341), .B2(KEYINPUT24), .ZN(new_n342));
  OAI21_X1  g141(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT23), .ZN(new_n344));
  INV_X1    g143(.A(G169gat), .ZN(new_n345));
  INV_X1    g144(.A(G176gat), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n344), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n342), .B1(new_n343), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n319), .A2(new_n323), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n349), .A2(KEYINPUT24), .A3(new_n341), .ZN(new_n350));
  AOI21_X1  g149(.A(KEYINPUT25), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  AND2_X1   g150(.A1(G183gat), .A2(G190gat), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT24), .ZN(new_n353));
  AOI22_X1  g152(.A1(new_n352), .A2(new_n353), .B1(G169gat), .B2(G176gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n347), .A2(new_n343), .ZN(new_n355));
  AND4_X1   g154(.A1(KEYINPUT25), .A2(new_n354), .A3(new_n355), .A4(new_n350), .ZN(new_n356));
  OAI21_X1  g155(.A(KEYINPUT64), .B1(new_n351), .B2(new_n356), .ZN(new_n357));
  AND2_X1   g156(.A1(G226gat), .A2(G233gat), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n348), .A2(KEYINPUT25), .A3(new_n350), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n354), .A2(new_n355), .A3(new_n350), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT25), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT64), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n359), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n339), .A2(new_n357), .A3(new_n358), .A4(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n359), .A2(new_n362), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(new_n334), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n358), .A2(KEYINPUT29), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n318), .B1(new_n365), .B2(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n339), .A2(new_n357), .A3(new_n364), .ZN(new_n371));
  INV_X1    g170(.A(new_n367), .ZN(new_n372));
  AOI22_X1  g171(.A1(new_n371), .A2(new_n368), .B1(new_n372), .B2(new_n358), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n370), .B1(new_n373), .B2(new_n318), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT74), .ZN(new_n375));
  XNOR2_X1  g174(.A(G8gat), .B(G36gat), .ZN(new_n376));
  XNOR2_X1  g175(.A(G64gat), .B(G92gat), .ZN(new_n377));
  XOR2_X1   g176(.A(new_n376), .B(new_n377), .Z(new_n378));
  NAND4_X1  g177(.A1(new_n374), .A2(new_n375), .A3(KEYINPUT30), .A4(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n371), .A2(new_n368), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n372), .A2(new_n358), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n380), .A2(new_n318), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n365), .A2(new_n369), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(new_n317), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n382), .A2(new_n384), .A3(KEYINPUT30), .A4(new_n378), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(KEYINPUT74), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n382), .A2(new_n384), .ZN(new_n387));
  INV_X1    g186(.A(new_n378), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  AND3_X1   g188(.A1(new_n379), .A2(new_n386), .A3(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT75), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n391), .B1(new_n387), .B2(new_n388), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n374), .A2(KEYINPUT75), .A3(new_n378), .ZN(new_n393));
  XOR2_X1   g192(.A(KEYINPUT76), .B(KEYINPUT30), .Z(new_n394));
  NAND3_X1  g193(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n312), .B1(new_n390), .B2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT40), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n292), .A2(KEYINPUT88), .A3(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n294), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  XOR2_X1   g198(.A(G78gat), .B(G106gat), .Z(new_n400));
  XNOR2_X1  g199(.A(new_n400), .B(KEYINPUT85), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n401), .B(G22gat), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT29), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT86), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n315), .A2(new_n405), .A3(new_n316), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n404), .B(new_n406), .C1(new_n317), .C2(new_n405), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n224), .B1(new_n407), .B2(new_n266), .ZN(new_n408));
  AND2_X1   g207(.A1(G228gat), .A2(G233gat), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n317), .B1(new_n404), .B2(new_n267), .ZN(new_n410));
  OR3_X1    g209(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n317), .A2(new_n404), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n224), .B1(new_n412), .B2(new_n266), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n409), .B1(new_n413), .B2(new_n410), .ZN(new_n414));
  XNOR2_X1  g213(.A(KEYINPUT31), .B(G50gat), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n411), .A2(new_n414), .A3(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n416), .B1(new_n411), .B2(new_n414), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n403), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n419), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n421), .A2(new_n402), .A3(new_n417), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n399), .A2(new_n423), .ZN(new_n424));
  AND2_X1   g223(.A1(new_n262), .A2(new_n270), .ZN(new_n425));
  AOI21_X1  g224(.A(KEYINPUT82), .B1(new_n425), .B2(new_n300), .ZN(new_n426));
  NOR3_X1   g225(.A1(new_n296), .A2(new_n295), .A3(new_n298), .ZN(new_n427));
  OAI211_X1 g226(.A(new_n291), .B(new_n311), .C1(new_n426), .C2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT83), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n302), .A2(new_n311), .ZN(new_n431));
  INV_X1    g230(.A(new_n291), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT6), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n302), .A2(KEYINPUT83), .A3(new_n291), .A4(new_n311), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n430), .A2(new_n433), .A3(new_n434), .A4(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n392), .A2(new_n393), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT37), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n378), .B1(new_n374), .B2(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n438), .B1(new_n373), .B2(new_n317), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n383), .A2(new_n318), .ZN(new_n441));
  AOI21_X1  g240(.A(KEYINPUT38), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n437), .B1(new_n439), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n312), .A2(KEYINPUT6), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n436), .A2(new_n443), .A3(KEYINPUT89), .A4(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT38), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n387), .A2(KEYINPUT37), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n446), .B1(new_n439), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n436), .A2(new_n444), .A3(new_n443), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT89), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n448), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n424), .B1(new_n445), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n371), .A2(new_n282), .ZN(new_n453));
  NAND2_X1  g252(.A1(G227gat), .A2(G233gat), .ZN(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n339), .A2(new_n263), .A3(new_n357), .A4(new_n364), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n453), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT33), .ZN(new_n458));
  XNOR2_X1  g257(.A(G15gat), .B(G43gat), .ZN(new_n459));
  XNOR2_X1  g258(.A(new_n459), .B(KEYINPUT70), .ZN(new_n460));
  XNOR2_X1  g259(.A(G71gat), .B(G99gat), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n460), .B(new_n461), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n457), .B(KEYINPUT32), .C1(new_n458), .C2(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n462), .B1(new_n457), .B2(KEYINPUT32), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n457), .A2(new_n458), .ZN(new_n465));
  AND3_X1   g264(.A1(new_n464), .A2(KEYINPUT71), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(KEYINPUT71), .B1(new_n464), .B2(new_n465), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n455), .B1(new_n453), .B2(new_n456), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT34), .ZN(new_n470));
  OAI21_X1  g269(.A(KEYINPUT72), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR3_X1   g270(.A1(new_n351), .A2(new_n356), .A3(KEYINPUT64), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n363), .B1(new_n359), .B2(new_n362), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n263), .B1(new_n474), .B2(new_n339), .ZN(new_n475));
  INV_X1    g274(.A(new_n456), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n454), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT72), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n477), .A2(new_n478), .A3(KEYINPUT34), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n470), .B(new_n454), .C1(new_n475), .C2(new_n476), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(KEYINPUT73), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT73), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n469), .A2(new_n482), .A3(new_n470), .ZN(new_n483));
  AOI22_X1  g282(.A1(new_n471), .A2(new_n479), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n468), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT36), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n484), .B(new_n463), .C1(new_n467), .C2(new_n466), .ZN(new_n488));
  AND3_X1   g287(.A1(new_n486), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n487), .B1(new_n486), .B2(new_n488), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n390), .A2(new_n395), .ZN(new_n492));
  INV_X1    g291(.A(new_n444), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n493), .B1(new_n436), .B2(KEYINPUT84), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n312), .A2(KEYINPUT6), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT84), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n495), .A2(new_n496), .A3(new_n435), .A4(new_n430), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n492), .B1(new_n494), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n491), .B1(new_n498), .B2(new_n423), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT35), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n486), .A2(new_n423), .A3(new_n488), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n500), .B1(new_n498), .B2(new_n501), .ZN(new_n502));
  AND2_X1   g301(.A1(new_n486), .A2(new_n488), .ZN(new_n503));
  INV_X1    g302(.A(new_n492), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n436), .A2(new_n444), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n506), .A2(new_n500), .A3(new_n423), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  OAI22_X1  g307(.A1(new_n452), .A2(new_n499), .B1(new_n502), .B2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(G36gat), .ZN(new_n510));
  AND2_X1   g309(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n511));
  NOR2_X1   g310(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(G29gat), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n514), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT15), .ZN(new_n517));
  XNOR2_X1  g316(.A(G43gat), .B(G50gat), .ZN(new_n518));
  OR2_X1    g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n516), .A2(KEYINPUT15), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n517), .A2(new_n518), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n522), .B(KEYINPUT17), .ZN(new_n523));
  XNOR2_X1  g322(.A(G15gat), .B(G22gat), .ZN(new_n524));
  INV_X1    g323(.A(G1gat), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n524), .A2(KEYINPUT16), .A3(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT91), .ZN(new_n527));
  OAI221_X1 g326(.A(new_n526), .B1(new_n527), .B2(G8gat), .C1(new_n525), .C2(new_n524), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(G8gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n528), .B(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n523), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(G229gat), .A2(G233gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n530), .A2(new_n522), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT18), .ZN(new_n536));
  OR2_X1    g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  XOR2_X1   g336(.A(new_n533), .B(KEYINPUT13), .Z(new_n538));
  INV_X1    g337(.A(new_n534), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n530), .A2(new_n522), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n535), .A2(new_n536), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n537), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(G113gat), .B(G141gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(KEYINPUT90), .B(KEYINPUT11), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  XOR2_X1   g345(.A(G169gat), .B(G197gat), .Z(new_n547));
  XNOR2_X1  g346(.A(new_n546), .B(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(KEYINPUT12), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n543), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n537), .A2(new_n541), .A3(new_n542), .A4(new_n549), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT97), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(KEYINPUT7), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT7), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(KEYINPUT97), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n555), .A2(new_n557), .A3(G85gat), .A4(G92gat), .ZN(new_n558));
  INV_X1    g357(.A(G85gat), .ZN(new_n559));
  INV_X1    g358(.A(G92gat), .ZN(new_n560));
  OAI211_X1 g359(.A(KEYINPUT97), .B(new_n556), .C1(new_n559), .C2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(G99gat), .A2(G106gat), .ZN(new_n562));
  AOI22_X1  g361(.A1(KEYINPUT8), .A2(new_n562), .B1(new_n559), .B2(new_n560), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n558), .A2(new_n561), .A3(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(G99gat), .B(G106gat), .ZN(new_n565));
  XOR2_X1   g364(.A(new_n564), .B(new_n565), .Z(new_n566));
  NAND2_X1  g365(.A1(new_n523), .A2(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n564), .B(new_n565), .ZN(new_n568));
  NAND2_X1  g367(.A1(G232gat), .A2(G233gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n569), .B(KEYINPUT96), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  AOI22_X1  g370(.A1(new_n522), .A2(new_n568), .B1(KEYINPUT41), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n567), .A2(new_n572), .ZN(new_n573));
  XOR2_X1   g372(.A(G190gat), .B(G218gat), .Z(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n573), .B(new_n575), .ZN(new_n576));
  OR2_X1    g375(.A1(new_n571), .A2(KEYINPUT41), .ZN(new_n577));
  XOR2_X1   g376(.A(G134gat), .B(G162gat), .Z(new_n578));
  XNOR2_X1  g377(.A(new_n577), .B(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n576), .B(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(G57gat), .B(G64gat), .ZN(new_n581));
  AOI21_X1  g380(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n582));
  OR2_X1    g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(G71gat), .B(G78gat), .ZN(new_n584));
  XOR2_X1   g383(.A(new_n583), .B(new_n584), .Z(new_n585));
  XNOR2_X1  g384(.A(KEYINPUT92), .B(KEYINPUT21), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  XOR2_X1   g386(.A(KEYINPUT94), .B(KEYINPUT19), .Z(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n583), .B(new_n584), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n530), .B1(KEYINPUT21), .B2(new_n590), .ZN(new_n591));
  XOR2_X1   g390(.A(new_n589), .B(new_n591), .Z(new_n592));
  XNOR2_X1  g391(.A(G127gat), .B(G155gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(KEYINPUT20), .ZN(new_n594));
  NAND2_X1  g393(.A1(G231gat), .A2(G233gat), .ZN(new_n595));
  XOR2_X1   g394(.A(new_n595), .B(KEYINPUT93), .Z(new_n596));
  XNOR2_X1  g395(.A(new_n594), .B(new_n596), .ZN(new_n597));
  XOR2_X1   g396(.A(G183gat), .B(G211gat), .Z(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(KEYINPUT95), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n597), .B(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n592), .B(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n580), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n568), .A2(new_n590), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT10), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(KEYINPUT100), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n566), .A2(new_n585), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n607), .A2(KEYINPUT98), .A3(new_n603), .ZN(new_n608));
  OR3_X1    g407(.A1(new_n568), .A2(new_n590), .A3(KEYINPUT98), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g409(.A(KEYINPUT99), .B1(new_n610), .B2(new_n604), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT99), .ZN(new_n612));
  AOI211_X1 g411(.A(new_n612), .B(KEYINPUT10), .C1(new_n608), .C2(new_n609), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n606), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(G230gat), .A2(G233gat), .ZN(new_n615));
  XOR2_X1   g414(.A(new_n615), .B(KEYINPUT101), .Z(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  OR2_X1    g417(.A1(new_n610), .A2(new_n615), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(G120gat), .B(G148gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(G176gat), .B(G204gat), .ZN(new_n622));
  XOR2_X1   g421(.A(new_n621), .B(new_n622), .Z(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n614), .A2(new_n615), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n626), .A2(new_n619), .A3(new_n623), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n602), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n509), .A2(new_n553), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(KEYINPUT102), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT102), .ZN(new_n632));
  NAND4_X1  g431(.A1(new_n509), .A2(new_n632), .A3(new_n553), .A4(new_n629), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n436), .A2(KEYINPUT84), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n635), .A2(new_n444), .A3(new_n497), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT103), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n494), .A2(KEYINPUT103), .A3(new_n497), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n634), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(G1gat), .ZN(G1324gat));
  INV_X1    g442(.A(KEYINPUT106), .ZN(new_n644));
  XOR2_X1   g443(.A(KEYINPUT104), .B(KEYINPUT42), .Z(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n553), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n449), .A2(new_n450), .ZN(new_n648));
  INV_X1    g447(.A(new_n448), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n648), .A2(new_n445), .A3(new_n649), .ZN(new_n650));
  AND2_X1   g449(.A1(new_n399), .A2(new_n423), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n504), .ZN(new_n653));
  INV_X1    g452(.A(new_n423), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n652), .A2(new_n655), .A3(new_n491), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n636), .A2(new_n504), .A3(new_n501), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n657), .A2(KEYINPUT35), .ZN(new_n658));
  OR2_X1    g457(.A1(new_n505), .A2(new_n507), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n647), .B1(new_n656), .B2(new_n660), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n632), .B1(new_n661), .B2(new_n629), .ZN(new_n662));
  AND4_X1   g461(.A1(new_n632), .A2(new_n509), .A3(new_n553), .A4(new_n629), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n492), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(KEYINPUT105), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT105), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n634), .A2(new_n666), .A3(new_n492), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g467(.A(KEYINPUT16), .B(G8gat), .Z(new_n669));
  AOI21_X1  g468(.A(new_n646), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n665), .A2(G8gat), .A3(new_n667), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n669), .A2(KEYINPUT42), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n664), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n644), .B1(new_n670), .B2(new_n675), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n666), .B1(new_n634), .B2(new_n492), .ZN(new_n677));
  AOI211_X1 g476(.A(KEYINPUT105), .B(new_n504), .C1(new_n631), .C2(new_n633), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n673), .B1(new_n679), .B2(G8gat), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n669), .B1(new_n677), .B2(new_n678), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(new_n645), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n680), .A2(new_n682), .A3(KEYINPUT106), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n676), .A2(new_n683), .ZN(G1325gat));
  INV_X1    g483(.A(new_n634), .ZN(new_n685));
  INV_X1    g484(.A(new_n503), .ZN(new_n686));
  OR3_X1    g485(.A1(new_n685), .A2(G15gat), .A3(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(G15gat), .B1(new_n685), .B2(new_n491), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(G1326gat));
  NAND2_X1  g488(.A1(new_n634), .A2(new_n654), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(KEYINPUT107), .ZN(new_n691));
  XOR2_X1   g490(.A(KEYINPUT43), .B(G22gat), .Z(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(G1327gat));
  INV_X1    g492(.A(new_n601), .ZN(new_n694));
  INV_X1    g493(.A(new_n579), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n576), .B(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n628), .ZN(new_n697));
  AND4_X1   g496(.A1(new_n661), .A2(new_n694), .A3(new_n696), .A4(new_n697), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n698), .A2(new_n514), .A3(new_n641), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(KEYINPUT45), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n580), .B1(new_n656), .B2(new_n660), .ZN(new_n701));
  OR2_X1    g500(.A1(new_n701), .A2(KEYINPUT44), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(KEYINPUT44), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n647), .A2(new_n628), .A3(new_n601), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(G29gat), .B1(new_n706), .B2(new_n640), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n700), .A2(new_n707), .ZN(G1328gat));
  NAND3_X1  g507(.A1(new_n698), .A2(new_n510), .A3(new_n492), .ZN(new_n709));
  XOR2_X1   g508(.A(new_n709), .B(KEYINPUT46), .Z(new_n710));
  OAI21_X1  g509(.A(G36gat), .B1(new_n706), .B2(new_n504), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(G1329gat));
  OAI21_X1  g511(.A(G43gat), .B1(new_n706), .B2(new_n491), .ZN(new_n713));
  INV_X1    g512(.A(G43gat), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n698), .A2(new_n714), .A3(new_n503), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT47), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n713), .A2(KEYINPUT47), .A3(new_n715), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(G1330gat));
  NAND2_X1  g519(.A1(new_n654), .A2(G50gat), .ZN(new_n721));
  AND2_X1   g520(.A1(new_n698), .A2(new_n654), .ZN(new_n722));
  OAI22_X1  g521(.A1(new_n706), .A2(new_n721), .B1(G50gat), .B2(new_n722), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT48), .ZN(G1331gat));
  NOR3_X1   g523(.A1(new_n602), .A2(new_n697), .A3(new_n553), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n509), .A2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(new_n641), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g528(.A(new_n504), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n727), .A2(new_n730), .ZN(new_n731));
  XOR2_X1   g530(.A(new_n731), .B(KEYINPUT108), .Z(new_n732));
  NOR2_X1   g531(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n732), .B(new_n733), .ZN(G1333gat));
  OR3_X1    g533(.A1(new_n726), .A2(G71gat), .A3(new_n686), .ZN(new_n735));
  OAI21_X1  g534(.A(G71gat), .B1(new_n726), .B2(new_n491), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  XOR2_X1   g536(.A(new_n737), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g537(.A1(new_n727), .A2(new_n654), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g539(.A1(new_n553), .A2(new_n601), .ZN(new_n741));
  INV_X1    g540(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n742), .A2(new_n697), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n704), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(G85gat), .B1(new_n744), .B2(new_n640), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT51), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n509), .A2(new_n696), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n746), .B1(new_n747), .B2(new_n742), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n701), .A2(KEYINPUT51), .A3(new_n741), .ZN(new_n749));
  AND2_X1   g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n641), .A2(new_n559), .A3(new_n628), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n745), .B1(new_n750), .B2(new_n751), .ZN(G1336gat));
  INV_X1    g551(.A(KEYINPUT110), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT109), .ZN(new_n754));
  OR2_X1    g553(.A1(new_n748), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n748), .A2(new_n754), .A3(new_n749), .ZN(new_n756));
  NOR3_X1   g555(.A1(new_n697), .A2(G92gat), .A3(new_n504), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n755), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n702), .A2(new_n492), .A3(new_n703), .A4(new_n743), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(G92gat), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n753), .B1(new_n761), .B2(KEYINPUT52), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT52), .ZN(new_n763));
  AOI211_X1 g562(.A(KEYINPUT110), .B(new_n763), .C1(new_n758), .C2(new_n760), .ZN(new_n764));
  INV_X1    g563(.A(new_n760), .ZN(new_n765));
  INV_X1    g564(.A(new_n757), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n763), .B1(new_n750), .B2(new_n766), .ZN(new_n767));
  OAI22_X1  g566(.A1(new_n762), .A2(new_n764), .B1(new_n765), .B2(new_n767), .ZN(G1337gat));
  OAI21_X1  g567(.A(G99gat), .B1(new_n744), .B2(new_n491), .ZN(new_n769));
  OR3_X1    g568(.A1(new_n686), .A2(new_n697), .A3(G99gat), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n769), .B1(new_n750), .B2(new_n770), .ZN(G1338gat));
  OAI21_X1  g570(.A(G106gat), .B1(new_n744), .B2(new_n423), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n697), .A2(G106gat), .A3(new_n423), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n755), .A2(new_n756), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(KEYINPUT53), .ZN(new_n776));
  INV_X1    g575(.A(new_n750), .ZN(new_n777));
  AOI21_X1  g576(.A(KEYINPUT53), .B1(new_n777), .B2(new_n773), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n772), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n776), .A2(new_n779), .ZN(G1339gat));
  INV_X1    g579(.A(KEYINPUT55), .ZN(new_n781));
  OAI211_X1 g580(.A(new_n616), .B(new_n606), .C1(new_n611), .C2(new_n613), .ZN(new_n782));
  AND3_X1   g581(.A1(new_n626), .A2(KEYINPUT54), .A3(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT54), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n614), .A2(new_n784), .A3(new_n617), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(new_n624), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n781), .B1(new_n783), .B2(new_n786), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n626), .A2(KEYINPUT54), .A3(new_n782), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n788), .A2(KEYINPUT55), .A3(new_n624), .A4(new_n785), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n787), .A2(new_n789), .A3(new_n553), .A4(new_n627), .ZN(new_n790));
  INV_X1    g589(.A(new_n552), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n539), .A2(new_n540), .ZN(new_n792));
  INV_X1    g591(.A(new_n538), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT113), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n794), .B(new_n795), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n533), .B1(new_n532), .B2(new_n534), .ZN(new_n797));
  OR2_X1    g596(.A1(new_n797), .A2(KEYINPUT112), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(KEYINPUT112), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n796), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n791), .B1(new_n548), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(new_n628), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n696), .B1(new_n790), .B2(new_n802), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n787), .A2(new_n789), .A3(new_n696), .A4(new_n627), .ZN(new_n804));
  INV_X1    g603(.A(new_n801), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n694), .B1(new_n803), .B2(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n697), .A2(new_n601), .A3(new_n580), .ZN(new_n808));
  OAI21_X1  g607(.A(KEYINPUT111), .B1(new_n808), .B2(new_n553), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT111), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n629), .A2(new_n810), .A3(new_n647), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n807), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(new_n423), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(KEYINPUT114), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n654), .B1(new_n807), .B2(new_n812), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT114), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n640), .A2(new_n505), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(G113gat), .B1(new_n821), .B2(new_n647), .ZN(new_n822));
  INV_X1    g621(.A(new_n820), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n814), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n824), .A2(new_n227), .A3(new_n553), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n822), .A2(new_n825), .ZN(new_n826));
  XNOR2_X1  g625(.A(new_n826), .B(KEYINPUT115), .ZN(G1340gat));
  NAND3_X1  g626(.A1(new_n824), .A2(new_n225), .A3(new_n628), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n823), .B1(new_n815), .B2(new_n818), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n225), .B1(new_n829), .B2(new_n628), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT116), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n830), .A2(new_n831), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n828), .B1(new_n832), .B2(new_n833), .ZN(G1341gat));
  OAI21_X1  g633(.A(G127gat), .B1(new_n821), .B2(new_n694), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n824), .A2(new_n248), .A3(new_n601), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(G1342gat));
  NAND4_X1  g636(.A1(new_n824), .A2(new_n234), .A3(new_n235), .A4(new_n696), .ZN(new_n838));
  XOR2_X1   g637(.A(new_n838), .B(KEYINPUT56), .Z(new_n839));
  OAI21_X1  g638(.A(G134gat), .B1(new_n821), .B2(new_n580), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(G1343gat));
  NOR3_X1   g640(.A1(new_n640), .A2(new_n490), .A3(new_n489), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(new_n504), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n423), .B1(new_n807), .B2(new_n812), .ZN(new_n844));
  OR2_X1    g643(.A1(new_n844), .A2(KEYINPUT57), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT57), .ZN(new_n846));
  AOI211_X1 g645(.A(new_n846), .B(new_n423), .C1(new_n807), .C2(new_n812), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n843), .B1(new_n845), .B2(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n203), .B1(new_n849), .B2(new_n553), .ZN(new_n850));
  XNOR2_X1  g649(.A(KEYINPUT118), .B(KEYINPUT58), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n553), .A2(new_n203), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n844), .A2(new_n842), .ZN(new_n854));
  OR2_X1    g653(.A1(new_n854), .A2(KEYINPUT117), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(KEYINPUT117), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n855), .A2(new_n504), .A3(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n852), .B1(new_n853), .B2(new_n857), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n854), .A2(new_n492), .A3(new_n853), .ZN(new_n859));
  OAI21_X1  g658(.A(KEYINPUT58), .B1(new_n850), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n858), .A2(new_n860), .ZN(G1344gat));
  NAND2_X1  g660(.A1(new_n849), .A2(new_n628), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT59), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n862), .A2(new_n863), .A3(G148gat), .ZN(new_n864));
  AND2_X1   g663(.A1(new_n789), .A2(new_n627), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT119), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n865), .A2(new_n866), .A3(new_n696), .A4(new_n787), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n804), .A2(KEYINPUT119), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n867), .A2(new_n868), .A3(new_n801), .ZN(new_n869));
  INV_X1    g668(.A(new_n803), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n601), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n808), .A2(new_n553), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n654), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n847), .B1(new_n846), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n842), .A2(new_n504), .A3(new_n628), .ZN(new_n875));
  OAI21_X1  g674(.A(G148gat), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n876), .A2(KEYINPUT120), .A3(KEYINPUT59), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(KEYINPUT120), .B1(new_n876), .B2(KEYINPUT59), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n864), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(new_n857), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n881), .A2(new_n205), .A3(new_n628), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n880), .A2(new_n882), .ZN(G1345gat));
  NAND3_X1  g682(.A1(new_n881), .A2(new_n213), .A3(new_n601), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n849), .A2(new_n601), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n884), .B1(new_n213), .B2(new_n885), .ZN(G1346gat));
  NAND2_X1  g685(.A1(new_n849), .A2(new_n696), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n214), .B1(new_n887), .B2(KEYINPUT121), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n888), .B1(KEYINPUT121), .B2(new_n887), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n881), .A2(new_n214), .A3(new_n696), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(G1347gat));
  AOI21_X1  g690(.A(new_n641), .B1(new_n807), .B2(new_n812), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n892), .A2(new_n492), .A3(new_n501), .ZN(new_n893));
  XNOR2_X1  g692(.A(new_n893), .B(KEYINPUT122), .ZN(new_n894));
  AOI21_X1  g693(.A(G169gat), .B1(new_n894), .B2(new_n553), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n640), .A2(new_n492), .A3(new_n503), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n896), .B1(new_n815), .B2(new_n818), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n647), .A2(new_n345), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n895), .B1(new_n897), .B2(new_n898), .ZN(G1348gat));
  NAND3_X1  g698(.A1(new_n894), .A2(new_n346), .A3(new_n628), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n897), .A2(new_n628), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n900), .B1(new_n901), .B2(new_n346), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(KEYINPUT123), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT123), .ZN(new_n904));
  OAI211_X1 g703(.A(new_n900), .B(new_n904), .C1(new_n901), .C2(new_n346), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n903), .A2(new_n905), .ZN(G1349gat));
  INV_X1    g705(.A(KEYINPUT125), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n601), .A2(new_n320), .A3(new_n322), .ZN(new_n908));
  OR2_X1    g707(.A1(new_n893), .A2(new_n908), .ZN(new_n909));
  AOI211_X1 g708(.A(new_n694), .B(new_n896), .C1(new_n815), .C2(new_n818), .ZN(new_n910));
  OAI211_X1 g709(.A(new_n907), .B(new_n909), .C1(new_n910), .C2(new_n319), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT124), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT60), .ZN(new_n914));
  OAI221_X1 g713(.A(new_n909), .B1(KEYINPUT124), .B2(new_n914), .C1(new_n910), .C2(new_n319), .ZN(new_n915));
  AOI22_X1  g714(.A1(new_n913), .A2(new_n915), .B1(new_n914), .B2(new_n911), .ZN(G1350gat));
  AOI21_X1  g715(.A(new_n323), .B1(new_n897), .B2(new_n696), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT126), .ZN(new_n918));
  OR2_X1    g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n917), .A2(new_n918), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n919), .A2(KEYINPUT61), .A3(new_n920), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n917), .A2(new_n918), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT61), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n580), .A2(G190gat), .ZN(new_n924));
  AOI22_X1  g723(.A1(new_n922), .A2(new_n923), .B1(new_n894), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n921), .A2(new_n925), .ZN(G1351gat));
  AND4_X1   g725(.A1(new_n654), .A2(new_n892), .A3(new_n492), .A4(new_n491), .ZN(new_n927));
  AOI21_X1  g726(.A(G197gat), .B1(new_n927), .B2(new_n553), .ZN(new_n928));
  INV_X1    g727(.A(new_n874), .ZN(new_n929));
  AND3_X1   g728(.A1(new_n640), .A2(new_n492), .A3(new_n491), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(new_n931), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n553), .A2(G197gat), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n928), .B1(new_n932), .B2(new_n933), .ZN(G1352gat));
  INV_X1    g733(.A(G204gat), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n927), .A2(new_n935), .A3(new_n628), .ZN(new_n936));
  XOR2_X1   g735(.A(new_n936), .B(KEYINPUT62), .Z(new_n937));
  OAI21_X1  g736(.A(G204gat), .B1(new_n931), .B2(new_n697), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(G1353gat));
  INV_X1    g738(.A(G211gat), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n927), .A2(new_n940), .A3(new_n601), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n929), .A2(new_n601), .A3(new_n930), .ZN(new_n942));
  AND3_X1   g741(.A1(new_n942), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n943));
  AOI21_X1  g742(.A(KEYINPUT63), .B1(new_n942), .B2(G211gat), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n941), .B1(new_n943), .B2(new_n944), .ZN(G1354gat));
  AOI21_X1  g744(.A(G218gat), .B1(new_n927), .B2(new_n696), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n696), .A2(G218gat), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(KEYINPUT127), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n946), .B1(new_n932), .B2(new_n948), .ZN(G1355gat));
endmodule


