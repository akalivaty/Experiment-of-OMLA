//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 1 0 0 1 0 1 0 1 0 0 0 0 0 1 0 1 1 1 1 1 1 1 1 0 1 0 0 0 1 1 0 0 0 1 1 1 1 0 0 1 1 0 1 1 1 0 0 0 1 0 0 0 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:00 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n703, new_n704, new_n706,
    new_n707, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n749, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990;
  INV_X1    g000(.A(KEYINPUT75), .ZN(new_n187));
  INV_X1    g001(.A(G472), .ZN(new_n188));
  INV_X1    g002(.A(G902), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT70), .B(G953), .ZN(new_n191));
  INV_X1    g005(.A(G237), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n191), .A2(G210), .A3(new_n192), .ZN(new_n193));
  XOR2_X1   g007(.A(KEYINPUT71), .B(KEYINPUT27), .Z(new_n194));
  XNOR2_X1  g008(.A(new_n193), .B(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT26), .B(G101), .ZN(new_n196));
  XNOR2_X1  g010(.A(new_n195), .B(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G119), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G116), .ZN(new_n199));
  INV_X1    g013(.A(G116), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G119), .ZN(new_n201));
  INV_X1    g015(.A(G113), .ZN(new_n202));
  AND2_X1   g016(.A1(new_n202), .A2(KEYINPUT2), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n202), .A2(KEYINPUT2), .ZN(new_n204));
  OAI211_X1 g018(.A(new_n199), .B(new_n201), .C1(new_n203), .C2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n199), .A2(new_n201), .ZN(new_n206));
  XNOR2_X1  g020(.A(KEYINPUT2), .B(G113), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT68), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n205), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n206), .A2(new_n207), .A3(KEYINPUT68), .ZN(new_n211));
  AND2_X1   g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  XNOR2_X1  g027(.A(G143), .B(G146), .ZN(new_n214));
  XNOR2_X1  g028(.A(KEYINPUT0), .B(G128), .ZN(new_n215));
  OAI21_X1  g029(.A(KEYINPUT64), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G146), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G143), .ZN(new_n218));
  INV_X1    g032(.A(G143), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G146), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT64), .ZN(new_n222));
  NAND2_X1  g036(.A1(KEYINPUT0), .A2(G128), .ZN(new_n223));
  OR2_X1    g037(.A1(KEYINPUT0), .A2(G128), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n221), .A2(new_n222), .A3(new_n223), .A4(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n214), .A2(KEYINPUT0), .A3(G128), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n216), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT11), .ZN(new_n229));
  INV_X1    g043(.A(G134), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n229), .B1(new_n230), .B2(G137), .ZN(new_n231));
  INV_X1    g045(.A(G137), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n232), .A2(KEYINPUT11), .A3(G134), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n230), .A2(G137), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n231), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G131), .ZN(new_n236));
  INV_X1    g050(.A(G131), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n231), .A2(new_n233), .A3(new_n237), .A4(new_n234), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n228), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G128), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n241), .A2(KEYINPUT1), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n242), .A2(new_n218), .A3(new_n220), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT66), .ZN(new_n245));
  OAI211_X1 g059(.A(new_n245), .B(KEYINPUT1), .C1(new_n219), .C2(G146), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G128), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n245), .B1(new_n218), .B2(KEYINPUT1), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n221), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(KEYINPUT67), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT67), .ZN(new_n251));
  OAI211_X1 g065(.A(new_n251), .B(new_n221), .C1(new_n247), .C2(new_n248), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n244), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n234), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n230), .A2(G137), .ZN(new_n255));
  OAI21_X1  g069(.A(G131), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(new_n238), .ZN(new_n257));
  OAI211_X1 g071(.A(new_n213), .B(new_n240), .C1(new_n253), .C2(new_n257), .ZN(new_n258));
  OAI211_X1 g072(.A(new_n240), .B(KEYINPUT30), .C1(new_n253), .C2(new_n257), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n259), .A2(KEYINPUT69), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT69), .ZN(new_n261));
  AND2_X1   g075(.A1(new_n236), .A2(new_n238), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n262), .A2(new_n227), .ZN(new_n263));
  INV_X1    g077(.A(new_n252), .ZN(new_n264));
  OAI21_X1  g078(.A(KEYINPUT1), .B1(new_n219), .B2(G146), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(KEYINPUT66), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n266), .A2(G128), .A3(new_n246), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n251), .B1(new_n267), .B2(new_n221), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n243), .B1(new_n264), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n257), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n263), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n261), .B1(new_n271), .B2(KEYINPUT30), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT30), .ZN(new_n273));
  OAI21_X1  g087(.A(KEYINPUT65), .B1(new_n262), .B2(new_n227), .ZN(new_n274));
  AND2_X1   g088(.A1(new_n225), .A2(new_n226), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT65), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n275), .A2(new_n276), .A3(new_n239), .A4(new_n216), .ZN(new_n277));
  AND2_X1   g091(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n253), .A2(new_n257), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n273), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n260), .B1(new_n272), .B2(new_n280), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n197), .B(new_n258), .C1(new_n281), .C2(new_n213), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT31), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(new_n258), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n271), .A2(new_n261), .A3(KEYINPUT30), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n259), .A2(KEYINPUT69), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n269), .A2(new_n270), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n274), .A2(new_n277), .ZN(new_n289));
  AOI21_X1  g103(.A(KEYINPUT30), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n286), .B1(new_n287), .B2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n285), .B1(new_n291), .B2(new_n212), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n292), .A2(KEYINPUT31), .A3(new_n197), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n284), .A2(new_n293), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n285), .A2(KEYINPUT28), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n213), .B1(new_n288), .B2(new_n289), .ZN(new_n296));
  OAI21_X1  g110(.A(KEYINPUT28), .B1(new_n296), .B2(new_n285), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT72), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n295), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  OAI211_X1 g113(.A(KEYINPUT72), .B(KEYINPUT28), .C1(new_n296), .C2(new_n285), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n197), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n190), .B1(new_n294), .B2(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n187), .B1(new_n304), .B2(KEYINPUT32), .ZN(new_n305));
  AOI22_X1  g119(.A1(new_n284), .A2(new_n293), .B1(new_n302), .B2(new_n301), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT32), .ZN(new_n307));
  NOR4_X1   g121(.A1(new_n306), .A2(KEYINPUT75), .A3(new_n307), .A4(new_n190), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n301), .A2(new_n197), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n292), .A2(new_n302), .ZN(new_n311));
  AOI21_X1  g125(.A(KEYINPUT29), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  XNOR2_X1  g126(.A(new_n271), .B(new_n213), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n295), .B1(new_n313), .B2(KEYINPUT28), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n314), .A2(KEYINPUT29), .A3(new_n197), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(new_n189), .ZN(new_n316));
  OAI21_X1  g130(.A(G472), .B1(new_n312), .B2(new_n316), .ZN(new_n317));
  XOR2_X1   g131(.A(KEYINPUT73), .B(KEYINPUT32), .Z(new_n318));
  OAI21_X1  g132(.A(KEYINPUT74), .B1(new_n304), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT74), .ZN(new_n320));
  INV_X1    g134(.A(new_n318), .ZN(new_n321));
  OAI211_X1 g135(.A(new_n320), .B(new_n321), .C1(new_n306), .C2(new_n190), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n309), .A2(new_n317), .A3(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(G217), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n325), .B1(G234), .B2(new_n189), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n191), .A2(G221), .A3(G234), .ZN(new_n328));
  OR2_X1    g142(.A1(new_n328), .A2(KEYINPUT79), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(KEYINPUT79), .ZN(new_n330));
  XNOR2_X1  g144(.A(KEYINPUT22), .B(G137), .ZN(new_n331));
  AND3_X1   g145(.A1(new_n329), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n331), .B1(new_n329), .B2(new_n330), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT16), .ZN(new_n336));
  INV_X1    g150(.A(G140), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n336), .A2(new_n337), .A3(G125), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(G125), .ZN(new_n339));
  INV_X1    g153(.A(G125), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(G140), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  OAI211_X1 g156(.A(G146), .B(new_n338), .C1(new_n342), .C2(new_n336), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT78), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n339), .A2(new_n341), .A3(KEYINPUT78), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n345), .A2(new_n217), .A3(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT76), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n348), .B1(new_n198), .B2(G128), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n198), .A2(G128), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n241), .A2(KEYINPUT76), .A3(G119), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  XNOR2_X1  g166(.A(KEYINPUT24), .B(G110), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n241), .A2(KEYINPUT23), .A3(G119), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n198), .A2(G128), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n355), .B(new_n350), .C1(new_n356), .C2(KEYINPUT23), .ZN(new_n357));
  OAI22_X1  g171(.A1(new_n354), .A2(KEYINPUT77), .B1(G110), .B2(new_n357), .ZN(new_n358));
  AND2_X1   g172(.A1(new_n354), .A2(KEYINPUT77), .ZN(new_n359));
  OAI211_X1 g173(.A(new_n343), .B(new_n347), .C1(new_n358), .C2(new_n359), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n338), .B1(new_n342), .B2(new_n336), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(new_n217), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(new_n343), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n357), .A2(G110), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n363), .B(new_n364), .C1(new_n353), .C2(new_n352), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n360), .A2(new_n365), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n335), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n334), .B1(new_n360), .B2(new_n365), .ZN(new_n368));
  OR2_X1    g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n369), .A2(KEYINPUT25), .A3(new_n189), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n189), .B1(new_n367), .B2(new_n368), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT25), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n327), .B1(new_n370), .B2(new_n373), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n326), .A2(G902), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n374), .B1(new_n369), .B2(new_n375), .ZN(new_n376));
  AND2_X1   g190(.A1(new_n324), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n191), .A2(G227), .ZN(new_n378));
  XOR2_X1   g192(.A(G110), .B(G140), .Z(new_n379));
  XNOR2_X1  g193(.A(new_n378), .B(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT84), .ZN(new_n381));
  INV_X1    g195(.A(G101), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT3), .ZN(new_n383));
  INV_X1    g197(.A(G104), .ZN(new_n384));
  AOI22_X1  g198(.A1(KEYINPUT80), .A2(new_n383), .B1(new_n384), .B2(G107), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT80), .ZN(new_n386));
  INV_X1    g200(.A(G107), .ZN(new_n387));
  AND4_X1   g201(.A1(new_n386), .A2(new_n387), .A3(KEYINPUT3), .A4(G104), .ZN(new_n388));
  AOI22_X1  g202(.A1(new_n386), .A2(KEYINPUT3), .B1(new_n387), .B2(G104), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n382), .B(new_n385), .C1(new_n388), .C2(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n241), .B1(new_n218), .B2(KEYINPUT1), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n243), .B1(new_n391), .B2(new_n214), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n384), .A2(G107), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n387), .A2(G104), .ZN(new_n394));
  OAI21_X1  g208(.A(G101), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n390), .A2(new_n392), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(KEYINPUT82), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT82), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n390), .A2(new_n392), .A3(new_n398), .A4(new_n395), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  XNOR2_X1  g214(.A(KEYINPUT83), .B(KEYINPUT10), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n390), .A2(new_n395), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n269), .A2(KEYINPUT10), .A3(new_n404), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n385), .B1(new_n388), .B2(new_n389), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(G101), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT4), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n408), .A2(KEYINPUT81), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n407), .A2(new_n390), .A3(new_n409), .ZN(new_n410));
  OAI211_X1 g224(.A(new_n406), .B(G101), .C1(KEYINPUT81), .C2(new_n408), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n410), .A2(new_n228), .A3(new_n411), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n402), .A2(new_n405), .A3(new_n262), .A4(new_n412), .ZN(new_n413));
  OAI211_X1 g227(.A(new_n243), .B(new_n403), .C1(new_n264), .C2(new_n268), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n400), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(KEYINPUT12), .B1(new_n415), .B2(new_n239), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT12), .ZN(new_n417));
  AOI211_X1 g231(.A(new_n417), .B(new_n262), .C1(new_n400), .C2(new_n414), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n381), .B(new_n413), .C1(new_n416), .C2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  AOI22_X1  g234(.A1(new_n253), .A2(new_n403), .B1(new_n397), .B2(new_n399), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n417), .B1(new_n421), .B2(new_n262), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n415), .A2(KEYINPUT12), .A3(new_n239), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n381), .B1(new_n424), .B2(new_n413), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n380), .B1(new_n420), .B2(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n402), .A2(new_n405), .A3(new_n412), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(new_n239), .ZN(new_n428));
  INV_X1    g242(.A(new_n380), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n428), .A2(new_n413), .A3(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n426), .A2(G469), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(G469), .A2(G902), .ZN(new_n432));
  INV_X1    g246(.A(G469), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n413), .A2(new_n429), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n434), .B1(new_n423), .B2(new_n422), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n429), .B1(new_n428), .B2(new_n413), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n433), .B(new_n189), .C1(new_n435), .C2(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n431), .A2(new_n432), .A3(new_n437), .ZN(new_n438));
  XNOR2_X1  g252(.A(KEYINPUT9), .B(G234), .ZN(new_n439));
  OAI21_X1  g253(.A(G221), .B1(new_n439), .B2(G902), .ZN(new_n440));
  AND2_X1   g254(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  OAI21_X1  g255(.A(G214), .B1(G237), .B2(G902), .ZN(new_n442));
  OAI21_X1  g256(.A(G210), .B1(G237), .B2(G902), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n228), .A2(G125), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n445), .B1(new_n253), .B2(G125), .ZN(new_n446));
  INV_X1    g260(.A(G224), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n447), .A2(G953), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  AND2_X1   g263(.A1(new_n449), .A2(KEYINPUT7), .ZN(new_n450));
  OR2_X1    g264(.A1(new_n446), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n212), .A2(new_n410), .A3(new_n411), .ZN(new_n452));
  INV_X1    g266(.A(new_n205), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n199), .A2(new_n201), .A3(KEYINPUT5), .ZN(new_n454));
  OAI21_X1  g268(.A(G113), .B1(new_n199), .B2(KEYINPUT5), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n453), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(new_n404), .ZN(new_n458));
  XNOR2_X1  g272(.A(G110), .B(G122), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n452), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n446), .A2(new_n450), .ZN(new_n461));
  AND2_X1   g275(.A1(new_n455), .A2(KEYINPUT87), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n454), .B1(new_n455), .B2(KEYINPUT87), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n205), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n404), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n457), .A2(new_n403), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n459), .B(KEYINPUT8), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n451), .A2(new_n460), .A3(new_n461), .A4(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(new_n189), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n460), .A2(KEYINPUT6), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n452), .A2(new_n458), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT85), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n459), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n452), .A2(KEYINPUT85), .A3(new_n458), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n471), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n472), .A2(new_n473), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT6), .ZN(new_n478));
  INV_X1    g292(.A(new_n459), .ZN(new_n479));
  NAND4_X1  g293(.A1(new_n477), .A2(new_n478), .A3(new_n475), .A4(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(KEYINPUT86), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT86), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n474), .A2(new_n482), .A3(new_n478), .A4(new_n475), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n476), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  OR2_X1    g298(.A1(new_n446), .A2(new_n448), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n446), .A2(new_n448), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  AOI211_X1 g302(.A(new_n444), .B(new_n470), .C1(new_n484), .C2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n481), .A2(new_n483), .ZN(new_n490));
  INV_X1    g304(.A(new_n476), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n490), .A2(new_n491), .A3(new_n488), .ZN(new_n492));
  INV_X1    g306(.A(new_n470), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n443), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n442), .B1(new_n489), .B2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  AND2_X1   g310(.A1(new_n441), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT97), .ZN(new_n498));
  INV_X1    g312(.A(G953), .ZN(new_n499));
  INV_X1    g313(.A(G952), .ZN(new_n500));
  AND2_X1   g314(.A1(new_n500), .A2(KEYINPUT96), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n500), .A2(KEYINPUT96), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n499), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n503), .B1(G234), .B2(G237), .ZN(new_n504));
  AOI211_X1 g318(.A(new_n189), .B(new_n191), .C1(G234), .C2(G237), .ZN(new_n505));
  XNOR2_X1  g319(.A(KEYINPUT21), .B(G898), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(G475), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n499), .A2(KEYINPUT70), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT70), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(G953), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n509), .A2(new_n511), .A3(G214), .A4(new_n192), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(new_n219), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n191), .A2(G143), .A3(G214), .A4(new_n192), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(KEYINPUT88), .A2(KEYINPUT18), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n515), .A2(G131), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n342), .A2(G146), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n347), .A2(new_n519), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n513), .B(new_n514), .C1(new_n237), .C2(new_n516), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n518), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n515), .A2(G131), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT17), .ZN(new_n524));
  OAI211_X1 g338(.A(new_n362), .B(new_n343), .C1(new_n523), .C2(new_n524), .ZN(new_n525));
  AND3_X1   g339(.A1(new_n513), .A2(new_n514), .A3(new_n237), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n237), .B1(new_n513), .B2(new_n514), .ZN(new_n527));
  NOR3_X1   g341(.A1(new_n526), .A2(new_n527), .A3(KEYINPUT17), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n522), .B1(new_n525), .B2(new_n528), .ZN(new_n529));
  XNOR2_X1  g343(.A(G113), .B(G122), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n530), .B(new_n384), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n531), .B(new_n522), .C1(new_n525), .C2(new_n528), .ZN(new_n534));
  AOI21_X1  g348(.A(G902), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n508), .B1(new_n535), .B2(KEYINPUT89), .ZN(new_n536));
  INV_X1    g350(.A(new_n534), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n363), .B1(KEYINPUT17), .B2(new_n527), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n513), .A2(new_n514), .A3(new_n237), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n523), .A2(new_n524), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n531), .B1(new_n541), .B2(new_n522), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n189), .B1(new_n537), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT89), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n536), .A2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT20), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT19), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n345), .A2(new_n548), .A3(new_n346), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n342), .A2(KEYINPUT19), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n549), .A2(new_n217), .A3(new_n550), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n551), .B(new_n343), .C1(new_n526), .C2(new_n527), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n522), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(new_n532), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(new_n534), .ZN(new_n555));
  NOR2_X1   g369(.A1(G475), .A2(G902), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n547), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n556), .ZN(new_n558));
  AOI211_X1 g372(.A(KEYINPUT20), .B(new_n558), .C1(new_n554), .C2(new_n534), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n546), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n200), .A2(G122), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n561), .B(KEYINPUT14), .ZN(new_n562));
  INV_X1    g376(.A(G122), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(KEYINPUT90), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT90), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(G122), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n200), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  OAI21_X1  g381(.A(G107), .B1(new_n562), .B2(new_n567), .ZN(new_n568));
  XNOR2_X1  g382(.A(KEYINPUT90), .B(G122), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n387), .B(new_n561), .C1(new_n569), .C2(new_n200), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n219), .A2(G128), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n241), .A2(G143), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n573), .A2(G134), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n230), .B1(new_n571), .B2(new_n572), .ZN(new_n575));
  OAI211_X1 g389(.A(new_n568), .B(new_n570), .C1(new_n574), .C2(new_n575), .ZN(new_n576));
  NOR3_X1   g390(.A1(new_n439), .A2(new_n325), .A3(G953), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT13), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n578), .B1(new_n241), .B2(G143), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(KEYINPUT92), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT92), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n571), .A2(new_n581), .A3(new_n578), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n219), .A2(KEYINPUT13), .A3(G128), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n580), .A2(new_n582), .A3(new_n572), .A4(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n574), .B1(new_n584), .B2(G134), .ZN(new_n585));
  INV_X1    g399(.A(new_n561), .ZN(new_n586));
  OAI21_X1  g400(.A(G107), .B1(new_n567), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n587), .A2(KEYINPUT91), .A3(new_n570), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(KEYINPUT91), .B1(new_n587), .B2(new_n570), .ZN(new_n590));
  OAI211_X1 g404(.A(new_n576), .B(new_n577), .C1(new_n589), .C2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n587), .A2(new_n570), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT91), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n595), .A2(new_n588), .A3(new_n585), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n577), .B1(new_n596), .B2(new_n576), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n189), .B1(new_n592), .B2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT93), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(G478), .ZN(new_n601));
  NOR2_X1   g415(.A1(KEYINPUT94), .A2(KEYINPUT15), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(KEYINPUT94), .A2(KEYINPUT15), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n601), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  OAI211_X1 g419(.A(KEYINPUT93), .B(new_n189), .C1(new_n592), .C2(new_n597), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n600), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  OR2_X1    g421(.A1(new_n598), .A2(new_n605), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OR2_X1    g423(.A1(new_n609), .A2(KEYINPUT95), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(KEYINPUT95), .ZN(new_n611));
  AOI211_X1 g425(.A(new_n507), .B(new_n560), .C1(new_n610), .C2(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n497), .A2(new_n498), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n497), .A2(new_n612), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(KEYINPUT97), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n377), .A2(new_n613), .A3(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(KEYINPUT98), .B(G101), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G3));
  NAND2_X1  g432(.A1(new_n441), .A2(new_n376), .ZN(new_n619));
  OAI21_X1  g433(.A(G472), .B1(new_n306), .B2(G902), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n620), .B1(new_n306), .B2(new_n190), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n600), .A2(new_n601), .A3(new_n606), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n596), .A2(new_n576), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n577), .B(KEYINPUT99), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n592), .B1(new_n626), .B2(KEYINPUT100), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n627), .B1(KEYINPUT100), .B2(new_n626), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(KEYINPUT33), .ZN(new_n629));
  OR3_X1    g443(.A1(new_n592), .A2(new_n597), .A3(KEYINPUT33), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n189), .A2(G478), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n623), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n560), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n495), .A2(new_n635), .A3(new_n507), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n622), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(KEYINPUT34), .B(G104), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G6));
  NAND2_X1  g453(.A1(new_n610), .A2(new_n611), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT101), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n641), .B1(new_n557), .B2(new_n559), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n531), .B1(new_n552), .B2(new_n522), .ZN(new_n643));
  AND2_X1   g457(.A1(new_n520), .A2(new_n521), .ZN(new_n644));
  AOI22_X1  g458(.A1(new_n538), .A2(new_n540), .B1(new_n644), .B2(new_n518), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n643), .B1(new_n645), .B2(new_n531), .ZN(new_n646));
  OAI21_X1  g460(.A(KEYINPUT20), .B1(new_n646), .B2(new_n558), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n555), .A2(new_n547), .A3(new_n556), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n647), .A2(KEYINPUT101), .A3(new_n648), .ZN(new_n649));
  AOI22_X1  g463(.A1(new_n642), .A2(new_n649), .B1(new_n545), .B2(new_n536), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NOR4_X1   g465(.A1(new_n495), .A2(new_n640), .A3(new_n507), .A4(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n622), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(KEYINPUT102), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT35), .B(G107), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G9));
  OR2_X1    g470(.A1(new_n334), .A2(KEYINPUT36), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(new_n366), .ZN(new_n658));
  NOR3_X1   g472(.A1(new_n658), .A2(G902), .A3(new_n326), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n374), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n621), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n615), .A2(new_n613), .A3(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT37), .B(G110), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(KEYINPUT103), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n662), .B(new_n664), .ZN(G12));
  INV_X1    g479(.A(G900), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n504), .B1(new_n505), .B2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  NOR3_X1   g482(.A1(new_n557), .A2(new_n559), .A3(new_n641), .ZN(new_n669));
  AOI21_X1  g483(.A(KEYINPUT101), .B1(new_n647), .B2(new_n648), .ZN(new_n670));
  OAI211_X1 g484(.A(new_n546), .B(new_n668), .C1(new_n669), .C2(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n640), .A2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n660), .ZN(new_n673));
  AND3_X1   g487(.A1(new_n441), .A2(new_n496), .A3(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n324), .A2(new_n672), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G128), .ZN(G30));
  XOR2_X1   g490(.A(new_n667), .B(KEYINPUT39), .Z(new_n677));
  NAND2_X1  g491(.A1(new_n441), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g492(.A(new_n678), .B(KEYINPUT40), .Z(new_n679));
  NOR2_X1   g493(.A1(new_n292), .A2(new_n302), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n189), .B1(new_n313), .B2(new_n197), .ZN(new_n681));
  OAI21_X1  g495(.A(G472), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n309), .A2(new_n323), .A3(new_n682), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n489), .A2(new_n494), .ZN(new_n684));
  XOR2_X1   g498(.A(new_n684), .B(KEYINPUT38), .Z(new_n685));
  NAND3_X1  g499(.A1(new_n610), .A2(new_n611), .A3(new_n560), .ZN(new_n686));
  INV_X1    g500(.A(new_n442), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n686), .A2(new_n673), .A3(new_n687), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n679), .A2(new_n683), .A3(new_n685), .A4(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G143), .ZN(G45));
  NOR2_X1   g504(.A1(new_n635), .A2(new_n667), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n324), .A2(new_n674), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G146), .ZN(G48));
  NOR2_X1   g507(.A1(new_n435), .A2(new_n436), .ZN(new_n694));
  OAI21_X1  g508(.A(G469), .B1(new_n694), .B2(G902), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n695), .A2(new_n440), .A3(new_n437), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n324), .A2(new_n636), .A3(new_n376), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(KEYINPUT41), .B(G113), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(G15));
  NAND4_X1  g514(.A1(new_n324), .A2(new_n652), .A3(new_n376), .A4(new_n697), .ZN(new_n701));
  AND2_X1   g515(.A1(new_n701), .A2(KEYINPUT104), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n701), .A2(KEYINPUT104), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(new_n200), .ZN(G18));
  NOR3_X1   g519(.A1(new_n495), .A2(new_n660), .A3(new_n696), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n324), .A2(new_n612), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G119), .ZN(G21));
  NOR2_X1   g522(.A1(new_n495), .A2(new_n686), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n696), .A2(new_n507), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n294), .B1(new_n197), .B2(new_n314), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n712), .A2(new_n188), .A3(new_n189), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n713), .A2(new_n376), .A3(new_n620), .ZN(new_n714));
  OAI21_X1  g528(.A(KEYINPUT105), .B1(new_n711), .B2(new_n714), .ZN(new_n715));
  AND3_X1   g529(.A1(new_n713), .A2(new_n376), .A3(new_n620), .ZN(new_n716));
  NOR4_X1   g530(.A1(new_n495), .A2(new_n686), .A3(new_n696), .A4(new_n507), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT105), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n716), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n715), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G122), .ZN(G24));
  AND2_X1   g535(.A1(new_n713), .A2(new_n620), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n722), .A2(new_n691), .A3(new_n706), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G125), .ZN(G27));
  XOR2_X1   g538(.A(new_n432), .B(KEYINPUT106), .Z(new_n725));
  NAND3_X1  g539(.A1(new_n431), .A2(new_n437), .A3(new_n725), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n726), .A2(KEYINPUT107), .A3(new_n440), .ZN(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  AOI21_X1  g542(.A(KEYINPUT107), .B1(new_n726), .B2(new_n440), .ZN(new_n729));
  AOI211_X1 g543(.A(new_n487), .B(new_n476), .C1(new_n481), .C2(new_n483), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n444), .B1(new_n730), .B2(new_n470), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n492), .A2(new_n443), .A3(new_n493), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n731), .A2(new_n442), .A3(new_n732), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n728), .A2(new_n729), .A3(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n324), .A2(new_n376), .A3(new_n691), .A4(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT42), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT108), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n734), .A2(new_n691), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n304), .A2(KEYINPUT32), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n307), .B1(new_n306), .B2(new_n190), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n740), .A2(new_n317), .A3(new_n741), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n742), .A2(KEYINPUT42), .A3(new_n376), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n738), .B1(new_n739), .B2(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(new_n743), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n745), .A2(KEYINPUT108), .A3(new_n691), .A4(new_n734), .ZN(new_n746));
  AND3_X1   g560(.A1(new_n737), .A2(new_n744), .A3(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(new_n237), .ZN(G33));
  XNOR2_X1  g562(.A(new_n672), .B(KEYINPUT109), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n324), .A2(new_n376), .A3(new_n749), .A4(new_n734), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G134), .ZN(G36));
  AND2_X1   g565(.A1(new_n426), .A2(new_n430), .ZN(new_n752));
  OR2_X1    g566(.A1(new_n752), .A2(KEYINPUT45), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(KEYINPUT45), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n753), .A2(G469), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(new_n725), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT46), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n755), .A2(KEYINPUT46), .A3(new_n725), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n758), .A2(new_n437), .A3(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n760), .A2(new_n440), .A3(new_n677), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT110), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n760), .A2(KEYINPUT110), .A3(new_n440), .A4(new_n677), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(new_n765), .ZN(new_n766));
  OR2_X1    g580(.A1(new_n560), .A2(KEYINPUT111), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n560), .A2(KEYINPUT111), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n767), .A2(new_n634), .A3(new_n768), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n560), .A2(KEYINPUT43), .ZN(new_n770));
  AOI22_X1  g584(.A1(new_n769), .A2(KEYINPUT43), .B1(new_n634), .B2(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n771), .A2(new_n621), .A3(new_n673), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT44), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(new_n733), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n775), .B1(new_n772), .B2(new_n773), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n766), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G137), .ZN(G39));
  INV_X1    g593(.A(new_n376), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n691), .A2(new_n780), .A3(new_n775), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n324), .A2(new_n781), .ZN(new_n782));
  AND3_X1   g596(.A1(new_n760), .A2(KEYINPUT47), .A3(new_n440), .ZN(new_n783));
  AOI21_X1  g597(.A(KEYINPUT47), .B1(new_n760), .B2(new_n440), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n782), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G140), .ZN(G42));
  OR2_X1    g600(.A1(new_n683), .A2(new_n780), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n695), .A2(new_n437), .ZN(new_n788));
  XOR2_X1   g602(.A(new_n788), .B(KEYINPUT49), .Z(new_n789));
  INV_X1    g603(.A(new_n440), .ZN(new_n790));
  OR3_X1    g604(.A1(new_n769), .A2(new_n687), .A3(new_n790), .ZN(new_n791));
  OR4_X1    g605(.A1(new_n685), .A2(new_n787), .A3(new_n789), .A4(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n742), .A2(new_n376), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n697), .A2(new_n504), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n795), .A2(new_n775), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n794), .A2(new_n771), .A3(new_n796), .ZN(new_n797));
  XOR2_X1   g611(.A(new_n797), .B(KEYINPUT48), .Z(new_n798));
  INV_X1    g612(.A(new_n796), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n787), .A2(new_n799), .A3(new_n635), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n771), .A2(new_n716), .A3(new_n504), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n801), .A2(new_n496), .A3(new_n697), .ZN(new_n802));
  NOR4_X1   g616(.A1(new_n798), .A2(new_n503), .A3(new_n800), .A4(new_n802), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n788), .A2(new_n790), .ZN(new_n804));
  OR3_X1    g618(.A1(new_n783), .A2(new_n784), .A3(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n805), .A2(new_n775), .A3(new_n801), .ZN(new_n806));
  OR4_X1    g620(.A1(new_n560), .A2(new_n787), .A3(new_n634), .A4(new_n799), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n796), .A2(new_n673), .A3(new_n722), .A4(new_n771), .ZN(new_n808));
  XOR2_X1   g622(.A(new_n808), .B(KEYINPUT119), .Z(new_n809));
  NOR3_X1   g623(.A1(new_n685), .A2(new_n442), .A3(new_n696), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(new_n801), .ZN(new_n811));
  XOR2_X1   g625(.A(new_n811), .B(KEYINPUT50), .Z(new_n812));
  NAND4_X1  g626(.A1(new_n806), .A2(new_n807), .A3(new_n809), .A4(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT51), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n803), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n495), .A2(new_n507), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n609), .A2(KEYINPUT113), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT113), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n607), .A2(new_n608), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(new_n820), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n635), .B1(new_n560), .B2(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n622), .A2(new_n816), .A3(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n616), .A2(new_n662), .A3(new_n823), .ZN(new_n824));
  AND3_X1   g638(.A1(new_n698), .A2(new_n720), .A3(new_n707), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n825), .B1(new_n702), .B2(new_n703), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n824), .B1(new_n826), .B2(KEYINPUT112), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT112), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n825), .B(new_n828), .C1(new_n702), .C2(new_n703), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT53), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n820), .A2(new_n671), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n832), .A2(new_n684), .A3(KEYINPUT114), .A4(new_n442), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT114), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n650), .A2(new_n817), .A3(new_n668), .A4(new_n819), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n834), .B1(new_n733), .B2(new_n835), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n438), .A2(new_n673), .A3(new_n440), .ZN(new_n837));
  AND3_X1   g651(.A1(new_n833), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n324), .A2(new_n838), .A3(KEYINPUT115), .ZN(new_n839));
  AOI21_X1  g653(.A(KEYINPUT115), .B1(new_n324), .B2(new_n838), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n734), .A2(new_n673), .A3(new_n691), .A4(new_n722), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n750), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g657(.A(KEYINPUT116), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n750), .A2(new_n842), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n324), .A2(new_n838), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT115), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n324), .A2(new_n838), .A3(KEYINPUT115), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT116), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n845), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n747), .B1(new_n844), .B2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT118), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n854), .B1(new_n673), .B2(new_n667), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n660), .A2(KEYINPUT118), .A3(new_n668), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n709), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n683), .A2(new_n440), .A3(new_n857), .A4(new_n726), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n858), .A2(new_n675), .A3(new_n692), .A4(new_n723), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n859), .A2(KEYINPUT52), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n675), .A2(new_n723), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(KEYINPUT117), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT117), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n675), .A2(new_n863), .A3(new_n723), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n862), .A2(new_n692), .A3(new_n858), .A4(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n860), .B1(new_n865), .B2(KEYINPUT52), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n830), .A2(new_n831), .A3(new_n853), .A4(new_n866), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n859), .A2(KEYINPUT52), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n868), .A2(new_n860), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n827), .A2(new_n853), .A3(new_n829), .A4(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(KEYINPUT53), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n867), .A2(KEYINPUT54), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n870), .A2(new_n831), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT54), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n826), .A2(new_n831), .A3(new_n824), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n875), .A2(new_n866), .A3(new_n853), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n873), .A2(new_n874), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n872), .A2(new_n877), .ZN(new_n878));
  AOI211_X1 g692(.A(new_n815), .B(new_n878), .C1(new_n814), .C2(new_n813), .ZN(new_n879));
  NOR2_X1   g693(.A1(G952), .A2(G953), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n792), .B1(new_n879), .B2(new_n880), .ZN(G75));
  XNOR2_X1  g695(.A(new_n484), .B(KEYINPUT120), .ZN(new_n882));
  XOR2_X1   g696(.A(new_n882), .B(KEYINPUT55), .Z(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n189), .B1(new_n873), .B2(new_n876), .ZN(new_n885));
  AOI211_X1 g699(.A(KEYINPUT56), .B(new_n487), .C1(new_n885), .C2(G210), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n873), .A2(new_n876), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n887), .A2(G210), .A3(G902), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT56), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n488), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n884), .B1(new_n886), .B2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(G210), .ZN(new_n892));
  AOI211_X1 g706(.A(new_n892), .B(new_n189), .C1(new_n873), .C2(new_n876), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n487), .B1(new_n893), .B2(KEYINPUT56), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n888), .A2(new_n889), .A3(new_n488), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n894), .A2(new_n895), .A3(new_n883), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n191), .A2(G952), .ZN(new_n897));
  INV_X1    g711(.A(new_n897), .ZN(new_n898));
  AND3_X1   g712(.A1(new_n891), .A2(new_n896), .A3(new_n898), .ZN(G51));
  XOR2_X1   g713(.A(new_n725), .B(KEYINPUT57), .Z(new_n900));
  AND3_X1   g714(.A1(new_n873), .A2(new_n874), .A3(new_n876), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n874), .B1(new_n873), .B2(new_n876), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n900), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n694), .B1(new_n903), .B2(KEYINPUT121), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT121), .ZN(new_n905));
  OAI211_X1 g719(.A(new_n905), .B(new_n900), .C1(new_n901), .C2(new_n902), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n885), .A2(G469), .A3(new_n754), .A4(new_n753), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n897), .B1(new_n907), .B2(new_n908), .ZN(G54));
  AND3_X1   g723(.A1(new_n885), .A2(KEYINPUT58), .A3(G475), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n898), .B1(new_n910), .B2(new_n555), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n911), .B1(new_n555), .B2(new_n910), .ZN(G60));
  NAND2_X1  g726(.A1(G478), .A2(G902), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n913), .B(KEYINPUT59), .Z(new_n914));
  AOI21_X1  g728(.A(new_n914), .B1(new_n872), .B2(new_n877), .ZN(new_n915));
  OR3_X1    g729(.A1(new_n915), .A2(KEYINPUT122), .A3(new_n631), .ZN(new_n916));
  OAI21_X1  g730(.A(KEYINPUT122), .B1(new_n915), .B2(new_n631), .ZN(new_n917));
  OR2_X1    g731(.A1(new_n901), .A2(new_n902), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n632), .A2(new_n914), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n897), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  AND3_X1   g734(.A1(new_n916), .A2(new_n917), .A3(new_n920), .ZN(G63));
  NAND2_X1  g735(.A1(G217), .A2(G902), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT60), .ZN(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n887), .A2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(new_n369), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n897), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n925), .A2(KEYINPUT123), .A3(new_n658), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT123), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n923), .B1(new_n873), .B2(new_n876), .ZN(new_n930));
  INV_X1    g744(.A(new_n658), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n929), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n927), .B1(new_n928), .B2(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT61), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  OAI211_X1 g749(.A(KEYINPUT61), .B(new_n927), .C1(new_n928), .C2(new_n932), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(G66));
  OAI21_X1  g751(.A(G953), .B1(new_n506), .B2(new_n447), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n938), .B(KEYINPUT124), .Z(new_n939));
  INV_X1    g753(.A(new_n191), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n939), .B1(new_n830), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n882), .B1(G898), .B2(new_n191), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n941), .B(new_n942), .ZN(G69));
  AND3_X1   g757(.A1(new_n862), .A2(new_n692), .A3(new_n864), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(new_n689), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT62), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n944), .A2(KEYINPUT62), .A3(new_n689), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(new_n678), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n377), .A2(new_n950), .A3(new_n775), .A4(new_n822), .ZN(new_n951));
  AND3_X1   g765(.A1(new_n778), .A2(new_n785), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n949), .A2(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT125), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n949), .A2(new_n952), .A3(KEYINPUT125), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n549), .A2(new_n550), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n291), .B(new_n958), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n957), .A2(new_n191), .A3(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(G227), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n959), .B1(new_n961), .B2(new_n940), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n785), .A2(new_n750), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n794), .A2(new_n709), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n964), .B1(new_n774), .B2(new_n776), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n963), .B1(new_n766), .B2(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(new_n747), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n966), .A2(new_n967), .A3(new_n944), .ZN(new_n968));
  INV_X1    g782(.A(new_n968), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n962), .B1(new_n969), .B2(new_n940), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n666), .B1(new_n959), .B2(new_n961), .ZN(new_n971));
  OAI211_X1 g785(.A(new_n960), .B(new_n970), .C1(new_n191), .C2(new_n971), .ZN(G72));
  NAND3_X1  g786(.A1(new_n955), .A2(new_n830), .A3(new_n956), .ZN(new_n973));
  NAND2_X1  g787(.A1(G472), .A2(G902), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n974), .B(KEYINPUT63), .Z(new_n975));
  NAND2_X1  g789(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(new_n680), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT127), .ZN(new_n978));
  INV_X1    g792(.A(new_n680), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n979), .A2(new_n311), .A3(new_n975), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n980), .B(KEYINPUT126), .Z(new_n981));
  NAND3_X1  g795(.A1(new_n867), .A2(new_n871), .A3(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(new_n830), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n975), .B1(new_n968), .B2(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(new_n311), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n897), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n977), .A2(new_n978), .A3(new_n982), .A4(new_n986), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n979), .B1(new_n973), .B2(new_n975), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n986), .A2(new_n982), .ZN(new_n989));
  OAI21_X1  g803(.A(KEYINPUT127), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n987), .A2(new_n990), .ZN(G57));
endmodule


