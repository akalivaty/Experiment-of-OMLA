//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 1 1 0 1 1 0 0 1 1 0 1 1 1 0 0 0 0 0 0 0 1 1 0 0 1 1 0 0 1 0 0 1 1 1 1 0 1 0 1 1 1 0 0 0 1 1 0 0 0 0 1 0 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n755, new_n756,
    new_n757, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n768, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n836, new_n838, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n889, new_n890, new_n892, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n964, new_n965;
  INV_X1    g000(.A(KEYINPUT72), .ZN(new_n202));
  INV_X1    g001(.A(G227gat), .ZN(new_n203));
  INV_X1    g002(.A(G233gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT69), .ZN(new_n206));
  OR2_X1    g005(.A1(KEYINPUT68), .A2(G183gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(KEYINPUT68), .A2(G183gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n207), .A2(KEYINPUT27), .A3(new_n208), .ZN(new_n209));
  NOR2_X1   g008(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  AOI21_X1  g010(.A(G190gat), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n206), .B1(new_n212), .B2(KEYINPUT28), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT28), .ZN(new_n214));
  AND2_X1   g013(.A1(KEYINPUT68), .A2(G183gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(KEYINPUT68), .A2(G183gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n210), .B1(new_n217), .B2(KEYINPUT27), .ZN(new_n218));
  OAI211_X1 g017(.A(KEYINPUT69), .B(new_n214), .C1(new_n218), .C2(G190gat), .ZN(new_n219));
  XNOR2_X1  g018(.A(KEYINPUT27), .B(G183gat), .ZN(new_n220));
  INV_X1    g019(.A(G190gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n220), .A2(KEYINPUT28), .A3(new_n221), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n213), .A2(new_n219), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(G183gat), .A2(G190gat), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(G169gat), .ZN(new_n226));
  INV_X1    g025(.A(G176gat), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT26), .ZN(new_n229));
  NOR2_X1   g028(.A1(G169gat), .A2(G176gat), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n228), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(new_n230), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(KEYINPUT26), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n225), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n223), .A2(new_n234), .ZN(new_n235));
  XOR2_X1   g034(.A(G127gat), .B(G134gat), .Z(new_n236));
  NOR2_X1   g035(.A1(new_n236), .A2(KEYINPUT1), .ZN(new_n237));
  INV_X1    g036(.A(G120gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(G113gat), .ZN(new_n239));
  XNOR2_X1  g038(.A(KEYINPUT70), .B(G113gat), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n239), .B1(new_n240), .B2(new_n238), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT1), .ZN(new_n242));
  INV_X1    g041(.A(new_n239), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n238), .A2(G113gat), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n242), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  AOI22_X1  g044(.A1(new_n237), .A2(new_n241), .B1(new_n245), .B2(new_n236), .ZN(new_n246));
  XNOR2_X1  g045(.A(KEYINPUT66), .B(KEYINPUT24), .ZN(new_n247));
  OAI21_X1  g046(.A(KEYINPUT67), .B1(new_n247), .B2(new_n225), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT67), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT24), .ZN(new_n250));
  AND2_X1   g049(.A1(new_n250), .A2(KEYINPUT66), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n250), .A2(KEYINPUT66), .ZN(new_n252));
  OAI211_X1 g051(.A(new_n249), .B(new_n224), .C1(new_n251), .C2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n225), .A2(KEYINPUT24), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n207), .A2(new_n208), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(new_n221), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n248), .A2(new_n253), .A3(new_n254), .A4(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n230), .A2(KEYINPUT23), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT23), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n228), .B1(new_n259), .B2(new_n232), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n257), .A2(KEYINPUT25), .A3(new_n258), .A4(new_n260), .ZN(new_n261));
  XOR2_X1   g060(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n262));
  OAI21_X1  g061(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n254), .B1(new_n264), .B2(new_n225), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(new_n260), .ZN(new_n266));
  XNOR2_X1  g065(.A(KEYINPUT65), .B(G176gat), .ZN(new_n267));
  NOR3_X1   g066(.A1(new_n267), .A2(new_n259), .A3(G169gat), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n262), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n261), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n235), .A2(new_n246), .A3(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n246), .B1(new_n235), .B2(new_n270), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n205), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT33), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(G15gat), .B(G43gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n277), .B(G71gat), .ZN(new_n278));
  INV_X1    g077(.A(G99gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n278), .B(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n276), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n274), .A2(KEYINPUT32), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n235), .A2(new_n270), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n237), .A2(new_n241), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n245), .A2(new_n236), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n283), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT34), .ZN(new_n288));
  INV_X1    g087(.A(new_n205), .ZN(new_n289));
  NAND4_X1  g088(.A1(new_n287), .A2(new_n288), .A3(new_n289), .A4(new_n271), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n287), .A2(new_n289), .A3(new_n271), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(KEYINPUT34), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n282), .A2(new_n290), .A3(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n282), .B1(new_n292), .B2(new_n290), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n281), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n292), .A2(new_n290), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n297), .A2(KEYINPUT32), .A3(new_n274), .ZN(new_n298));
  INV_X1    g097(.A(new_n281), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n298), .A2(new_n299), .A3(new_n293), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n202), .B1(new_n296), .B2(new_n300), .ZN(new_n301));
  NOR3_X1   g100(.A1(new_n301), .A2(KEYINPUT71), .A3(KEYINPUT36), .ZN(new_n302));
  NOR3_X1   g101(.A1(new_n294), .A2(new_n295), .A3(new_n281), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n299), .B1(new_n298), .B2(new_n293), .ZN(new_n304));
  OAI21_X1  g103(.A(KEYINPUT71), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  AND2_X1   g104(.A1(new_n305), .A2(KEYINPUT36), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT71), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n303), .A2(new_n304), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n307), .B1(new_n308), .B2(new_n202), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n302), .B1(new_n306), .B2(new_n309), .ZN(new_n310));
  XOR2_X1   g109(.A(G197gat), .B(G204gat), .Z(new_n311));
  INV_X1    g110(.A(KEYINPUT22), .ZN(new_n312));
  INV_X1    g111(.A(G218gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(KEYINPUT73), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT73), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(G218gat), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n314), .A2(new_n316), .A3(G211gat), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n311), .B1(new_n312), .B2(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(G211gat), .B(G218gat), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n319), .A2(KEYINPUT74), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n318), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(KEYINPUT73), .B(G218gat), .ZN(new_n323));
  AOI21_X1  g122(.A(KEYINPUT22), .B1(new_n323), .B2(G211gat), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n320), .B1(new_n324), .B2(new_n311), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n322), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT81), .ZN(new_n327));
  INV_X1    g126(.A(G148gat), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n327), .B1(new_n328), .B2(G141gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(G141gat), .ZN(new_n330));
  INV_X1    g129(.A(G141gat), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n331), .A2(KEYINPUT81), .A3(G148gat), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n329), .A2(new_n330), .A3(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(G155gat), .ZN(new_n334));
  INV_X1    g133(.A(G162gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(G155gat), .A2(G162gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(KEYINPUT2), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(KEYINPUT82), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT82), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n337), .A2(new_n341), .A3(KEYINPUT2), .ZN(new_n342));
  NAND4_X1  g141(.A1(new_n333), .A2(new_n338), .A3(new_n340), .A4(new_n342), .ZN(new_n343));
  XNOR2_X1  g142(.A(G141gat), .B(G148gat), .ZN(new_n344));
  OAI211_X1 g143(.A(new_n337), .B(new_n336), .C1(new_n344), .C2(KEYINPUT2), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(KEYINPUT83), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT29), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT83), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n343), .A2(new_n349), .A3(new_n345), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n326), .A2(new_n347), .A3(new_n348), .A4(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n347), .A2(KEYINPUT3), .A3(new_n350), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n351), .A2(KEYINPUT91), .A3(new_n352), .ZN(new_n353));
  AND3_X1   g152(.A1(new_n343), .A2(new_n349), .A3(new_n345), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n349), .B1(new_n343), .B2(new_n345), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT91), .ZN(new_n357));
  AOI21_X1  g156(.A(KEYINPUT29), .B1(new_n322), .B2(new_n325), .ZN(new_n358));
  OAI211_X1 g157(.A(new_n356), .B(new_n357), .C1(KEYINPUT3), .C2(new_n358), .ZN(new_n359));
  AND2_X1   g158(.A1(new_n322), .A2(new_n325), .ZN(new_n360));
  XOR2_X1   g159(.A(KEYINPUT76), .B(KEYINPUT29), .Z(new_n361));
  OAI21_X1  g160(.A(new_n361), .B1(new_n346), .B2(KEYINPUT3), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT92), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT92), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n360), .A2(new_n362), .A3(new_n365), .ZN(new_n366));
  NAND4_X1  g165(.A1(new_n353), .A2(new_n359), .A3(new_n364), .A4(new_n366), .ZN(new_n367));
  AND2_X1   g166(.A1(G228gat), .A2(G233gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT3), .ZN(new_n370));
  INV_X1    g169(.A(new_n319), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n361), .B1(new_n318), .B2(new_n371), .ZN(new_n372));
  NOR3_X1   g171(.A1(new_n324), .A2(new_n319), .A3(new_n311), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n370), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT85), .ZN(new_n375));
  AND3_X1   g174(.A1(new_n343), .A2(new_n375), .A3(new_n345), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n375), .B1(new_n343), .B2(new_n345), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n374), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n368), .B1(new_n360), .B2(new_n362), .ZN(new_n380));
  AND2_X1   g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n369), .A2(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(G78gat), .B(G106gat), .ZN(new_n384));
  XOR2_X1   g183(.A(new_n384), .B(KEYINPUT90), .Z(new_n385));
  NAND2_X1  g184(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(KEYINPUT31), .B(G50gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n387), .B(G22gat), .ZN(new_n388));
  INV_X1    g187(.A(new_n385), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n369), .A2(new_n382), .A3(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n386), .A2(new_n388), .A3(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n388), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n389), .B1(new_n369), .B2(new_n382), .ZN(new_n393));
  AOI211_X1 g192(.A(new_n385), .B(new_n381), .C1(new_n367), .C2(new_n368), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n392), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n391), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n352), .A2(KEYINPUT84), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT84), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n347), .A2(new_n399), .A3(KEYINPUT3), .A4(new_n350), .ZN(new_n400));
  AND2_X1   g199(.A1(new_n343), .A2(new_n345), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(new_n370), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n398), .A2(new_n400), .A3(new_n286), .A4(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT4), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n404), .B(new_n246), .C1(new_n376), .C2(new_n377), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n401), .A2(new_n246), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  OAI211_X1 g206(.A(new_n405), .B(KEYINPUT89), .C1(new_n407), .C2(new_n404), .ZN(new_n408));
  OAI211_X1 g207(.A(new_n403), .B(new_n408), .C1(KEYINPUT89), .C2(new_n405), .ZN(new_n409));
  NAND2_X1  g208(.A1(G225gat), .A2(G233gat), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT5), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  OR2_X1    g211(.A1(new_n409), .A2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT87), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n406), .A2(new_n404), .ZN(new_n415));
  OAI211_X1 g214(.A(KEYINPUT4), .B(new_n246), .C1(new_n376), .C2(new_n377), .ZN(new_n416));
  AND3_X1   g215(.A1(new_n415), .A2(new_n416), .A3(new_n410), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n347), .A2(new_n350), .A3(new_n286), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n410), .B1(new_n418), .B2(new_n406), .ZN(new_n419));
  OAI21_X1  g218(.A(KEYINPUT86), .B1(new_n419), .B2(new_n411), .ZN(new_n420));
  INV_X1    g219(.A(new_n410), .ZN(new_n421));
  NOR3_X1   g220(.A1(new_n354), .A2(new_n355), .A3(new_n246), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n421), .B1(new_n422), .B2(new_n407), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT86), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n423), .A2(new_n424), .A3(KEYINPUT5), .ZN(new_n425));
  AOI221_X4 g224(.A(new_n414), .B1(new_n403), .B2(new_n417), .C1(new_n420), .C2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n420), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n403), .A2(new_n417), .ZN(new_n428));
  AOI21_X1  g227(.A(KEYINPUT87), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n413), .B1(new_n426), .B2(new_n429), .ZN(new_n430));
  XNOR2_X1  g229(.A(KEYINPUT88), .B(KEYINPUT0), .ZN(new_n431));
  XNOR2_X1  g230(.A(G57gat), .B(G85gat), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n431), .B(new_n432), .ZN(new_n433));
  XNOR2_X1  g232(.A(G1gat), .B(G29gat), .ZN(new_n434));
  XOR2_X1   g233(.A(new_n433), .B(new_n434), .Z(new_n435));
  NAND2_X1  g234(.A1(new_n430), .A2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT6), .ZN(new_n437));
  INV_X1    g236(.A(new_n435), .ZN(new_n438));
  OAI211_X1 g237(.A(new_n413), .B(new_n438), .C1(new_n426), .C2(new_n429), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n436), .A2(new_n437), .A3(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n430), .A2(KEYINPUT6), .A3(new_n435), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT77), .ZN(new_n444));
  NAND2_X1  g243(.A1(G226gat), .A2(G233gat), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT75), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n283), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n235), .A2(KEYINPUT75), .A3(new_n270), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n445), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(KEYINPUT29), .B1(new_n235), .B2(new_n270), .ZN(new_n450));
  INV_X1    g249(.A(new_n445), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n326), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n444), .B1(new_n449), .B2(new_n452), .ZN(new_n453));
  AND2_X1   g252(.A1(new_n361), .A2(new_n445), .ZN(new_n454));
  AND3_X1   g253(.A1(new_n235), .A2(KEYINPUT75), .A3(new_n270), .ZN(new_n455));
  AOI21_X1  g254(.A(KEYINPUT75), .B1(new_n235), .B2(new_n270), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n454), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n235), .A2(new_n451), .A3(new_n270), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n457), .A2(new_n360), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n283), .A2(new_n348), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n360), .B1(new_n460), .B2(new_n445), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n451), .B1(new_n455), .B2(new_n456), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n461), .A2(new_n462), .A3(KEYINPUT77), .ZN(new_n463));
  AND3_X1   g262(.A1(new_n453), .A2(new_n459), .A3(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT79), .ZN(new_n465));
  XNOR2_X1  g264(.A(G8gat), .B(G36gat), .ZN(new_n466));
  XNOR2_X1  g265(.A(G64gat), .B(G92gat), .ZN(new_n467));
  XNOR2_X1  g266(.A(new_n466), .B(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n464), .A2(new_n465), .A3(KEYINPUT30), .A4(new_n469), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n453), .A2(new_n463), .A3(new_n469), .A4(new_n459), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT30), .ZN(new_n472));
  OAI21_X1  g271(.A(KEYINPUT79), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n453), .A2(new_n463), .A3(new_n459), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT78), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n453), .A2(new_n463), .A3(KEYINPUT78), .A4(new_n459), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(new_n468), .ZN(new_n480));
  NOR3_X1   g279(.A1(new_n449), .A2(new_n452), .A3(new_n444), .ZN(new_n481));
  AOI21_X1  g280(.A(KEYINPUT77), .B1(new_n461), .B2(new_n462), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n483), .A2(KEYINPUT80), .A3(new_n469), .A4(new_n459), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT80), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n471), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n484), .A2(new_n472), .A3(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n474), .A2(new_n480), .A3(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n397), .B1(new_n443), .B2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT37), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n453), .A2(new_n463), .A3(new_n490), .A4(new_n459), .ZN(new_n491));
  AND2_X1   g290(.A1(new_n491), .A2(new_n468), .ZN(new_n492));
  OAI211_X1 g291(.A(new_n462), .B(new_n360), .C1(new_n451), .C2(new_n450), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n457), .A2(new_n326), .A3(new_n458), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n493), .A2(KEYINPUT37), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(KEYINPUT38), .B1(new_n492), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n491), .A2(new_n468), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n497), .B1(new_n479), .B2(KEYINPUT37), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n496), .B1(new_n498), .B2(KEYINPUT38), .ZN(new_n499));
  XNOR2_X1  g298(.A(new_n471), .B(KEYINPUT80), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  NOR3_X1   g300(.A1(new_n499), .A2(new_n442), .A3(new_n501), .ZN(new_n502));
  AND3_X1   g301(.A1(new_n474), .A2(new_n480), .A3(new_n487), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT39), .ZN(new_n504));
  NOR3_X1   g303(.A1(new_n422), .A2(new_n421), .A3(new_n407), .ZN(new_n505));
  AOI211_X1 g304(.A(new_n504), .B(new_n505), .C1(new_n409), .C2(new_n421), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n409), .A2(new_n504), .A3(new_n421), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(new_n438), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  OR2_X1    g308(.A1(new_n509), .A2(KEYINPUT40), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(KEYINPUT40), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n510), .A2(new_n436), .A3(new_n511), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n396), .B1(new_n503), .B2(new_n512), .ZN(new_n513));
  OAI211_X1 g312(.A(new_n310), .B(new_n489), .C1(new_n502), .C2(new_n513), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n469), .B1(new_n477), .B2(new_n478), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n515), .B1(new_n500), .B2(new_n472), .ZN(new_n516));
  AND3_X1   g315(.A1(new_n396), .A2(new_n296), .A3(new_n300), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n516), .A2(new_n442), .A3(new_n474), .A4(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT35), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n503), .A2(KEYINPUT35), .A3(new_n442), .A4(new_n517), .ZN(new_n521));
  AND2_X1   g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n514), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(G230gat), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n524), .A2(new_n204), .ZN(new_n525));
  XOR2_X1   g324(.A(G57gat), .B(G64gat), .Z(new_n526));
  INV_X1    g325(.A(G71gat), .ZN(new_n527));
  INV_X1    g326(.A(G78gat), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT9), .ZN(new_n530));
  NOR3_X1   g329(.A1(new_n530), .A2(G71gat), .A3(G78gat), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n526), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(G57gat), .B(G64gat), .ZN(new_n533));
  OAI22_X1  g332(.A1(new_n533), .A2(new_n530), .B1(new_n527), .B2(new_n528), .ZN(new_n534));
  NOR2_X1   g333(.A1(G71gat), .A2(G78gat), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n535), .B(KEYINPUT101), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n532), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n537), .B(KEYINPUT102), .ZN(new_n538));
  INV_X1    g337(.A(G85gat), .ZN(new_n539));
  INV_X1    g338(.A(G92gat), .ZN(new_n540));
  OAI21_X1  g339(.A(KEYINPUT107), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT107), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n542), .A2(G85gat), .A3(G92gat), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n541), .A2(new_n543), .A3(KEYINPUT7), .ZN(new_n544));
  NAND2_X1  g343(.A1(G99gat), .A2(G106gat), .ZN(new_n545));
  AOI22_X1  g344(.A1(KEYINPUT8), .A2(new_n545), .B1(new_n539), .B2(new_n540), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT7), .ZN(new_n547));
  OAI211_X1 g346(.A(KEYINPUT107), .B(new_n547), .C1(new_n539), .C2(new_n540), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n544), .A2(new_n546), .A3(new_n548), .ZN(new_n549));
  XOR2_X1   g348(.A(G99gat), .B(G106gat), .Z(new_n550));
  OR3_X1    g349(.A1(new_n549), .A2(KEYINPUT108), .A3(new_n550), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n549), .A2(new_n550), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n549), .A2(new_n550), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n553), .A2(KEYINPUT108), .A3(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n538), .A2(new_n551), .A3(new_n555), .ZN(new_n556));
  XOR2_X1   g355(.A(KEYINPUT109), .B(KEYINPUT10), .Z(new_n557));
  NOR2_X1   g356(.A1(new_n552), .A2(new_n537), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(new_n554), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n556), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n555), .A2(new_n551), .ZN(new_n561));
  XOR2_X1   g360(.A(new_n537), .B(KEYINPUT102), .Z(new_n562));
  NAND3_X1  g361(.A1(new_n561), .A2(new_n562), .A3(KEYINPUT10), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n525), .B1(new_n560), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n556), .A2(new_n559), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n564), .B1(new_n525), .B2(new_n565), .ZN(new_n566));
  XOR2_X1   g365(.A(G120gat), .B(G148gat), .Z(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(G204gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(KEYINPUT110), .B(G176gat), .ZN(new_n569));
  XOR2_X1   g368(.A(new_n568), .B(new_n569), .Z(new_n570));
  OR2_X1    g369(.A1(new_n566), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n564), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n565), .A2(new_n525), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n572), .A2(new_n573), .A3(new_n570), .ZN(new_n574));
  AND2_X1   g373(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n523), .A2(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(G113gat), .B(G141gat), .ZN(new_n577));
  INV_X1    g376(.A(G197gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n577), .B(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(KEYINPUT11), .B(G169gat), .ZN(new_n580));
  XOR2_X1   g379(.A(new_n579), .B(new_n580), .Z(new_n581));
  XOR2_X1   g380(.A(new_n581), .B(KEYINPUT12), .Z(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT99), .ZN(new_n584));
  XNOR2_X1  g383(.A(G15gat), .B(G22gat), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT16), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n585), .B1(new_n586), .B2(G1gat), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n587), .B1(G1gat), .B2(new_n585), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(G8gat), .ZN(new_n589));
  INV_X1    g388(.A(G43gat), .ZN(new_n590));
  OAI21_X1  g389(.A(KEYINPUT15), .B1(new_n590), .B2(G50gat), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n591), .B1(new_n590), .B2(G50gat), .ZN(new_n592));
  OR3_X1    g391(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n593));
  OAI21_X1  g392(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n592), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  XOR2_X1   g394(.A(KEYINPUT95), .B(G36gat), .Z(new_n596));
  XNOR2_X1  g395(.A(KEYINPUT94), .B(G29gat), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n590), .A2(G50gat), .ZN(new_n599));
  XOR2_X1   g398(.A(KEYINPUT96), .B(G50gat), .Z(new_n600));
  AOI21_X1  g399(.A(new_n599), .B1(new_n600), .B2(new_n590), .ZN(new_n601));
  OAI211_X1 g400(.A(new_n595), .B(new_n598), .C1(KEYINPUT15), .C2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT93), .ZN(new_n603));
  AND2_X1   g402(.A1(new_n593), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n594), .B1(new_n593), .B2(new_n603), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n598), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(new_n592), .ZN(new_n607));
  AND2_X1   g406(.A1(new_n602), .A2(new_n607), .ZN(new_n608));
  OR2_X1    g407(.A1(KEYINPUT97), .A2(KEYINPUT17), .ZN(new_n609));
  NAND2_X1  g408(.A1(KEYINPUT97), .A2(KEYINPUT17), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n602), .A2(new_n607), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n612), .A2(KEYINPUT97), .A3(KEYINPUT17), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n589), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT18), .ZN(new_n615));
  INV_X1    g414(.A(new_n589), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n608), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(G229gat), .A2(G233gat), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NOR4_X1   g418(.A1(new_n614), .A2(new_n615), .A3(new_n617), .A4(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n616), .B(new_n612), .ZN(new_n621));
  XNOR2_X1  g420(.A(KEYINPUT98), .B(KEYINPUT13), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(new_n618), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n584), .B1(new_n620), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n611), .A2(new_n613), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n617), .B1(new_n627), .B2(new_n616), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(new_n618), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(new_n615), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n626), .A2(new_n630), .ZN(new_n631));
  NOR3_X1   g430(.A1(new_n620), .A2(new_n584), .A3(new_n625), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n583), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  AOI21_X1  g432(.A(KEYINPUT18), .B1(new_n628), .B2(new_n618), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n583), .B1(new_n634), .B2(KEYINPUT100), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n620), .A2(new_n625), .ZN(new_n636));
  OAI211_X1 g435(.A(new_n635), .B(new_n636), .C1(KEYINPUT100), .C2(new_n634), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n640));
  OR2_X1    g439(.A1(new_n562), .A2(KEYINPUT21), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(KEYINPUT103), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n589), .B1(new_n562), .B2(KEYINPUT21), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(G183gat), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT103), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n641), .B(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(G183gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n643), .B(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  NAND4_X1  g449(.A1(new_n645), .A2(new_n650), .A3(G231gat), .A4(G233gat), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  AOI22_X1  g451(.A1(new_n645), .A2(new_n650), .B1(G231gat), .B2(G233gat), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n640), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(KEYINPUT104), .B(KEYINPUT105), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(G211gat), .ZN(new_n656));
  XOR2_X1   g455(.A(G127gat), .B(G155gat), .Z(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n645), .A2(new_n650), .ZN(new_n659));
  INV_X1    g458(.A(G231gat), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n659), .B1(new_n660), .B2(new_n204), .ZN(new_n661));
  INV_X1    g460(.A(new_n640), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n661), .A2(new_n662), .A3(new_n651), .ZN(new_n663));
  AND3_X1   g462(.A1(new_n654), .A2(new_n658), .A3(new_n663), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n658), .B1(new_n654), .B2(new_n663), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(G134gat), .B(G162gat), .ZN(new_n668));
  AOI21_X1  g467(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n669));
  XOR2_X1   g468(.A(new_n668), .B(new_n669), .Z(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n627), .A2(new_n551), .A3(new_n555), .ZN(new_n672));
  NAND3_X1  g471(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n561), .A2(new_n612), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n672), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(KEYINPUT106), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n675), .A2(KEYINPUT106), .ZN(new_n678));
  XNOR2_X1  g477(.A(G190gat), .B(G218gat), .ZN(new_n679));
  NOR3_X1   g478(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n679), .ZN(new_n681));
  OR2_X1    g480(.A1(new_n675), .A2(KEYINPUT106), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n681), .B1(new_n682), .B2(new_n676), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n671), .B1(new_n680), .B2(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n679), .B1(new_n677), .B2(new_n678), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n682), .A2(new_n681), .A3(new_n676), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n685), .A2(new_n670), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  NOR4_X1   g487(.A1(new_n576), .A2(new_n639), .A3(new_n667), .A4(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(new_n443), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g490(.A1(new_n689), .A2(new_n488), .ZN(new_n692));
  NAND2_X1  g491(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n693));
  INV_X1    g492(.A(G8gat), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n586), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n692), .A2(new_n693), .A3(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT42), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND4_X1  g497(.A1(new_n692), .A2(KEYINPUT42), .A3(new_n693), .A4(new_n695), .ZN(new_n699));
  OAI211_X1 g498(.A(new_n698), .B(new_n699), .C1(new_n694), .C2(new_n692), .ZN(G1325gat));
  AOI21_X1  g499(.A(G15gat), .B1(new_n689), .B2(new_n308), .ZN(new_n701));
  INV_X1    g500(.A(G15gat), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n310), .A2(new_n702), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n701), .B1(new_n689), .B2(new_n703), .ZN(G1326gat));
  NAND2_X1  g503(.A1(new_n689), .A2(new_n397), .ZN(new_n705));
  XNOR2_X1  g504(.A(KEYINPUT43), .B(G22gat), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n705), .B(new_n706), .ZN(G1327gat));
  INV_X1    g506(.A(new_n688), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n708), .A2(KEYINPUT44), .ZN(new_n709));
  AND3_X1   g508(.A1(new_n514), .A2(new_n522), .A3(KEYINPUT111), .ZN(new_n710));
  AOI21_X1  g509(.A(KEYINPUT111), .B1(new_n514), .B2(new_n522), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n709), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n523), .A2(new_n688), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(KEYINPUT44), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n667), .A2(new_n638), .A3(new_n575), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n715), .A2(new_n443), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(KEYINPUT112), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT112), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n715), .A2(new_n720), .A3(new_n443), .A4(new_n717), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n719), .A2(new_n597), .A3(new_n721), .ZN(new_n722));
  NOR4_X1   g521(.A1(new_n713), .A2(new_n442), .A3(new_n597), .A4(new_n716), .ZN(new_n723));
  XOR2_X1   g522(.A(new_n723), .B(KEYINPUT45), .Z(new_n724));
  NAND2_X1  g523(.A1(new_n722), .A2(new_n724), .ZN(G1328gat));
  NAND3_X1  g524(.A1(new_n715), .A2(new_n488), .A3(new_n717), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT113), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n715), .A2(KEYINPUT113), .A3(new_n488), .A4(new_n717), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n728), .A2(new_n596), .A3(new_n729), .ZN(new_n730));
  NOR4_X1   g529(.A1(new_n713), .A2(new_n596), .A3(new_n503), .A4(new_n716), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(KEYINPUT46), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n730), .A2(new_n732), .ZN(G1329gat));
  INV_X1    g532(.A(KEYINPUT114), .ZN(new_n734));
  AOI211_X1 g533(.A(new_n310), .B(new_n716), .C1(new_n712), .C2(new_n714), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n734), .B1(new_n735), .B2(new_n590), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n708), .B1(new_n514), .B2(new_n522), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n737), .A2(new_n590), .A3(new_n308), .A4(new_n717), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n738), .B1(new_n735), .B2(new_n590), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT47), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n736), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  OAI221_X1 g540(.A(new_n738), .B1(new_n734), .B2(KEYINPUT47), .C1(new_n735), .C2(new_n590), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(G1330gat));
  NOR4_X1   g542(.A1(new_n713), .A2(new_n600), .A3(new_n396), .A4(new_n716), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n715), .A2(new_n397), .A3(new_n717), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n744), .B1(new_n745), .B2(new_n600), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(KEYINPUT48), .ZN(G1331gat));
  OR2_X1    g546(.A1(new_n710), .A2(new_n711), .ZN(new_n748));
  INV_X1    g547(.A(new_n575), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n666), .A2(new_n639), .A3(new_n708), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n748), .A2(new_n749), .A3(new_n751), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n752), .A2(new_n442), .ZN(new_n753));
  XOR2_X1   g552(.A(new_n753), .B(G57gat), .Z(G1332gat));
  AND2_X1   g553(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n755));
  NOR3_X1   g554(.A1(new_n752), .A2(new_n503), .A3(new_n755), .ZN(new_n756));
  NOR2_X1   g555(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n756), .B(new_n757), .ZN(G1333gat));
  INV_X1    g557(.A(new_n308), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n527), .B1(new_n752), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n310), .A2(new_n527), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n748), .A2(new_n749), .A3(new_n751), .A4(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(KEYINPUT50), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT50), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n760), .A2(new_n765), .A3(new_n762), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n764), .A2(new_n766), .ZN(G1334gat));
  NOR2_X1   g566(.A1(new_n752), .A2(new_n396), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(new_n528), .ZN(G1335gat));
  NOR2_X1   g568(.A1(new_n666), .A2(new_n638), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n715), .A2(new_n749), .A3(new_n770), .ZN(new_n771));
  NOR3_X1   g570(.A1(new_n771), .A2(new_n539), .A3(new_n442), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n523), .A2(new_n688), .A3(new_n770), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT51), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n775), .A2(new_n443), .A3(new_n749), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n772), .B1(new_n539), .B2(new_n776), .ZN(G1336gat));
  INV_X1    g576(.A(new_n770), .ZN(new_n778));
  AOI211_X1 g577(.A(new_n575), .B(new_n778), .C1(new_n712), .C2(new_n714), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n540), .B1(new_n779), .B2(new_n488), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n503), .A2(G92gat), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n775), .A2(new_n749), .A3(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(KEYINPUT52), .B1(new_n780), .B2(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(G92gat), .B1(new_n771), .B2(new_n503), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT52), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n785), .A2(new_n786), .A3(new_n782), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n784), .A2(new_n787), .ZN(G1337gat));
  NOR2_X1   g587(.A1(new_n773), .A2(new_n774), .ZN(new_n789));
  AOI21_X1  g588(.A(KEYINPUT51), .B1(new_n737), .B2(new_n770), .ZN(new_n790));
  OAI211_X1 g589(.A(new_n749), .B(new_n308), .C1(new_n789), .C2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(new_n279), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n310), .A2(new_n279), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n715), .A2(new_n749), .A3(new_n770), .A4(new_n793), .ZN(new_n794));
  AND3_X1   g593(.A1(new_n792), .A2(KEYINPUT115), .A3(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(KEYINPUT115), .B1(new_n792), .B2(new_n794), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n795), .A2(new_n796), .ZN(G1338gat));
  NAND4_X1  g596(.A1(new_n715), .A2(new_n749), .A3(new_n397), .A4(new_n770), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(G106gat), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n575), .A2(new_n396), .A3(G106gat), .ZN(new_n800));
  AOI21_X1  g599(.A(KEYINPUT53), .B1(new_n775), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  XOR2_X1   g601(.A(new_n800), .B(KEYINPUT116), .Z(new_n803));
  AOI22_X1  g602(.A1(new_n798), .A2(G106gat), .B1(new_n775), .B2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT53), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n802), .B1(new_n804), .B2(new_n805), .ZN(G1339gat));
  INV_X1    g605(.A(new_n517), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n560), .A2(new_n525), .A3(new_n563), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n572), .A2(KEYINPUT54), .A3(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT54), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n570), .B1(new_n564), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT55), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n809), .A2(KEYINPUT55), .A3(new_n811), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n814), .A2(new_n574), .A3(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT117), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n814), .A2(KEYINPUT117), .A3(new_n574), .A4(new_n815), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n638), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n628), .A2(new_n618), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n821), .B1(new_n621), .B2(new_n624), .ZN(new_n822));
  OR2_X1    g621(.A1(new_n822), .A2(new_n581), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n749), .A2(new_n637), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n688), .B1(new_n820), .B2(new_n824), .ZN(new_n825));
  AND2_X1   g624(.A1(new_n823), .A2(new_n637), .ZN(new_n826));
  AND4_X1   g625(.A1(new_n688), .A2(new_n826), .A3(new_n818), .A4(new_n819), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n667), .B1(new_n825), .B2(new_n827), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n666), .A2(new_n639), .A3(new_n708), .A4(new_n575), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n807), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n488), .A2(new_n442), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(new_n638), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(G113gat), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n834), .B1(new_n240), .B2(new_n833), .ZN(G1340gat));
  NAND2_X1  g634(.A1(new_n832), .A2(new_n749), .ZN(new_n836));
  XNOR2_X1  g635(.A(new_n836), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g636(.A1(new_n832), .A2(new_n666), .ZN(new_n838));
  XNOR2_X1  g637(.A(new_n838), .B(G127gat), .ZN(G1342gat));
  INV_X1    g638(.A(new_n830), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n688), .A2(new_n503), .ZN(new_n841));
  XNOR2_X1  g640(.A(new_n841), .B(KEYINPUT118), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(new_n443), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n840), .A2(G134gat), .A3(new_n843), .ZN(new_n844));
  XNOR2_X1  g643(.A(KEYINPUT119), .B(KEYINPUT56), .ZN(new_n845));
  XNOR2_X1  g644(.A(new_n844), .B(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(new_n832), .ZN(new_n847));
  OAI21_X1  g646(.A(G134gat), .B1(new_n847), .B2(new_n708), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n846), .A2(new_n848), .ZN(G1343gat));
  AOI21_X1  g648(.A(new_n396), .B1(new_n828), .B2(new_n829), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n310), .A2(new_n831), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n638), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(new_n331), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT58), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(KEYINPUT121), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n828), .A2(new_n829), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n396), .A2(KEYINPUT57), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n824), .B1(new_n639), .B2(new_n816), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT120), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  OAI211_X1 g661(.A(KEYINPUT120), .B(new_n824), .C1(new_n639), .C2(new_n816), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n688), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n667), .B1(new_n864), .B2(new_n827), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n396), .B1(new_n865), .B2(new_n829), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT57), .ZN(new_n867));
  OAI211_X1 g666(.A(new_n851), .B(new_n859), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n638), .A2(G141gat), .ZN(new_n869));
  OAI211_X1 g668(.A(new_n854), .B(new_n856), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  OR2_X1    g669(.A1(new_n855), .A2(KEYINPUT121), .ZN(new_n871));
  XNOR2_X1  g670(.A(new_n870), .B(new_n871), .ZN(G1344gat));
  INV_X1    g671(.A(KEYINPUT59), .ZN(new_n873));
  AOI211_X1 g672(.A(new_n873), .B(G148gat), .C1(new_n852), .C2(new_n749), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n873), .B1(new_n868), .B2(new_n575), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n862), .A2(new_n863), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(new_n708), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n688), .A2(new_n826), .ZN(new_n878));
  OR2_X1    g677(.A1(new_n878), .A2(new_n816), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n666), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(new_n829), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n858), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  OR2_X1    g681(.A1(new_n850), .A2(new_n867), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(new_n749), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n851), .A2(KEYINPUT59), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n875), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n874), .B1(new_n887), .B2(G148gat), .ZN(G1345gat));
  NOR3_X1   g687(.A1(new_n868), .A2(new_n334), .A3(new_n667), .ZN(new_n889));
  AOI21_X1  g688(.A(G155gat), .B1(new_n852), .B2(new_n666), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n889), .A2(new_n890), .ZN(G1346gat));
  OAI21_X1  g690(.A(G162gat), .B1(new_n868), .B2(new_n708), .ZN(new_n892));
  INV_X1    g691(.A(new_n843), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n893), .A2(new_n850), .A3(new_n335), .A4(new_n310), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n892), .A2(new_n894), .ZN(G1347gat));
  NOR2_X1   g694(.A1(new_n503), .A2(new_n443), .ZN(new_n896));
  AND3_X1   g695(.A1(new_n857), .A2(new_n517), .A3(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(G169gat), .B1(new_n898), .B2(new_n639), .ZN(new_n899));
  AOI21_X1  g698(.A(KEYINPUT122), .B1(new_n857), .B2(new_n442), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT122), .ZN(new_n901));
  AOI211_X1 g700(.A(new_n901), .B(new_n443), .C1(new_n828), .C2(new_n829), .ZN(new_n902));
  OAI211_X1 g701(.A(new_n488), .B(new_n517), .C1(new_n900), .C2(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n638), .A2(new_n226), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n899), .B1(new_n903), .B2(new_n904), .ZN(G1348gat));
  OAI21_X1  g704(.A(new_n227), .B1(new_n903), .B2(new_n575), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n897), .A2(new_n749), .A3(new_n267), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT123), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n906), .A2(KEYINPUT123), .A3(new_n907), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(G1349gat));
  INV_X1    g711(.A(KEYINPUT125), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT60), .ZN(new_n914));
  INV_X1    g713(.A(new_n220), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n903), .A2(new_n667), .A3(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT124), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n897), .A2(new_n917), .A3(new_n666), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n830), .A2(new_n666), .A3(new_n896), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(KEYINPUT124), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n255), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  OAI211_X1 g720(.A(new_n913), .B(new_n914), .C1(new_n916), .C2(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(new_n900), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n857), .A2(KEYINPUT122), .A3(new_n442), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n807), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND4_X1  g724(.A1(new_n925), .A2(new_n666), .A3(new_n220), .A4(new_n488), .ZN(new_n926));
  INV_X1    g725(.A(new_n920), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n919), .A2(KEYINPUT124), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n217), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(new_n930));
  NAND2_X1  g729(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n931));
  NAND4_X1  g730(.A1(new_n926), .A2(new_n929), .A3(new_n930), .A4(new_n931), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n922), .A2(new_n932), .ZN(G1350gat));
  AOI21_X1  g732(.A(new_n221), .B1(new_n897), .B2(new_n688), .ZN(new_n934));
  XOR2_X1   g733(.A(new_n934), .B(KEYINPUT61), .Z(new_n935));
  NOR3_X1   g734(.A1(new_n903), .A2(G190gat), .A3(new_n708), .ZN(new_n936));
  AND2_X1   g735(.A1(new_n936), .A2(KEYINPUT126), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n936), .A2(KEYINPUT126), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n935), .B1(new_n937), .B2(new_n938), .ZN(G1351gat));
  AND2_X1   g738(.A1(new_n310), .A2(new_n488), .ZN(new_n940));
  OAI211_X1 g739(.A(new_n397), .B(new_n940), .C1(new_n900), .C2(new_n902), .ZN(new_n941));
  INV_X1    g740(.A(new_n941), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n942), .A2(new_n578), .A3(new_n638), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n310), .A2(new_n896), .ZN(new_n944));
  INV_X1    g743(.A(new_n944), .ZN(new_n945));
  NAND4_X1  g744(.A1(new_n882), .A2(new_n638), .A3(new_n883), .A4(new_n945), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(G197gat), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n943), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(KEYINPUT127), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT127), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n943), .A2(new_n950), .A3(new_n947), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n949), .A2(new_n951), .ZN(G1352gat));
  NOR3_X1   g751(.A1(new_n941), .A2(G204gat), .A3(new_n575), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT62), .ZN(new_n954));
  OR2_X1    g753(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g754(.A(G204gat), .B1(new_n885), .B2(new_n944), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n953), .A2(new_n954), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n955), .A2(new_n956), .A3(new_n957), .ZN(G1353gat));
  OR3_X1    g757(.A1(new_n941), .A2(G211gat), .A3(new_n667), .ZN(new_n959));
  NAND4_X1  g758(.A1(new_n882), .A2(new_n666), .A3(new_n883), .A4(new_n945), .ZN(new_n960));
  AND3_X1   g759(.A1(new_n960), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n961));
  AOI21_X1  g760(.A(KEYINPUT63), .B1(new_n960), .B2(G211gat), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n959), .B1(new_n961), .B2(new_n962), .ZN(G1354gat));
  NAND4_X1  g762(.A1(new_n884), .A2(new_n688), .A3(new_n323), .A4(new_n945), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n313), .B1(new_n941), .B2(new_n708), .ZN(new_n965));
  AND2_X1   g764(.A1(new_n964), .A2(new_n965), .ZN(G1355gat));
endmodule


