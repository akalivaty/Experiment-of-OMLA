//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 1 1 0 1 0 1 1 1 1 0 0 0 1 0 0 0 1 1 0 0 1 0 0 0 0 1 0 1 1 1 1 0 0 0 0 0 1 1 1 1 1 0 0 0 0 1 0 0 0 0 0 1 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:04 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1303, new_n1304, new_n1305, new_n1306, new_n1307, new_n1308,
    new_n1310, new_n1311, new_n1312, new_n1313, new_n1314, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1367, new_n1368, new_n1369, new_n1370, new_n1371,
    new_n1372, new_n1373, new_n1374;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n207));
  XOR2_X1   g0007(.A(new_n207), .B(KEYINPUT64), .Z(new_n208));
  AOI22_X1  g0008(.A1(G58), .A2(G232), .B1(G116), .B2(G270), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n211));
  NAND3_X1  g0011(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  OAI21_X1  g0012(.A(new_n206), .B1(new_n208), .B2(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(KEYINPUT1), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT65), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n206), .A2(G13), .ZN(new_n216));
  OAI211_X1 g0016(.A(new_n216), .B(G250), .C1(G257), .C2(G264), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT0), .ZN(new_n218));
  OAI21_X1  g0018(.A(G50), .B1(G58), .B2(G68), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G13), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n221), .A2(new_n204), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n218), .B(new_n223), .C1(KEYINPUT1), .C2(new_n213), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n215), .A2(new_n224), .ZN(G361));
  XOR2_X1   g0025(.A(G238), .B(G244), .Z(new_n226));
  XNOR2_X1  g0026(.A(G226), .B(G232), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT67), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G264), .B(G270), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n231), .B(new_n234), .ZN(G358));
  XNOR2_X1  g0035(.A(G68), .B(G77), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT68), .ZN(new_n237));
  XOR2_X1   g0037(.A(G50), .B(G58), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XOR2_X1   g0040(.A(G107), .B(G116), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  XNOR2_X1  g0043(.A(KEYINPUT3), .B(G33), .ZN(new_n244));
  NOR2_X1   g0044(.A1(G232), .A2(G1698), .ZN(new_n245));
  INV_X1    g0045(.A(G1698), .ZN(new_n246));
  NOR2_X1   g0046(.A1(new_n246), .A2(G238), .ZN(new_n247));
  OAI21_X1  g0047(.A(new_n244), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  AOI21_X1  g0048(.A(new_n221), .B1(G33), .B2(G41), .ZN(new_n249));
  OAI211_X1 g0049(.A(new_n248), .B(new_n249), .C1(G107), .C2(new_n244), .ZN(new_n250));
  OR2_X1    g0050(.A1(KEYINPUT69), .A2(G45), .ZN(new_n251));
  INV_X1    g0051(.A(G41), .ZN(new_n252));
  NAND2_X1  g0052(.A1(KEYINPUT69), .A2(G45), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n251), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n203), .A2(G274), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G45), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n252), .A2(new_n258), .ZN(new_n259));
  AND2_X1   g0059(.A1(G1), .A2(G13), .ZN(new_n260));
  NAND2_X1  g0060(.A1(G33), .A2(G41), .ZN(new_n261));
  AOI22_X1  g0061(.A1(new_n203), .A2(new_n259), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G244), .ZN(new_n263));
  AND3_X1   g0063(.A1(new_n250), .A2(new_n257), .A3(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G179), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g0066(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(new_n221), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT72), .ZN(new_n269));
  INV_X1    g0069(.A(G33), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n269), .B1(new_n270), .B2(G20), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n204), .A2(KEYINPUT72), .A3(G33), .ZN(new_n272));
  AND2_X1   g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  XNOR2_X1  g0073(.A(KEYINPUT15), .B(G87), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g0075(.A(KEYINPUT8), .B(G58), .ZN(new_n276));
  NOR2_X1   g0076(.A1(G20), .A2(G33), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G77), .ZN(new_n279));
  OAI22_X1  g0079(.A1(new_n276), .A2(new_n278), .B1(new_n204), .B2(new_n279), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n268), .B1(new_n275), .B2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G13), .ZN(new_n282));
  NOR3_X1   g0082(.A1(new_n282), .A2(new_n204), .A3(G1), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n283), .A2(new_n268), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n279), .B1(new_n203), .B2(G20), .ZN(new_n285));
  AOI22_X1  g0085(.A1(new_n284), .A2(new_n285), .B1(new_n279), .B2(new_n283), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n281), .A2(new_n286), .ZN(new_n287));
  OAI211_X1 g0087(.A(new_n266), .B(new_n287), .C1(G169), .C2(new_n264), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n287), .B1(G190), .B2(new_n264), .ZN(new_n289));
  INV_X1    g0089(.A(G200), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n289), .B1(new_n290), .B2(new_n264), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n262), .A2(G226), .B1(new_n254), .B2(new_n256), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n244), .A2(G223), .A3(G1698), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n293), .B1(new_n279), .B2(new_n244), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n244), .A2(G222), .A3(new_n246), .ZN(new_n295));
  OR2_X1    g0095(.A1(new_n295), .A2(KEYINPUT70), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(KEYINPUT70), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n294), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n261), .A2(G1), .A3(G13), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n292), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G169), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  AND3_X1   g0102(.A1(new_n267), .A2(KEYINPUT71), .A3(new_n221), .ZN(new_n303));
  AOI21_X1  g0103(.A(KEYINPUT71), .B1(new_n267), .B2(new_n221), .ZN(new_n304));
  NOR3_X1   g0104(.A1(new_n303), .A2(new_n304), .A3(new_n283), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n305), .B(G50), .C1(G1), .C2(new_n204), .ZN(new_n306));
  INV_X1    g0106(.A(G50), .ZN(new_n307));
  INV_X1    g0107(.A(G58), .ZN(new_n308));
  INV_X1    g0108(.A(G68), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  AOI22_X1  g0110(.A1(new_n310), .A2(G20), .B1(G150), .B2(new_n277), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n311), .B1(new_n273), .B2(new_n276), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT71), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n268), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n267), .A2(KEYINPUT71), .A3(new_n221), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n312), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n283), .A2(new_n307), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n306), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  OAI211_X1 g0119(.A(new_n292), .B(new_n265), .C1(new_n298), .C2(new_n299), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n302), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT73), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n319), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n324), .B1(new_n300), .B2(new_n301), .ZN(new_n325));
  AOI21_X1  g0125(.A(KEYINPUT73), .B1(new_n325), .B2(new_n320), .ZN(new_n326));
  OAI211_X1 g0126(.A(new_n288), .B(new_n291), .C1(new_n323), .C2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT9), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n319), .A2(new_n328), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n306), .A2(new_n317), .A3(KEYINPUT9), .A4(new_n318), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT74), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(KEYINPUT10), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n329), .A2(new_n330), .A3(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n331), .A2(KEYINPUT10), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n300), .A2(G200), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n292), .B(G190), .C1(new_n298), .C2(new_n299), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n334), .A2(new_n336), .A3(new_n337), .A4(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n337), .A2(new_n338), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n335), .B1(new_n340), .B2(new_n333), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  OAI21_X1  g0142(.A(KEYINPUT75), .B1(new_n327), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n291), .A2(new_n288), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n321), .A2(new_n322), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n325), .A2(KEYINPUT73), .A3(new_n320), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n344), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT75), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n347), .A2(new_n348), .A3(new_n341), .A4(new_n339), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT16), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT7), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n351), .B1(new_n244), .B2(G20), .ZN(new_n352));
  AND2_X1   g0152(.A1(KEYINPUT3), .A2(G33), .ZN(new_n353));
  NOR2_X1   g0153(.A1(KEYINPUT3), .A2(G33), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n355), .A2(KEYINPUT7), .A3(new_n204), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n309), .B1(new_n352), .B2(new_n356), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n308), .A2(new_n309), .ZN(new_n358));
  NOR2_X1   g0158(.A1(G58), .A2(G68), .ZN(new_n359));
  OAI21_X1  g0159(.A(G20), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n277), .A2(G159), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n350), .B1(new_n357), .B2(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(KEYINPUT7), .B1(new_n355), .B2(new_n204), .ZN(new_n364));
  NOR4_X1   g0164(.A1(new_n353), .A2(new_n354), .A3(new_n351), .A4(G20), .ZN(new_n365));
  OAI21_X1  g0165(.A(G68), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n362), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n366), .A2(KEYINPUT16), .A3(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n363), .A2(new_n368), .A3(new_n268), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n276), .B1(new_n203), .B2(G20), .ZN(new_n370));
  AOI22_X1  g0170(.A1(new_n305), .A2(new_n370), .B1(new_n283), .B2(new_n276), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(G223), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(new_n246), .ZN(new_n374));
  INV_X1    g0174(.A(G226), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(G1698), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n374), .B(new_n376), .C1(new_n353), .C2(new_n354), .ZN(new_n377));
  NAND2_X1  g0177(.A1(G33), .A2(G87), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n299), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n299), .A2(G232), .A3(new_n380), .ZN(new_n381));
  AND2_X1   g0181(.A1(KEYINPUT69), .A2(G45), .ZN(new_n382));
  NOR2_X1   g0182(.A1(KEYINPUT69), .A2(G45), .ZN(new_n383));
  NOR3_X1   g0183(.A1(new_n382), .A2(new_n383), .A3(G41), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n381), .B1(new_n384), .B2(new_n255), .ZN(new_n385));
  NOR3_X1   g0185(.A1(new_n379), .A2(new_n385), .A3(G179), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n377), .A2(new_n378), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n249), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT76), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n262), .A2(G232), .B1(new_n254), .B2(new_n256), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  OAI21_X1  g0191(.A(KEYINPUT76), .B1(new_n379), .B2(new_n385), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n386), .B1(new_n393), .B2(new_n301), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n372), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(KEYINPUT18), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT18), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n372), .A2(new_n394), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT77), .ZN(new_n400));
  AOI21_X1  g0200(.A(G200), .B1(new_n391), .B2(new_n392), .ZN(new_n401));
  NOR3_X1   g0201(.A1(new_n379), .A2(new_n385), .A3(G190), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n369), .B(new_n371), .C1(new_n401), .C2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT17), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n371), .ZN(new_n406));
  INV_X1    g0206(.A(new_n268), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n366), .A2(new_n367), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n407), .B1(new_n408), .B2(new_n350), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n406), .B1(new_n409), .B2(new_n368), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n389), .B1(new_n388), .B2(new_n390), .ZN(new_n411));
  NOR3_X1   g0211(.A1(new_n379), .A2(new_n385), .A3(KEYINPUT76), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n290), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n402), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(KEYINPUT17), .B1(new_n410), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n400), .B1(new_n405), .B2(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n410), .A2(new_n415), .A3(KEYINPUT17), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n402), .B1(new_n393), .B2(new_n290), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n404), .B1(new_n372), .B2(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n418), .A2(new_n420), .A3(KEYINPUT77), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n399), .B1(new_n417), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n375), .A2(new_n246), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n244), .B(new_n423), .C1(G232), .C2(new_n246), .ZN(new_n424));
  NAND2_X1  g0224(.A1(G33), .A2(G97), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n299), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n262), .A2(G238), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(new_n257), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT13), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OAI21_X1  g0231(.A(KEYINPUT13), .B1(new_n426), .B2(new_n428), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(G190), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n273), .A2(new_n279), .ZN(new_n436));
  OAI22_X1  g0236(.A1(new_n278), .A2(new_n307), .B1(new_n204), .B2(G68), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n316), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT11), .ZN(new_n439));
  OR2_X1    g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n438), .A2(new_n439), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n282), .A2(G1), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(G20), .ZN(new_n443));
  OR3_X1    g0243(.A1(new_n443), .A2(KEYINPUT12), .A3(G68), .ZN(new_n444));
  OAI21_X1  g0244(.A(KEYINPUT12), .B1(new_n443), .B2(G68), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n309), .B1(new_n203), .B2(G20), .ZN(new_n446));
  AOI22_X1  g0246(.A1(new_n444), .A2(new_n445), .B1(new_n284), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n440), .A2(new_n441), .A3(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n290), .B1(new_n431), .B2(new_n432), .ZN(new_n449));
  NOR3_X1   g0249(.A1(new_n435), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n432), .ZN(new_n451));
  NOR3_X1   g0251(.A1(new_n426), .A2(new_n428), .A3(KEYINPUT13), .ZN(new_n452));
  OAI21_X1  g0252(.A(G169), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(KEYINPUT14), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT14), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n455), .B(G169), .C1(new_n451), .C2(new_n452), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n454), .B(new_n456), .C1(new_n265), .C2(new_n433), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n450), .B1(new_n457), .B2(new_n448), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n343), .A2(new_n349), .A3(new_n422), .A4(new_n458), .ZN(new_n459));
  OAI211_X1 g0259(.A(G257), .B(G1698), .C1(new_n353), .C2(new_n354), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT85), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n244), .A2(KEYINPUT85), .A3(G257), .A4(G1698), .ZN(new_n463));
  NAND2_X1  g0263(.A1(G33), .A2(G294), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n244), .A2(G250), .A3(new_n246), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n462), .A2(new_n463), .A3(new_n464), .A4(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n249), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n203), .A2(G45), .ZN(new_n468));
  NOR2_X1   g0268(.A1(KEYINPUT5), .A2(G41), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(KEYINPUT5), .A2(G41), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n468), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(G274), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n258), .A2(G1), .ZN(new_n474));
  INV_X1    g0274(.A(new_n471), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n474), .B1(new_n475), .B2(new_n469), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n476), .A2(G264), .A3(new_n299), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n473), .A2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n467), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(new_n301), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n478), .B1(new_n466), .B2(new_n249), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n265), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n204), .B(G87), .C1(new_n353), .C2(new_n354), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(KEYINPUT22), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT22), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n244), .A2(new_n486), .A3(new_n204), .A4(G87), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(G116), .ZN(new_n489));
  NOR3_X1   g0289(.A1(new_n270), .A2(new_n489), .A3(G20), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT23), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n491), .B1(new_n204), .B2(G107), .ZN(new_n492));
  INV_X1    g0292(.A(G107), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n493), .A2(KEYINPUT23), .A3(G20), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n490), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n488), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(KEYINPUT24), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT24), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n488), .A2(new_n498), .A3(new_n495), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n407), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n283), .A2(new_n493), .ZN(new_n501));
  XNOR2_X1  g0301(.A(new_n501), .B(KEYINPUT25), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n203), .A2(G33), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n314), .A2(new_n443), .A3(new_n315), .A4(new_n503), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n504), .A2(new_n493), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n481), .B(new_n483), .C1(new_n500), .C2(new_n507), .ZN(new_n508));
  AND3_X1   g0308(.A1(new_n482), .A2(KEYINPUT86), .A3(new_n434), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n482), .A2(new_n434), .ZN(new_n510));
  OAI21_X1  g0310(.A(KEYINPUT86), .B1(new_n482), .B2(G200), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(new_n499), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n498), .B1(new_n488), .B2(new_n495), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n268), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(new_n506), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n508), .B1(new_n512), .B2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(G97), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n283), .A2(new_n518), .ZN(new_n519));
  XNOR2_X1  g0319(.A(new_n519), .B(KEYINPUT78), .ZN(new_n520));
  OAI21_X1  g0320(.A(G107), .B1(new_n364), .B2(new_n365), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT6), .ZN(new_n522));
  AND2_X1   g0322(.A1(G97), .A2(G107), .ZN(new_n523));
  NOR2_X1   g0323(.A1(G97), .A2(G107), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n493), .A2(KEYINPUT6), .A3(G97), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  AOI22_X1  g0327(.A1(new_n527), .A2(G20), .B1(G77), .B2(new_n277), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n521), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n520), .B1(new_n529), .B2(new_n268), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n305), .A2(G97), .A3(new_n503), .ZN(new_n531));
  OAI211_X1 g0331(.A(G244), .B(new_n246), .C1(new_n353), .C2(new_n354), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT4), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(G33), .A2(G283), .ZN(new_n535));
  INV_X1    g0335(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(G250), .A2(G1698), .ZN(new_n537));
  NAND2_X1  g0337(.A1(KEYINPUT4), .A2(G244), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n537), .B1(new_n538), .B2(G1698), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n536), .B1(new_n244), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n534), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(new_n249), .ZN(new_n542));
  XNOR2_X1  g0342(.A(KEYINPUT5), .B(G41), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n543), .A2(new_n474), .B1(new_n260), .B2(new_n261), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n544), .A2(G257), .B1(G274), .B2(new_n472), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  AOI22_X1  g0346(.A1(new_n530), .A2(new_n531), .B1(new_n301), .B2(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(KEYINPUT79), .B1(new_n541), .B2(new_n249), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT79), .ZN(new_n549));
  AOI211_X1 g0349(.A(new_n549), .B(new_n299), .C1(new_n534), .C2(new_n540), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n265), .B(new_n545), .C1(new_n548), .C2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n542), .A2(G190), .A3(new_n545), .ZN(new_n552));
  AND3_X1   g0352(.A1(new_n493), .A2(KEYINPUT6), .A3(G97), .ZN(new_n553));
  XNOR2_X1  g0353(.A(G97), .B(G107), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n553), .B1(new_n554), .B2(new_n522), .ZN(new_n555));
  OAI22_X1  g0355(.A1(new_n555), .A2(new_n204), .B1(new_n279), .B2(new_n278), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n493), .B1(new_n352), .B2(new_n356), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n268), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(new_n520), .ZN(new_n559));
  AND4_X1   g0359(.A1(new_n552), .A2(new_n558), .A3(new_n531), .A4(new_n559), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n545), .B1(new_n548), .B2(new_n550), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(G200), .ZN(new_n562));
  AOI22_X1  g0362(.A1(new_n547), .A2(new_n551), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  OAI211_X1 g0363(.A(G257), .B(new_n246), .C1(new_n353), .C2(new_n354), .ZN(new_n564));
  OAI211_X1 g0364(.A(G264), .B(G1698), .C1(new_n353), .C2(new_n354), .ZN(new_n565));
  XNOR2_X1  g0365(.A(KEYINPUT83), .B(G303), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n564), .B(new_n565), .C1(new_n244), .C2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n249), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n544), .A2(G270), .B1(G274), .B2(new_n472), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(G200), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n489), .B1(new_n203), .B2(G33), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n204), .A2(G116), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n284), .A2(new_n572), .B1(new_n442), .B2(new_n573), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n535), .B(new_n204), .C1(G33), .C2(new_n518), .ZN(new_n575));
  INV_X1    g0375(.A(new_n573), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n575), .A2(new_n576), .A3(new_n268), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT20), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n573), .B1(new_n221), .B2(new_n267), .ZN(new_n580));
  AOI21_X1  g0380(.A(KEYINPUT20), .B1(new_n580), .B2(new_n575), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n574), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n568), .A2(new_n569), .A3(G190), .ZN(new_n584));
  AND3_X1   g0384(.A1(new_n571), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT84), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT21), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n570), .A2(new_n582), .A3(G169), .A4(new_n588), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n582), .A2(G179), .A3(new_n568), .A4(new_n569), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n301), .B1(new_n568), .B2(new_n569), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n588), .B1(new_n592), .B2(new_n582), .ZN(new_n593));
  NOR3_X1   g0393(.A1(new_n585), .A2(new_n591), .A3(new_n593), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n305), .A2(KEYINPUT82), .A3(G87), .A4(new_n503), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT82), .ZN(new_n596));
  INV_X1    g0396(.A(G87), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n596), .B1(new_n504), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n274), .A2(new_n283), .ZN(new_n600));
  NAND3_X1  g0400(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n601));
  AND2_X1   g0401(.A1(new_n601), .A2(new_n204), .ZN(new_n602));
  NOR3_X1   g0402(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n603));
  OAI21_X1  g0403(.A(KEYINPUT80), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  AOI22_X1  g0404(.A1(new_n204), .A2(new_n601), .B1(new_n524), .B2(new_n597), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT80), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n244), .A2(new_n204), .A3(G68), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n518), .B1(new_n271), .B2(new_n272), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n609), .B1(new_n610), .B2(KEYINPUT19), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n268), .B1(new_n608), .B2(new_n611), .ZN(new_n612));
  AND3_X1   g0412(.A1(new_n599), .A2(new_n600), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n468), .A2(G250), .ZN(new_n614));
  OAI22_X1  g0414(.A1(new_n249), .A2(new_n614), .B1(new_n258), .B2(new_n255), .ZN(new_n615));
  OAI211_X1 g0415(.A(G244), .B(G1698), .C1(new_n353), .C2(new_n354), .ZN(new_n616));
  OAI211_X1 g0416(.A(G238), .B(new_n246), .C1(new_n353), .C2(new_n354), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n616), .B(new_n617), .C1(new_n270), .C2(new_n489), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n615), .B1(new_n618), .B2(new_n249), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n434), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n620), .B1(G200), .B2(new_n619), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n613), .A2(new_n621), .ZN(new_n622));
  OR2_X1    g0422(.A1(new_n504), .A2(new_n274), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n612), .A2(new_n600), .A3(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT81), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n612), .A2(KEYINPUT81), .A3(new_n600), .A4(new_n623), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n618), .A2(new_n249), .ZN(new_n628));
  INV_X1    g0428(.A(new_n615), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n628), .A2(new_n629), .A3(G179), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n630), .B1(new_n301), .B2(new_n619), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n626), .A2(new_n627), .A3(new_n631), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n563), .A2(new_n594), .A3(new_n622), .A4(new_n632), .ZN(new_n633));
  NOR3_X1   g0433(.A1(new_n459), .A2(new_n517), .A3(new_n633), .ZN(G372));
  OAI21_X1  g0434(.A(new_n456), .B1(new_n265), .B2(new_n433), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n455), .B1(new_n433), .B2(G169), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n448), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n637), .B1(new_n450), .B2(new_n288), .ZN(new_n638));
  AOI21_X1  g0438(.A(KEYINPUT77), .B1(new_n418), .B2(new_n420), .ZN(new_n639));
  AND3_X1   g0439(.A1(new_n418), .A2(new_n420), .A3(KEYINPUT77), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n638), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n396), .A2(new_n398), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n342), .ZN(new_n644));
  AOI22_X1  g0444(.A1(new_n643), .A2(new_n644), .B1(new_n345), .B2(new_n346), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n631), .A2(new_n624), .ZN(new_n646));
  INV_X1    g0446(.A(new_n509), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n511), .A2(new_n510), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n500), .A2(new_n507), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n591), .A2(new_n593), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n508), .ZN(new_n653));
  AOI22_X1  g0453(.A1(new_n613), .A2(new_n621), .B1(new_n624), .B2(new_n631), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n651), .A2(new_n653), .A3(new_n563), .A4(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n558), .A2(new_n531), .A3(new_n559), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n546), .A2(new_n301), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n551), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT87), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n551), .A2(new_n656), .A3(KEYINPUT87), .A4(new_n657), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n660), .A2(new_n654), .A3(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT26), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  AND3_X1   g0464(.A1(new_n551), .A2(new_n656), .A3(new_n657), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n665), .A2(new_n632), .A3(new_n622), .ZN(new_n666));
  XNOR2_X1  g0466(.A(KEYINPUT88), .B(KEYINPUT26), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  OAI211_X1 g0468(.A(new_n646), .B(new_n655), .C1(new_n664), .C2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n645), .B1(new_n459), .B2(new_n670), .ZN(G369));
  NAND2_X1  g0471(.A1(new_n442), .A2(new_n204), .ZN(new_n672));
  OR2_X1    g0472(.A1(new_n672), .A2(KEYINPUT27), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(KEYINPUT27), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(G213), .A3(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(G343), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n508), .A2(new_n677), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n516), .B1(new_n647), .B2(new_n648), .ZN(new_n679));
  INV_X1    g0479(.A(new_n508), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT89), .ZN(new_n682));
  INV_X1    g0482(.A(new_n677), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n516), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n681), .A2(new_n682), .A3(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n650), .A2(new_n677), .ZN(new_n686));
  OAI21_X1  g0486(.A(KEYINPUT89), .B1(new_n517), .B2(new_n686), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n678), .B1(new_n685), .B2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n677), .A2(new_n583), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n690), .B1(new_n591), .B2(new_n593), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n571), .A2(new_n583), .A3(new_n584), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n652), .A2(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n691), .B1(new_n693), .B2(new_n690), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(G330), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n689), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n680), .A2(new_n677), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n652), .A2(new_n683), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n685), .A2(new_n687), .A3(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n697), .A2(new_n698), .A3(new_n700), .ZN(G399));
  NAND3_X1  g0501(.A1(new_n216), .A2(KEYINPUT90), .A3(new_n252), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(KEYINPUT90), .B1(new_n216), .B2(new_n252), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n603), .A2(new_n489), .ZN(new_n706));
  NOR3_X1   g0506(.A1(new_n705), .A2(new_n203), .A3(new_n706), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n707), .B1(new_n220), .B2(new_n705), .ZN(new_n708));
  XOR2_X1   g0508(.A(new_n708), .B(KEYINPUT28), .Z(new_n709));
  INV_X1    g0509(.A(KEYINPUT29), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n655), .A2(new_n646), .ZN(new_n711));
  INV_X1    g0511(.A(new_n666), .ZN(new_n712));
  INV_X1    g0512(.A(new_n667), .ZN(new_n713));
  AOI22_X1  g0513(.A1(new_n712), .A2(new_n713), .B1(new_n662), .B2(new_n663), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n677), .B1(new_n711), .B2(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n710), .B1(new_n715), .B2(KEYINPUT93), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n666), .A2(new_n667), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n660), .A2(new_n654), .A3(KEYINPUT26), .A4(new_n661), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT94), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n717), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  AND2_X1   g0520(.A1(new_n718), .A2(new_n719), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n677), .B1(new_n722), .B2(new_n711), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT93), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n715), .A2(new_n724), .ZN(new_n725));
  AOI22_X1  g0525(.A1(new_n716), .A2(new_n723), .B1(new_n725), .B2(new_n710), .ZN(new_n726));
  INV_X1    g0526(.A(G330), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n560), .A2(new_n562), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n728), .A2(new_n632), .A3(new_n658), .A4(new_n622), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n730), .A2(new_n681), .A3(new_n594), .A4(new_n677), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT92), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n729), .A2(new_n693), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n734), .A2(KEYINPUT92), .A3(new_n681), .A4(new_n677), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  AND2_X1   g0536(.A1(new_n467), .A2(new_n619), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n570), .A2(new_n265), .ZN(new_n738));
  AND3_X1   g0538(.A1(new_n542), .A2(new_n477), .A3(new_n545), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n737), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT30), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n619), .A2(G179), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n561), .A2(new_n480), .A3(new_n570), .A4(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n740), .A2(new_n741), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n683), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  OR2_X1    g0547(.A1(KEYINPUT91), .A2(KEYINPUT31), .ZN(new_n748));
  NAND2_X1  g0548(.A1(KEYINPUT91), .A2(KEYINPUT31), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n747), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n750), .B1(new_n748), .B2(new_n747), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n727), .B1(new_n736), .B2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n726), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n709), .B1(new_n755), .B2(G1), .ZN(G364));
  NOR2_X1   g0556(.A1(new_n282), .A2(G20), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n203), .B1(new_n757), .B2(G45), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n705), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n216), .A2(new_n244), .ZN(new_n761));
  INV_X1    g0561(.A(G355), .ZN(new_n762));
  OAI22_X1  g0562(.A1(new_n761), .A2(new_n762), .B1(G116), .B2(new_n216), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n239), .A2(G45), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n216), .A2(new_n355), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n382), .A2(new_n383), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n765), .B1(new_n220), .B2(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n763), .B1(new_n764), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(G13), .A2(G33), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(G20), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n221), .B1(G20), .B2(new_n301), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n760), .B1(new_n768), .B2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n204), .A2(G190), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n776), .A2(new_n265), .A3(G200), .ZN(new_n777));
  INV_X1    g0577(.A(G283), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n204), .A2(new_n434), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n780), .A2(new_n265), .A3(G200), .ZN(new_n781));
  INV_X1    g0581(.A(G303), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n265), .A2(G200), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(new_n776), .ZN(new_n784));
  INV_X1    g0584(.A(G311), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n781), .A2(new_n782), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(G179), .A2(G200), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n776), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  AOI211_X1 g0589(.A(new_n779), .B(new_n786), .C1(G329), .C2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n204), .A2(new_n265), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n791), .A2(G190), .A3(G200), .ZN(new_n792));
  AND2_X1   g0592(.A1(new_n792), .A2(KEYINPUT95), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n792), .A2(KEYINPUT95), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(G326), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n791), .A2(new_n434), .A3(G200), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(G317), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(KEYINPUT33), .ZN(new_n801));
  OR2_X1    g0601(.A1(new_n800), .A2(KEYINPUT33), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n799), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n780), .A2(new_n783), .ZN(new_n804));
  INV_X1    g0604(.A(G322), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n355), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n204), .B1(new_n787), .B2(G190), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n806), .B1(G294), .B2(new_n808), .ZN(new_n809));
  NAND4_X1  g0609(.A1(new_n790), .A2(new_n797), .A3(new_n803), .A4(new_n809), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n804), .A2(new_n308), .B1(new_n784), .B2(new_n279), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n811), .B1(new_n796), .B2(G50), .ZN(new_n812));
  XOR2_X1   g0612(.A(new_n812), .B(KEYINPUT96), .Z(new_n813));
  NAND2_X1  g0613(.A1(new_n789), .A2(G159), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n814), .B(KEYINPUT32), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n244), .B1(new_n777), .B2(new_n493), .C1(new_n597), .C2(new_n781), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n798), .A2(new_n309), .B1(new_n807), .B2(new_n518), .ZN(new_n817));
  OR3_X1    g0617(.A1(new_n815), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n810), .B1(new_n813), .B2(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n775), .B1(new_n819), .B2(new_n772), .ZN(new_n820));
  INV_X1    g0620(.A(new_n771), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n820), .B1(new_n694), .B2(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n694), .A2(G330), .ZN(new_n823));
  INV_X1    g0623(.A(new_n760), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n695), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n822), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n826), .B(KEYINPUT97), .ZN(G396));
  NOR2_X1   g0627(.A1(new_n344), .A2(new_n683), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n828), .B1(new_n711), .B2(new_n714), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n683), .A2(new_n287), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n291), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(new_n288), .ZN(new_n833));
  OR2_X1    g0633(.A1(new_n288), .A2(new_n683), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n830), .B1(new_n715), .B2(new_n835), .ZN(new_n836));
  OR2_X1    g0636(.A1(new_n836), .A2(new_n752), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(new_n752), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n837), .A2(new_n824), .A3(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n772), .A2(new_n769), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n824), .B1(new_n279), .B2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n772), .ZN(new_n842));
  INV_X1    g0642(.A(new_n804), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n244), .B1(new_n843), .B2(G294), .ZN(new_n844));
  OAI221_X1 g0644(.A(new_n844), .B1(new_n518), .B2(new_n807), .C1(new_n778), .C2(new_n798), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n795), .A2(new_n782), .ZN(new_n846));
  OAI22_X1  g0646(.A1(new_n777), .A2(new_n597), .B1(new_n788), .B2(new_n785), .ZN(new_n847));
  OAI22_X1  g0647(.A1(new_n781), .A2(new_n493), .B1(new_n784), .B2(new_n489), .ZN(new_n848));
  NOR4_X1   g0648(.A1(new_n845), .A2(new_n846), .A3(new_n847), .A4(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n784), .ZN(new_n850));
  AOI22_X1  g0650(.A1(G143), .A2(new_n843), .B1(new_n850), .B2(G159), .ZN(new_n851));
  INV_X1    g0651(.A(G150), .ZN(new_n852));
  INV_X1    g0652(.A(G137), .ZN(new_n853));
  OAI221_X1 g0653(.A(new_n851), .B1(new_n852), .B2(new_n798), .C1(new_n795), .C2(new_n853), .ZN(new_n854));
  XNOR2_X1  g0654(.A(new_n854), .B(KEYINPUT34), .ZN(new_n855));
  INV_X1    g0655(.A(G132), .ZN(new_n856));
  OAI22_X1  g0656(.A1(new_n777), .A2(new_n309), .B1(new_n788), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n244), .B1(new_n781), .B2(new_n307), .ZN(new_n858));
  AOI211_X1 g0658(.A(new_n857), .B(new_n858), .C1(G58), .C2(new_n808), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n849), .B1(new_n855), .B2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n835), .ZN(new_n861));
  OAI221_X1 g0661(.A(new_n841), .B1(new_n842), .B2(new_n860), .C1(new_n861), .C2(new_n770), .ZN(new_n862));
  AND2_X1   g0662(.A1(new_n839), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(G384));
  OR2_X1    g0664(.A1(new_n527), .A2(KEYINPUT35), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n527), .A2(KEYINPUT35), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n865), .A2(new_n866), .A3(G116), .A4(new_n222), .ZN(new_n867));
  XOR2_X1   g0667(.A(new_n867), .B(KEYINPUT36), .Z(new_n868));
  OAI211_X1 g0668(.A(new_n220), .B(G77), .C1(new_n308), .C2(new_n309), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n307), .A2(G68), .ZN(new_n870));
  AOI211_X1 g0670(.A(new_n203), .B(G13), .C1(new_n869), .C2(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  OR2_X1    g0672(.A1(KEYINPUT102), .A2(KEYINPUT31), .ZN(new_n873));
  OR2_X1    g0673(.A1(new_n747), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n747), .A2(new_n873), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NOR3_X1   g0676(.A1(new_n517), .A2(new_n729), .A3(new_n693), .ZN(new_n877));
  AOI21_X1  g0677(.A(KEYINPUT92), .B1(new_n877), .B2(new_n677), .ZN(new_n878));
  NOR4_X1   g0678(.A1(new_n633), .A2(new_n517), .A3(new_n732), .A4(new_n683), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n876), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n450), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n448), .A2(new_n683), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n881), .A2(new_n637), .A3(new_n882), .ZN(new_n883));
  OAI211_X1 g0683(.A(new_n448), .B(new_n683), .C1(new_n457), .C2(new_n450), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n861), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n880), .A2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT37), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n363), .A2(new_n368), .A3(new_n316), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n371), .ZN(new_n891));
  AOI22_X1  g0691(.A1(new_n410), .A2(new_n415), .B1(new_n891), .B2(new_n676), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n394), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n889), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n372), .A2(new_n676), .ZN(new_n895));
  NAND4_X1  g0695(.A1(new_n395), .A2(new_n895), .A3(new_n889), .A4(new_n403), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(KEYINPUT38), .B1(new_n894), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n642), .B1(new_n640), .B2(new_n639), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n891), .A2(new_n676), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n898), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  XOR2_X1   g0702(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  AND2_X1   g0704(.A1(new_n395), .A2(new_n403), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT100), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n905), .A2(new_n906), .A3(new_n889), .A4(new_n895), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n395), .A2(new_n895), .A3(new_n403), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(KEYINPUT37), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n896), .A2(KEYINPUT100), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n907), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n418), .A2(new_n420), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n372), .B(new_n676), .C1(new_n399), .C2(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n904), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(KEYINPUT40), .B1(new_n902), .B2(new_n914), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n888), .A2(new_n915), .ZN(new_n916));
  OAI22_X1  g0716(.A1(new_n422), .A2(new_n900), .B1(new_n897), .B2(new_n894), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT38), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT98), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n900), .A2(new_n893), .A3(new_n403), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(KEYINPUT37), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n918), .B1(new_n922), .B2(new_n896), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n920), .B(new_n923), .C1(new_n422), .C2(new_n900), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n899), .A2(new_n901), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n920), .B1(new_n926), .B2(new_n923), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n919), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  AOI22_X1  g0728(.A1(new_n733), .A2(new_n735), .B1(new_n874), .B2(new_n875), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n929), .A2(new_n886), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  XNOR2_X1  g0731(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n916), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  NOR3_X1   g0734(.A1(new_n934), .A2(new_n459), .A3(new_n929), .ZN(new_n935));
  INV_X1    g0735(.A(new_n459), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n933), .B1(new_n936), .B2(new_n880), .ZN(new_n937));
  NOR3_X1   g0737(.A1(new_n935), .A2(new_n727), .A3(new_n937), .ZN(new_n938));
  AND2_X1   g0738(.A1(new_n883), .A2(new_n884), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n939), .B1(new_n829), .B2(new_n834), .ZN(new_n940));
  AOI22_X1  g0740(.A1(new_n928), .A2(new_n940), .B1(new_n399), .B2(new_n675), .ZN(new_n941));
  OAI211_X1 g0741(.A(KEYINPUT39), .B(new_n919), .C1(new_n925), .C2(new_n927), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n911), .A2(new_n913), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(new_n903), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n923), .B1(new_n422), .B2(new_n900), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT39), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n457), .A2(new_n448), .A3(new_n677), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n942), .A2(new_n948), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n941), .A2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n645), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n715), .A2(KEYINPUT93), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n954), .A2(new_n723), .A3(KEYINPUT29), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n725), .A2(new_n710), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n953), .B1(new_n957), .B2(new_n936), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n952), .B(new_n958), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n938), .A2(new_n959), .B1(new_n203), .B2(new_n757), .ZN(new_n960));
  AND2_X1   g0760(.A1(new_n938), .A2(new_n959), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n872), .B1(new_n960), .B2(new_n961), .ZN(G367));
  OAI21_X1  g0762(.A(new_n773), .B1(new_n216), .B2(new_n274), .ZN(new_n963));
  INV_X1    g0763(.A(new_n765), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n963), .B1(new_n234), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n796), .A2(G143), .ZN(new_n966));
  AOI22_X1  g0766(.A1(G50), .A2(new_n850), .B1(new_n789), .B2(G137), .ZN(new_n967));
  OAI221_X1 g0767(.A(new_n967), .B1(new_n308), .B2(new_n781), .C1(new_n852), .C2(new_n804), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n244), .B1(new_n777), .B2(new_n279), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(KEYINPUT108), .ZN(new_n970));
  INV_X1    g0770(.A(G159), .ZN(new_n971));
  OAI22_X1  g0771(.A1(new_n798), .A2(new_n971), .B1(new_n807), .B2(new_n309), .ZN(new_n972));
  NOR3_X1   g0772(.A1(new_n968), .A2(new_n970), .A3(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(G294), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n798), .A2(new_n974), .ZN(new_n975));
  OAI221_X1 g0775(.A(new_n355), .B1(new_n807), .B2(new_n493), .C1(new_n800), .C2(new_n788), .ZN(new_n976));
  AOI211_X1 g0776(.A(new_n975), .B(new_n976), .C1(new_n796), .C2(G311), .ZN(new_n977));
  INV_X1    g0777(.A(new_n566), .ZN(new_n978));
  AOI22_X1  g0778(.A1(new_n843), .A2(new_n978), .B1(new_n850), .B2(G283), .ZN(new_n979));
  INV_X1    g0779(.A(new_n777), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(G97), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT107), .ZN(new_n982));
  INV_X1    g0782(.A(new_n781), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n982), .B1(new_n983), .B2(G116), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT46), .ZN(new_n985));
  OAI211_X1 g0785(.A(new_n979), .B(new_n981), .C1(new_n984), .C2(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n986), .B1(new_n985), .B2(new_n984), .ZN(new_n987));
  AOI22_X1  g0787(.A1(new_n966), .A2(new_n973), .B1(new_n977), .B2(new_n987), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n988), .B(KEYINPUT47), .Z(new_n989));
  AOI211_X1 g0789(.A(new_n824), .B(new_n965), .C1(new_n989), .C2(new_n772), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n613), .A2(new_n677), .ZN(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(new_n654), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(new_n646), .B2(new_n992), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n990), .B1(new_n821), .B2(new_n994), .ZN(new_n995));
  OAI211_X1 g0795(.A(new_n695), .B(new_n700), .C1(new_n689), .C2(new_n699), .ZN(new_n996));
  AOI211_X1 g0796(.A(new_n678), .B(new_n699), .C1(new_n685), .C2(new_n687), .ZN(new_n997));
  INV_X1    g0797(.A(new_n700), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n696), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n996), .A2(new_n999), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n726), .A2(new_n1000), .A3(new_n753), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(KEYINPUT106), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT105), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT44), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n656), .A2(new_n683), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n728), .A2(new_n658), .A3(new_n1007), .ZN(new_n1008));
  OR2_X1    g0808(.A1(new_n1008), .A2(KEYINPUT103), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n665), .A2(new_n683), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1008), .A2(KEYINPUT103), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1009), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1012), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n700), .A2(new_n698), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1006), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT45), .ZN(new_n1017));
  AND3_X1   g0817(.A1(new_n1009), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1017), .B1(new_n1014), .B2(new_n1018), .ZN(new_n1019));
  NAND4_X1  g0819(.A1(new_n700), .A2(KEYINPUT45), .A3(new_n698), .A4(new_n1012), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1013), .A2(new_n1014), .A3(new_n1006), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1016), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n697), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT106), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n726), .A2(new_n1000), .A3(new_n1026), .A4(new_n753), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n1022), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n1028), .A2(new_n1015), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1029), .A2(new_n697), .A3(new_n1021), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n1002), .A2(new_n1025), .A3(new_n1027), .A4(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1031), .A2(new_n755), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n705), .B(KEYINPUT41), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n759), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n994), .A2(KEYINPUT43), .ZN(new_n1035));
  OAI21_X1  g0835(.A(KEYINPUT42), .B1(new_n1018), .B2(new_n700), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n508), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n677), .B1(new_n1037), .B2(new_n665), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1039));
  NOR3_X1   g0839(.A1(new_n1018), .A2(new_n700), .A3(KEYINPUT42), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1035), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(KEYINPUT104), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n994), .A2(KEYINPUT43), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT104), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n1044), .B(new_n1035), .C1(new_n1039), .C2(new_n1040), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1042), .A2(new_n1043), .A3(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1043), .B1(new_n1042), .B2(new_n1045), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n1047), .A2(new_n1048), .B1(new_n697), .B2(new_n1018), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1048), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n697), .A2(new_n1018), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1050), .A2(new_n1051), .A3(new_n1046), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1049), .A2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n995), .B1(new_n1034), .B2(new_n1053), .ZN(G387));
  NAND2_X1  g0854(.A1(new_n1000), .A2(new_n759), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n781), .A2(new_n279), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(G68), .B2(new_n850), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n1057), .B1(new_n307), .B2(new_n804), .C1(new_n852), .C2(new_n788), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n795), .A2(new_n971), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n807), .A2(new_n274), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n981), .B(new_n244), .C1(new_n276), .C2(new_n798), .ZN(new_n1061));
  NOR4_X1   g0861(.A1(new_n1058), .A2(new_n1059), .A3(new_n1060), .A4(new_n1061), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT110), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n796), .A2(G322), .B1(G311), .B2(new_n799), .ZN(new_n1064));
  OR2_X1    g0864(.A1(new_n1064), .A2(KEYINPUT111), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1064), .A2(KEYINPUT111), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n843), .A2(G317), .B1(new_n850), .B2(new_n978), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1065), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT48), .ZN(new_n1069));
  OR2_X1    g0869(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n781), .A2(new_n974), .B1(new_n807), .B2(new_n778), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1072));
  XOR2_X1   g0872(.A(KEYINPUT112), .B(KEYINPUT49), .Z(new_n1073));
  NAND3_X1  g0873(.A1(new_n1070), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n244), .B1(new_n789), .B2(G326), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1074), .B(new_n1075), .C1(new_n489), .C2(new_n777), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1073), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1063), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(new_n772), .ZN(new_n1079));
  AOI211_X1 g0879(.A(G45), .B(new_n706), .C1(G68), .C2(G77), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1080), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n1081), .A2(KEYINPUT109), .ZN(new_n1082));
  OAI21_X1  g0882(.A(KEYINPUT50), .B1(new_n276), .B2(G50), .ZN(new_n1083));
  OR3_X1    g0883(.A1(new_n276), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT109), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1083), .B(new_n1084), .C1(new_n1080), .C2(new_n1085), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n964), .B1(new_n1082), .B2(new_n1086), .C1(new_n230), .C2(new_n766), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n706), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n1087), .B1(G107), .B2(new_n216), .C1(new_n1088), .C2(new_n761), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n824), .B1(new_n1089), .B2(new_n773), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1079), .B(new_n1090), .C1(new_n689), .C2(new_n821), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1001), .A2(KEYINPUT113), .A3(new_n705), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1092), .B1(new_n755), .B2(new_n1000), .ZN(new_n1093));
  AOI21_X1  g0893(.A(KEYINPUT113), .B1(new_n1001), .B2(new_n705), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1055), .B(new_n1091), .C1(new_n1093), .C2(new_n1094), .ZN(G393));
  INV_X1    g0895(.A(KEYINPUT115), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n697), .B1(new_n1029), .B2(new_n1021), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1001), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n705), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1031), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1096), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n1099), .A2(new_n1031), .A3(KEYINPUT115), .A4(new_n705), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1018), .A2(new_n771), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n773), .B1(new_n518), .B2(new_n216), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1106), .B1(new_n242), .B2(new_n964), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n795), .A2(new_n800), .B1(new_n785), .B2(new_n804), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1108), .B(KEYINPUT52), .ZN(new_n1109));
  OAI221_X1 g0909(.A(new_n355), .B1(new_n777), .B2(new_n493), .C1(new_n566), .C2(new_n798), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n983), .A2(G283), .B1(new_n850), .B2(G294), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1111), .B1(new_n805), .B2(new_n788), .ZN(new_n1112));
  AOI211_X1 g0912(.A(new_n1110), .B(new_n1112), .C1(G116), .C2(new_n808), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1109), .A2(new_n1113), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n795), .A2(new_n852), .B1(new_n971), .B2(new_n804), .ZN(new_n1115));
  XOR2_X1   g0915(.A(new_n1115), .B(KEYINPUT51), .Z(new_n1116));
  NOR2_X1   g0916(.A1(new_n781), .A2(new_n309), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n244), .B1(new_n777), .B2(new_n597), .ZN(new_n1118));
  AOI211_X1 g0918(.A(new_n1117), .B(new_n1118), .C1(G143), .C2(new_n789), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n276), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n799), .A2(G50), .B1(new_n850), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT114), .ZN(new_n1122));
  OR2_X1    g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n807), .A2(new_n279), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1119), .A2(new_n1123), .A3(new_n1124), .A4(new_n1126), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1114), .B1(new_n1116), .B2(new_n1127), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n824), .B(new_n1107), .C1(new_n1128), .C2(new_n772), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1105), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1025), .A2(new_n1030), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1130), .B1(new_n1131), .B2(new_n758), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1104), .A2(new_n1133), .ZN(G390));
  INV_X1    g0934(.A(new_n834), .ZN(new_n1135));
  OR2_X1    g0935(.A1(new_n718), .A2(new_n719), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n718), .A2(new_n719), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1136), .A2(new_n1137), .A3(new_n717), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n711), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n683), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1135), .B1(new_n1140), .B2(new_n833), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n949), .B(new_n946), .C1(new_n1141), .C2(new_n939), .ZN(new_n1142));
  AOI21_X1  g0942(.A(KEYINPUT39), .B1(new_n944), .B2(new_n945), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n945), .A2(KEYINPUT98), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n1144), .A2(new_n924), .B1(new_n918), .B2(new_n917), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1143), .B1(new_n1145), .B2(KEYINPUT39), .ZN(new_n1146));
  OAI21_X1  g0946(.A(KEYINPUT116), .B1(new_n940), .B2(new_n950), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT116), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1135), .B1(new_n669), .B2(new_n828), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n1148), .B(new_n949), .C1(new_n1149), .C2(new_n939), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1147), .A2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1142), .B1(new_n1146), .B2(new_n1151), .ZN(new_n1152));
  NOR3_X1   g0952(.A1(new_n929), .A2(new_n727), .A3(new_n886), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n751), .B1(new_n878), .B2(new_n879), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n1155), .A2(new_n885), .A3(G330), .A4(new_n861), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n1142), .B(new_n1156), .C1(new_n1146), .C2(new_n1151), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1154), .A2(new_n1157), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1158), .A2(new_n758), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n942), .A2(new_n948), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1160), .A2(new_n769), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n840), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n760), .B1(new_n1120), .B2(new_n1162), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n355), .B1(new_n781), .B2(new_n597), .ZN(new_n1164));
  AOI211_X1 g0964(.A(new_n1125), .B(new_n1164), .C1(G107), .C2(new_n799), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n777), .A2(new_n309), .B1(new_n784), .B2(new_n518), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n804), .A2(new_n489), .B1(new_n788), .B2(new_n974), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n1165), .B(new_n1168), .C1(new_n778), .C2(new_n795), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n781), .A2(new_n852), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT53), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n1170), .A2(new_n1171), .B1(new_n853), .B2(new_n798), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(new_n1171), .B2(new_n1170), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n307), .A2(new_n777), .B1(new_n804), .B2(new_n856), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(G125), .B2(new_n789), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(KEYINPUT54), .B(G143), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n244), .B1(new_n784), .B2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(G159), .B2(new_n808), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1173), .A2(new_n1175), .A3(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(G128), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n795), .A2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1169), .B1(new_n1179), .B2(new_n1181), .ZN(new_n1182));
  OR2_X1    g0982(.A1(new_n1182), .A2(KEYINPUT118), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n842), .B1(new_n1182), .B2(KEYINPUT118), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1163), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1159), .B1(new_n1161), .B2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n705), .ZN(new_n1187));
  NOR3_X1   g0987(.A1(new_n929), .A2(new_n727), .A3(new_n835), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n1141), .B(new_n1156), .C1(new_n1188), .C2(new_n885), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1155), .A2(G330), .A3(new_n861), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n727), .B1(new_n736), .B2(new_n876), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n1190), .A2(new_n939), .B1(new_n1191), .B2(new_n887), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1189), .B1(new_n1149), .B2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1191), .A2(new_n936), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n645), .B(new_n1194), .C1(new_n726), .C2(new_n459), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1193), .A2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1187), .B1(new_n1158), .B2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n885), .B1(new_n752), .B2(new_n861), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n1199), .A2(new_n1153), .B1(new_n830), .B2(new_n1135), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1195), .B1(new_n1200), .B2(new_n1189), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1154), .A2(new_n1201), .A3(new_n1157), .ZN(new_n1202));
  AOI21_X1  g1002(.A(KEYINPUT117), .B1(new_n1198), .B2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1157), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1153), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1160), .A2(new_n1147), .A3(new_n1150), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1205), .B1(new_n1206), .B2(new_n1142), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1197), .B1(new_n1204), .B2(new_n1207), .ZN(new_n1208));
  AND4_X1   g1008(.A1(KEYINPUT117), .A2(new_n1208), .A3(new_n705), .A4(new_n1202), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1186), .B1(new_n1203), .B2(new_n1209), .ZN(G378));
  INV_X1    g1010(.A(KEYINPUT57), .ZN(new_n1211));
  AND2_X1   g1011(.A1(new_n1202), .A2(new_n1196), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n932), .B1(new_n1145), .B2(new_n888), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n930), .A2(KEYINPUT40), .A3(new_n946), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1213), .A2(G330), .A3(new_n1214), .ZN(new_n1215));
  XOR2_X1   g1015(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n339), .A2(new_n341), .A3(new_n321), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n324), .A2(new_n675), .ZN(new_n1219));
  OR2_X1    g1019(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT121), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1220), .A2(new_n1221), .A3(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1221), .B1(new_n1220), .B2(new_n1222), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1217), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1225), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1227), .A2(new_n1216), .A3(new_n1223), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1226), .A2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1215), .A2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n952), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1213), .A2(new_n1229), .A3(G330), .A4(new_n1214), .ZN(new_n1233));
  AND3_X1   g1033(.A1(new_n1231), .A2(new_n1232), .A3(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1232), .B1(new_n1231), .B2(new_n1233), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1211), .B1(new_n1212), .B2(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1229), .B1(new_n933), .B2(G330), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1233), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n952), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT122), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1231), .A2(new_n1232), .A3(new_n1233), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1240), .A2(new_n1241), .A3(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1202), .A2(new_n1196), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1235), .A2(KEYINPUT122), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1243), .A2(KEYINPUT57), .A3(new_n1244), .A4(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1237), .A2(new_n1246), .A3(new_n705), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1240), .A2(new_n1242), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1230), .A2(new_n769), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n760), .B1(G50), .B2(new_n1162), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n796), .A2(G116), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n777), .A2(new_n308), .ZN(new_n1252));
  OAI22_X1  g1052(.A1(new_n804), .A2(new_n493), .B1(new_n784), .B2(new_n274), .ZN(new_n1253));
  AOI211_X1 g1053(.A(new_n1252), .B(new_n1253), .C1(G283), .C2(new_n789), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n799), .A2(G97), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n355), .A2(new_n252), .ZN(new_n1256));
  AOI211_X1 g1056(.A(new_n1256), .B(new_n1056), .C1(G68), .C2(new_n808), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1251), .A2(new_n1254), .A3(new_n1255), .A4(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT58), .ZN(new_n1259));
  AOI21_X1  g1059(.A(G50), .B1(new_n270), .B2(new_n252), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(new_n1258), .A2(new_n1259), .B1(new_n1256), .B2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n796), .A2(G125), .ZN(new_n1262));
  OAI22_X1  g1062(.A1(new_n781), .A2(new_n1176), .B1(new_n804), .B2(new_n1180), .ZN(new_n1263));
  XNOR2_X1  g1063(.A(new_n1263), .B(KEYINPUT119), .ZN(new_n1264));
  OAI22_X1  g1064(.A1(new_n784), .A2(new_n853), .B1(new_n807), .B2(new_n852), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1265), .B1(G132), .B2(new_n799), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1262), .A2(new_n1264), .A3(new_n1266), .ZN(new_n1267));
  XOR2_X1   g1067(.A(new_n1267), .B(KEYINPUT120), .Z(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1269), .A2(KEYINPUT59), .ZN(new_n1270));
  OAI211_X1 g1070(.A(new_n270), .B(new_n252), .C1(new_n777), .C2(new_n971), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1271), .B1(G124), .B2(new_n789), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT59), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1272), .B1(new_n1268), .B2(new_n1273), .ZN(new_n1274));
  OAI221_X1 g1074(.A(new_n1261), .B1(new_n1259), .B2(new_n1258), .C1(new_n1270), .C2(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1250), .B1(new_n1275), .B2(new_n772), .ZN(new_n1276));
  AOI22_X1  g1076(.A1(new_n1248), .A2(new_n759), .B1(new_n1249), .B2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1247), .A2(new_n1277), .ZN(G375));
  NAND3_X1  g1078(.A1(new_n1200), .A2(new_n1195), .A3(new_n1189), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1197), .A2(new_n1033), .A3(new_n1279), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n760), .B1(G68), .B2(new_n1162), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n885), .A2(new_n770), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n355), .B1(new_n777), .B2(new_n279), .ZN(new_n1283));
  AOI211_X1 g1083(.A(new_n1060), .B(new_n1283), .C1(G116), .C2(new_n799), .ZN(new_n1284));
  OAI22_X1  g1084(.A1(new_n781), .A2(new_n518), .B1(new_n788), .B2(new_n782), .ZN(new_n1285));
  OAI22_X1  g1085(.A1(new_n804), .A2(new_n778), .B1(new_n784), .B2(new_n493), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  OAI211_X1 g1087(.A(new_n1284), .B(new_n1287), .C1(new_n974), .C2(new_n795), .ZN(new_n1288));
  OR2_X1    g1088(.A1(new_n1288), .A2(KEYINPUT123), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(KEYINPUT123), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n796), .A2(G132), .ZN(new_n1291));
  OAI22_X1  g1091(.A1(new_n781), .A2(new_n971), .B1(new_n788), .B2(new_n1180), .ZN(new_n1292));
  OAI22_X1  g1092(.A1(new_n804), .A2(new_n853), .B1(new_n784), .B2(new_n852), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n808), .A2(G50), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n798), .A2(new_n1176), .ZN(new_n1296));
  NOR3_X1   g1096(.A1(new_n1296), .A2(new_n1252), .A3(new_n355), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1291), .A2(new_n1294), .A3(new_n1295), .A4(new_n1297), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1289), .A2(new_n1290), .A3(new_n1298), .ZN(new_n1299));
  AOI211_X1 g1099(.A(new_n1281), .B(new_n1282), .C1(new_n772), .C2(new_n1299), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1300), .B1(new_n1193), .B2(new_n759), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1280), .A2(new_n1301), .ZN(G381));
  NAND2_X1  g1102(.A1(new_n1198), .A2(new_n1202), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1186), .A2(new_n1303), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1280), .A2(new_n863), .A3(new_n1301), .ZN(new_n1305));
  OR2_X1    g1105(.A1(G393), .A2(G396), .ZN(new_n1306));
  NOR4_X1   g1106(.A1(new_n1304), .A2(G390), .A3(new_n1305), .A4(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(G387), .ZN(new_n1308));
  NAND4_X1  g1108(.A1(new_n1307), .A2(new_n1308), .A3(new_n1247), .A4(new_n1277), .ZN(G407));
  INV_X1    g1109(.A(new_n1304), .ZN(new_n1310));
  INV_X1    g1110(.A(G213), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1311), .A2(G343), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1310), .A2(new_n1312), .ZN(new_n1313));
  OAI211_X1 g1113(.A(G407), .B(G213), .C1(G375), .C2(new_n1313), .ZN(new_n1314));
  XNOR2_X1  g1114(.A(new_n1314), .B(KEYINPUT124), .ZN(G409));
  INV_X1    g1115(.A(KEYINPUT60), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1279), .A2(new_n1316), .ZN(new_n1317));
  NAND4_X1  g1117(.A1(new_n1200), .A2(new_n1195), .A3(KEYINPUT60), .A4(new_n1189), .ZN(new_n1318));
  NAND4_X1  g1118(.A1(new_n1317), .A2(new_n705), .A3(new_n1197), .A4(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1319), .A2(new_n1301), .ZN(new_n1320));
  OR2_X1    g1120(.A1(new_n863), .A2(KEYINPUT125), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n863), .A2(KEYINPUT125), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1320), .A2(new_n1321), .A3(new_n1322), .ZN(new_n1323));
  NAND4_X1  g1123(.A1(new_n1319), .A2(KEYINPUT125), .A3(new_n863), .A4(new_n1301), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1325), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1247), .A2(G378), .A3(new_n1277), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1243), .A2(new_n759), .A3(new_n1245), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1248), .A2(new_n1244), .A3(new_n1033), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1249), .A2(new_n1276), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1328), .A2(new_n1329), .A3(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1310), .A2(new_n1331), .ZN(new_n1332));
  AOI211_X1 g1132(.A(new_n1312), .B(new_n1326), .C1(new_n1327), .C2(new_n1332), .ZN(new_n1333));
  OAI21_X1  g1133(.A(KEYINPUT63), .B1(new_n1333), .B2(KEYINPUT126), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1308), .A2(G390), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(G393), .A2(G396), .ZN(new_n1336));
  AOI21_X1  g1136(.A(new_n1132), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1337), .A2(G387), .ZN(new_n1338));
  NAND4_X1  g1138(.A1(new_n1335), .A2(new_n1306), .A3(new_n1336), .A4(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1306), .A2(new_n1336), .ZN(new_n1340));
  AND2_X1   g1140(.A1(new_n1337), .A2(G387), .ZN(new_n1341));
  NOR2_X1   g1141(.A1(new_n1337), .A2(G387), .ZN(new_n1342));
  OAI21_X1  g1142(.A(new_n1340), .B1(new_n1341), .B2(new_n1342), .ZN(new_n1343));
  INV_X1    g1143(.A(KEYINPUT61), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1339), .A2(new_n1343), .A3(new_n1344), .ZN(new_n1345));
  AOI21_X1  g1145(.A(new_n1312), .B1(new_n1327), .B2(new_n1332), .ZN(new_n1346));
  INV_X1    g1146(.A(new_n1346), .ZN(new_n1347));
  AOI21_X1  g1147(.A(new_n1325), .B1(G2897), .B2(new_n1312), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1312), .A2(G2897), .ZN(new_n1349));
  AOI21_X1  g1149(.A(new_n1349), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1350));
  NOR2_X1   g1150(.A1(new_n1348), .A2(new_n1350), .ZN(new_n1351));
  INV_X1    g1151(.A(new_n1351), .ZN(new_n1352));
  AOI21_X1  g1152(.A(new_n1345), .B1(new_n1347), .B2(new_n1352), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1346), .A2(new_n1325), .ZN(new_n1354));
  INV_X1    g1154(.A(KEYINPUT126), .ZN(new_n1355));
  INV_X1    g1155(.A(KEYINPUT63), .ZN(new_n1356));
  NAND3_X1  g1156(.A1(new_n1354), .A2(new_n1355), .A3(new_n1356), .ZN(new_n1357));
  NAND3_X1  g1157(.A1(new_n1334), .A2(new_n1353), .A3(new_n1357), .ZN(new_n1358));
  INV_X1    g1158(.A(KEYINPUT62), .ZN(new_n1359));
  AND3_X1   g1159(.A1(new_n1346), .A2(new_n1359), .A3(new_n1325), .ZN(new_n1360));
  XOR2_X1   g1160(.A(KEYINPUT127), .B(KEYINPUT61), .Z(new_n1361));
  OAI21_X1  g1161(.A(new_n1361), .B1(new_n1346), .B2(new_n1351), .ZN(new_n1362));
  AOI21_X1  g1162(.A(new_n1359), .B1(new_n1346), .B2(new_n1325), .ZN(new_n1363));
  NOR3_X1   g1163(.A1(new_n1360), .A2(new_n1362), .A3(new_n1363), .ZN(new_n1364));
  AND2_X1   g1164(.A1(new_n1339), .A2(new_n1343), .ZN(new_n1365));
  OAI21_X1  g1165(.A(new_n1358), .B1(new_n1364), .B2(new_n1365), .ZN(G405));
  INV_X1    g1166(.A(new_n1327), .ZN(new_n1367));
  AOI21_X1  g1167(.A(new_n1304), .B1(new_n1247), .B2(new_n1277), .ZN(new_n1368));
  OAI21_X1  g1168(.A(new_n1365), .B1(new_n1367), .B2(new_n1368), .ZN(new_n1369));
  NOR2_X1   g1169(.A1(new_n1367), .A2(new_n1368), .ZN(new_n1370));
  NAND2_X1  g1170(.A1(new_n1339), .A2(new_n1343), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1370), .A2(new_n1371), .ZN(new_n1372));
  AND3_X1   g1172(.A1(new_n1369), .A2(new_n1326), .A3(new_n1372), .ZN(new_n1373));
  AOI21_X1  g1173(.A(new_n1326), .B1(new_n1369), .B2(new_n1372), .ZN(new_n1374));
  NOR2_X1   g1174(.A1(new_n1373), .A2(new_n1374), .ZN(G402));
endmodule


