//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 0 0 0 0 1 0 0 0 0 0 0 1 1 0 0 0 0 1 1 1 0 0 1 1 1 0 0 0 1 0 1 0 1 0 1 1 0 0 1 1 0 1 1 1 0 0 0 1 1 1 1 0 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:12 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  INV_X1    g0001(.A(G97), .ZN(new_n202));
  INV_X1    g0002(.A(G107), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(G87), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n207), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT64), .ZN(new_n215));
  OAI21_X1  g0015(.A(G50), .B1(G58), .B2(G68), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT65), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  AND2_X1   g0020(.A1(new_n220), .A2(KEYINPUT66), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(KEYINPUT66), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n219), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  OR2_X1    g0023(.A1(new_n223), .A2(KEYINPUT67), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n223), .A2(KEYINPUT67), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n228));
  NAND3_X1  g0028(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n209), .B1(new_n225), .B2(new_n229), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n212), .B1(new_n215), .B2(new_n218), .C1(new_n230), .C2(KEYINPUT1), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n230), .ZN(G361));
  XOR2_X1   g0032(.A(G250), .B(G257), .Z(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(KEYINPUT69), .B(KEYINPUT70), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G238), .B(G244), .Z(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G226), .B(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n237), .B(new_n242), .ZN(G358));
  XOR2_X1   g0043(.A(G68), .B(G77), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT71), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G107), .B(G116), .Z(new_n248));
  XNOR2_X1  g0048(.A(G87), .B(G97), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n247), .B(new_n250), .Z(G351));
  NAND2_X1  g0051(.A1(new_n208), .A2(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(new_n213), .ZN(new_n253));
  INV_X1    g0053(.A(G13), .ZN(new_n254));
  NOR3_X1   g0054(.A1(new_n254), .A2(new_n207), .A3(G1), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(KEYINPUT72), .ZN(new_n257));
  AOI22_X1  g0057(.A1(new_n208), .A2(G33), .B1(G1), .B2(G13), .ZN(new_n258));
  INV_X1    g0058(.A(new_n255), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT72), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  AND2_X1   g0062(.A1(new_n257), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n206), .A2(G20), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n263), .A2(G68), .A3(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G68), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n255), .A2(new_n266), .ZN(new_n267));
  XOR2_X1   g0067(.A(new_n267), .B(KEYINPUT12), .Z(new_n268));
  INV_X1    g0068(.A(G33), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n269), .A2(G20), .ZN(new_n270));
  AOI22_X1  g0070(.A1(new_n270), .A2(G77), .B1(G20), .B2(new_n266), .ZN(new_n271));
  INV_X1    g0071(.A(G50), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n207), .A2(new_n269), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n271), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  AND2_X1   g0074(.A1(new_n274), .A2(new_n253), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n268), .B1(KEYINPUT11), .B2(new_n275), .ZN(new_n276));
  OAI211_X1 g0076(.A(new_n265), .B(new_n276), .C1(KEYINPUT11), .C2(new_n275), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT76), .ZN(new_n278));
  XNOR2_X1  g0078(.A(new_n277), .B(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(G33), .A2(G41), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n280), .A2(G1), .A3(G13), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G274), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G232), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G1698), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n286), .B1(G226), .B2(G1698), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n269), .A2(KEYINPUT3), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT3), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G33), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  OAI22_X1  g0091(.A1(new_n287), .A2(new_n291), .B1(new_n269), .B2(new_n202), .ZN(new_n292));
  INV_X1    g0092(.A(new_n281), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n284), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n281), .A2(new_n283), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  AND2_X1   g0096(.A1(new_n296), .A2(KEYINPUT75), .ZN(new_n297));
  OAI21_X1  g0097(.A(G238), .B1(new_n296), .B2(KEYINPUT75), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n294), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  XNOR2_X1  g0099(.A(new_n299), .B(KEYINPUT13), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(G200), .ZN(new_n301));
  INV_X1    g0101(.A(G190), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n301), .B1(new_n302), .B2(new_n300), .ZN(new_n303));
  OR2_X1    g0103(.A1(new_n279), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n300), .A2(G169), .ZN(new_n305));
  INV_X1    g0105(.A(G179), .ZN(new_n306));
  OAI22_X1  g0106(.A1(new_n305), .A2(KEYINPUT14), .B1(new_n306), .B2(new_n300), .ZN(new_n307));
  AND2_X1   g0107(.A1(new_n305), .A2(KEYINPUT14), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n279), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  AND2_X1   g0109(.A1(new_n304), .A2(new_n309), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n284), .B1(G244), .B2(new_n296), .ZN(new_n311));
  XNOR2_X1  g0111(.A(KEYINPUT3), .B(G33), .ZN(new_n312));
  NOR2_X1   g0112(.A1(G232), .A2(G1698), .ZN(new_n313));
  INV_X1    g0113(.A(G1698), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n314), .A2(G238), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n312), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n316), .B(new_n293), .C1(G107), .C2(new_n312), .ZN(new_n317));
  AND2_X1   g0117(.A1(new_n311), .A2(new_n317), .ZN(new_n318));
  OAI21_X1  g0118(.A(KEYINPUT73), .B1(new_n318), .B2(G169), .ZN(new_n319));
  INV_X1    g0119(.A(new_n318), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n319), .B1(G179), .B2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n318), .A2(KEYINPUT73), .A3(new_n306), .ZN(new_n322));
  AND2_X1   g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n263), .A2(G77), .A3(new_n264), .ZN(new_n324));
  XNOR2_X1  g0124(.A(KEYINPUT15), .B(G87), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n326), .A2(new_n270), .B1(G20), .B2(G77), .ZN(new_n327));
  XNOR2_X1  g0127(.A(KEYINPUT8), .B(G58), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n327), .B1(new_n273), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(G77), .ZN(new_n330));
  AOI22_X1  g0130(.A1(new_n329), .A2(new_n253), .B1(new_n330), .B2(new_n255), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n324), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n323), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n320), .A2(G200), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n318), .A2(G190), .ZN(new_n335));
  NAND4_X1  g0135(.A1(new_n334), .A2(new_n324), .A3(new_n331), .A4(new_n335), .ZN(new_n336));
  AND2_X1   g0136(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  NOR2_X1   g0137(.A1(G50), .A2(G58), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n207), .B1(new_n338), .B2(new_n266), .ZN(new_n339));
  INV_X1    g0139(.A(G150), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n273), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n328), .ZN(new_n342));
  AOI211_X1 g0142(.A(new_n339), .B(new_n341), .C1(new_n342), .C2(new_n270), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n343), .A2(new_n258), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n264), .A2(G50), .ZN(new_n345));
  OAI22_X1  g0145(.A1(new_n260), .A2(new_n345), .B1(G50), .B2(new_n259), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  XOR2_X1   g0147(.A(new_n347), .B(KEYINPUT9), .Z(new_n348));
  INV_X1    g0148(.A(G226), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n295), .A2(new_n349), .ZN(new_n350));
  NOR2_X1   g0150(.A1(G222), .A2(G1698), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n314), .A2(G223), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n312), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n281), .B1(new_n291), .B2(new_n330), .ZN(new_n354));
  AOI211_X1 g0154(.A(new_n284), .B(new_n350), .C1(new_n353), .C2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(G200), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT74), .ZN(new_n358));
  AOI22_X1  g0158(.A1(new_n357), .A2(new_n358), .B1(G190), .B2(new_n355), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n348), .B(new_n359), .C1(new_n358), .C2(new_n357), .ZN(new_n360));
  XNOR2_X1  g0160(.A(new_n360), .B(KEYINPUT10), .ZN(new_n361));
  AND2_X1   g0161(.A1(new_n355), .A2(new_n306), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n355), .A2(G169), .ZN(new_n363));
  NOR3_X1   g0163(.A1(new_n362), .A2(new_n363), .A3(new_n347), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  AND4_X1   g0165(.A1(new_n310), .A2(new_n337), .A3(new_n361), .A4(new_n365), .ZN(new_n366));
  NOR2_X1   g0166(.A1(G223), .A2(G1698), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n367), .B1(new_n349), .B2(G1698), .ZN(new_n368));
  OAI21_X1  g0168(.A(KEYINPUT77), .B1(new_n289), .B2(G33), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT77), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n370), .A2(new_n269), .A3(KEYINPUT3), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n368), .A2(new_n369), .A3(new_n290), .A4(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(G33), .A2(G87), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n281), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  OAI22_X1  g0174(.A1(new_n285), .A2(new_n295), .B1(new_n282), .B2(new_n283), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n356), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n369), .A2(new_n371), .A3(new_n290), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n349), .A2(G1698), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n378), .B1(G223), .B2(G1698), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n373), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(new_n293), .ZN(new_n381));
  INV_X1    g0181(.A(new_n375), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n381), .A2(new_n382), .A3(new_n302), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n376), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n328), .B1(new_n206), .B2(G20), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n256), .A2(new_n385), .B1(new_n255), .B2(new_n328), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT16), .ZN(new_n387));
  INV_X1    g0187(.A(G58), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n388), .A2(new_n266), .ZN(new_n389));
  NOR2_X1   g0189(.A1(G58), .A2(G68), .ZN(new_n390));
  OAI21_X1  g0190(.A(G20), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n207), .A2(new_n269), .A3(G159), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n377), .A2(new_n207), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n266), .B1(new_n394), .B2(KEYINPUT7), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT7), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n377), .A2(new_n396), .A3(new_n207), .ZN(new_n397));
  AOI211_X1 g0197(.A(new_n387), .B(new_n393), .C1(new_n395), .C2(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n396), .B1(new_n312), .B2(G20), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n291), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n266), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n387), .B1(new_n401), .B2(new_n393), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(new_n253), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n384), .B(new_n386), .C1(new_n398), .C2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(KEYINPUT79), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n394), .A2(KEYINPUT7), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n406), .A2(G68), .A3(new_n397), .ZN(new_n407));
  INV_X1    g0207(.A(new_n393), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n407), .A2(KEYINPUT16), .A3(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n409), .A2(new_n253), .A3(new_n402), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT79), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n410), .A2(new_n411), .A3(new_n386), .A4(new_n384), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n405), .A2(KEYINPUT17), .A3(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT17), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n410), .A2(new_n414), .A3(new_n386), .A4(new_n384), .ZN(new_n415));
  AND2_X1   g0215(.A1(new_n415), .A2(KEYINPUT80), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n386), .B1(new_n398), .B2(new_n403), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n374), .A2(new_n375), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(G179), .ZN(new_n420));
  INV_X1    g0220(.A(G169), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n420), .B1(new_n421), .B2(new_n419), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n418), .A2(KEYINPUT18), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(KEYINPUT78), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT78), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n418), .A2(new_n422), .A3(new_n425), .A4(KEYINPUT18), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n418), .A2(new_n422), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT18), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n424), .A2(new_n426), .A3(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT80), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n405), .A2(new_n431), .A3(KEYINPUT17), .A4(new_n412), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n417), .A2(new_n430), .A3(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n366), .A2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT92), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n369), .A2(new_n371), .A3(new_n207), .A4(new_n290), .ZN(new_n437));
  NAND2_X1  g0237(.A1(KEYINPUT22), .A2(G87), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(G87), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n440), .A2(G20), .ZN(new_n441));
  AOI21_X1  g0241(.A(KEYINPUT22), .B1(new_n312), .B2(new_n441), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n436), .B1(new_n439), .B2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT22), .ZN(new_n444));
  INV_X1    g0244(.A(new_n441), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n444), .B1(new_n291), .B2(new_n445), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n446), .B(KEYINPUT92), .C1(new_n437), .C2(new_n438), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n443), .A2(new_n447), .ZN(new_n448));
  NOR3_X1   g0248(.A1(new_n207), .A2(KEYINPUT23), .A3(G107), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT23), .ZN(new_n450));
  OAI22_X1  g0250(.A1(new_n449), .A2(KEYINPUT93), .B1(new_n450), .B2(new_n203), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n450), .A2(new_n203), .A3(G20), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT93), .ZN(new_n453));
  AOI21_X1  g0253(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n454));
  OAI22_X1  g0254(.A1(new_n452), .A2(new_n453), .B1(new_n454), .B2(G20), .ZN(new_n455));
  OAI21_X1  g0255(.A(KEYINPUT94), .B1(new_n451), .B2(new_n455), .ZN(new_n456));
  AOI22_X1  g0256(.A1(new_n452), .A2(new_n453), .B1(KEYINPUT23), .B2(G107), .ZN(new_n457));
  OR2_X1    g0257(.A1(new_n454), .A2(G20), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT94), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n449), .A2(KEYINPUT93), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n457), .A2(new_n458), .A3(new_n459), .A4(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n456), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n448), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(KEYINPUT24), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT24), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n448), .A2(new_n465), .A3(new_n462), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n258), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n206), .A2(G33), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n256), .A2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT95), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(KEYINPUT25), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n203), .B1(new_n471), .B2(KEYINPUT25), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n472), .B1(new_n473), .B2(new_n259), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n255), .A2(new_n471), .A3(KEYINPUT25), .A4(new_n203), .ZN(new_n475));
  AOI22_X1  g0275(.A1(new_n470), .A2(G107), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n467), .A2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(G41), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n206), .B(G45), .C1(new_n479), .C2(KEYINPUT5), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT85), .ZN(new_n481));
  AND2_X1   g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n479), .A2(KEYINPUT5), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n483), .B1(new_n480), .B2(new_n481), .ZN(new_n484));
  OR3_X1    g0284(.A1(new_n482), .A2(new_n484), .A3(new_n282), .ZN(new_n485));
  OAI211_X1 g0285(.A(G264), .B(new_n281), .C1(new_n482), .C2(new_n484), .ZN(new_n486));
  INV_X1    g0286(.A(G257), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(G1698), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n488), .B1(G250), .B2(G1698), .ZN(new_n489));
  INV_X1    g0289(.A(G294), .ZN(new_n490));
  OAI22_X1  g0290(.A1(new_n377), .A2(new_n489), .B1(new_n269), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(new_n293), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n485), .A2(new_n486), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n421), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n494), .B1(G179), .B2(new_n493), .ZN(new_n495));
  OR2_X1    g0295(.A1(new_n478), .A2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT21), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n257), .A2(G116), .A3(new_n262), .A4(new_n468), .ZN(new_n498));
  INV_X1    g0298(.A(G116), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n255), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n258), .B1(G20), .B2(new_n499), .ZN(new_n501));
  NAND2_X1  g0301(.A1(G33), .A2(G283), .ZN(new_n502));
  OR2_X1    g0302(.A1(KEYINPUT81), .A2(G97), .ZN(new_n503));
  NAND2_X1  g0303(.A1(KEYINPUT81), .A2(G97), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n207), .B(new_n502), .C1(new_n506), .C2(G33), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n501), .A2(new_n507), .A3(KEYINPUT20), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(KEYINPUT20), .B1(new_n501), .B2(new_n507), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n498), .B(new_n500), .C1(new_n509), .C2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  OAI211_X1 g0312(.A(G270), .B(new_n281), .C1(new_n482), .C2(new_n484), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n487), .A2(new_n314), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n514), .B1(G264), .B2(new_n314), .ZN(new_n515));
  INV_X1    g0315(.A(G303), .ZN(new_n516));
  OAI22_X1  g0316(.A1(new_n377), .A2(new_n515), .B1(new_n516), .B2(new_n312), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n293), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n485), .A2(new_n513), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(G169), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n497), .B1(new_n512), .B2(new_n520), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n511), .A2(KEYINPUT21), .A3(G169), .A4(new_n519), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n519), .A2(new_n306), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n511), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n521), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n496), .A2(new_n526), .ZN(new_n527));
  AOI221_X4 g0327(.A(KEYINPUT24), .B1(new_n456), .B2(new_n461), .C1(new_n443), .C2(new_n447), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n465), .B1(new_n448), .B2(new_n462), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n253), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  AND2_X1   g0330(.A1(new_n492), .A2(new_n486), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n356), .B1(new_n531), .B2(new_n485), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n493), .A2(new_n302), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n530), .A2(new_n476), .A3(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(new_n535), .ZN(new_n536));
  OR2_X1    g0336(.A1(new_n519), .A2(new_n302), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n519), .A2(G200), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n512), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  NOR3_X1   g0340(.A1(new_n527), .A2(new_n536), .A3(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT90), .ZN(new_n542));
  OR2_X1    g0342(.A1(G238), .A2(G1698), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n543), .B1(G244), .B2(new_n314), .ZN(new_n544));
  OAI22_X1  g0344(.A1(new_n377), .A2(new_n544), .B1(new_n269), .B2(new_n499), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n293), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n206), .A2(G45), .ZN(new_n547));
  INV_X1    g0347(.A(G250), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n549), .B(new_n281), .C1(G274), .C2(new_n547), .ZN(new_n550));
  AND2_X1   g0350(.A1(new_n546), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n542), .B1(new_n551), .B2(G190), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n546), .A2(new_n550), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(G200), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n554), .B1(new_n302), .B2(new_n553), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n552), .B1(new_n555), .B2(new_n542), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n469), .A2(new_n440), .ZN(new_n557));
  XNOR2_X1  g0357(.A(new_n557), .B(KEYINPUT89), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT86), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT19), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n560), .A2(new_n207), .A3(G33), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n561), .B1(new_n503), .B2(new_n504), .ZN(new_n562));
  NOR2_X1   g0362(.A1(G87), .A2(G107), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n503), .A2(new_n504), .A3(new_n563), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n207), .B1(new_n269), .B2(new_n202), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n562), .B1(new_n566), .B2(KEYINPUT19), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n437), .A2(new_n266), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n559), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n560), .B1(new_n564), .B2(new_n565), .ZN(new_n570));
  OAI221_X1 g0370(.A(KEYINPUT86), .B1(new_n266), .B2(new_n437), .C1(new_n570), .C2(new_n562), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n569), .A2(new_n571), .A3(new_n253), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n326), .A2(new_n259), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(KEYINPUT87), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT87), .ZN(new_n576));
  OAI22_X1  g0376(.A1(new_n570), .A2(new_n562), .B1(new_n266), .B2(new_n437), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n258), .B1(new_n577), .B2(new_n559), .ZN(new_n578));
  AOI211_X1 g0378(.A(new_n576), .B(new_n573), .C1(new_n578), .C2(new_n571), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n556), .B(new_n558), .C1(new_n575), .C2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n470), .A2(new_n326), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n582), .B1(new_n579), .B2(new_n575), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(KEYINPUT88), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT88), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n585), .B(new_n582), .C1(new_n579), .C2(new_n575), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n551), .A2(new_n306), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n553), .A2(new_n421), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n581), .B1(new_n587), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n314), .A2(G244), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT4), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n312), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n502), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n548), .A2(new_n314), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n312), .A2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT84), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n312), .A2(KEYINPUT84), .A3(new_n598), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n597), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n594), .B1(new_n377), .B2(new_n593), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n281), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  OAI211_X1 g0405(.A(G257), .B(new_n281), .C1(new_n482), .C2(new_n484), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n485), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n421), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n601), .A2(new_n602), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n609), .A2(new_n596), .A3(new_n502), .ZN(new_n610));
  INV_X1    g0410(.A(new_n604), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n293), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n607), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n612), .A2(new_n613), .A3(new_n306), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n203), .B1(new_n399), .B2(new_n400), .ZN(new_n615));
  XNOR2_X1  g0415(.A(new_n615), .B(KEYINPUT83), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n273), .A2(new_n330), .ZN(new_n617));
  NAND2_X1  g0417(.A1(G97), .A2(G107), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n204), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(KEYINPUT6), .B1(new_n619), .B2(KEYINPUT82), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT82), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n204), .A2(new_n621), .A3(new_n618), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n505), .A2(KEYINPUT6), .A3(new_n203), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n617), .B1(new_n625), .B2(G20), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n258), .B1(new_n616), .B2(new_n626), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n259), .A2(G97), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n628), .B1(new_n470), .B2(G97), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n608), .B(new_n614), .C1(new_n627), .C2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT83), .ZN(new_n632));
  OR2_X1    g0432(.A1(new_n615), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n615), .A2(new_n632), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n626), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(new_n253), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n612), .A2(new_n613), .A3(G190), .ZN(new_n637));
  OAI21_X1  g0437(.A(G200), .B1(new_n605), .B2(new_n607), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n636), .A2(new_n629), .A3(new_n637), .A4(new_n638), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n631), .A2(new_n639), .ZN(new_n640));
  AOI21_X1  g0440(.A(KEYINPUT91), .B1(new_n592), .B2(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n590), .B1(new_n584), .B2(new_n586), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT91), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n631), .A2(new_n639), .ZN(new_n644));
  NOR4_X1   g0444(.A1(new_n642), .A2(new_n581), .A3(new_n643), .A4(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n541), .B1(new_n641), .B2(new_n645), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n435), .A2(new_n646), .ZN(G372));
  NOR2_X1   g0447(.A1(new_n279), .A2(new_n303), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n309), .B1(new_n648), .B2(new_n333), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n649), .A2(new_n417), .A3(new_n432), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n429), .A2(new_n423), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n364), .B1(new_n652), .B2(new_n361), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT97), .ZN(new_n654));
  INV_X1    g0454(.A(new_n555), .ZN(new_n655));
  OAI211_X1 g0455(.A(new_n655), .B(new_n558), .C1(new_n579), .C2(new_n575), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  OR2_X1    g0457(.A1(new_n589), .A2(KEYINPUT96), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n589), .A2(KEYINPUT96), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n658), .A2(new_n588), .A3(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n657), .B1(new_n587), .B2(new_n661), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n535), .A2(new_n631), .A3(new_n639), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n654), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n660), .B1(new_n584), .B2(new_n586), .ZN(new_n666));
  NOR4_X1   g0466(.A1(new_n666), .A2(KEYINPUT97), .A3(new_n663), .A4(new_n657), .ZN(new_n667));
  INV_X1    g0467(.A(new_n527), .ZN(new_n668));
  NOR3_X1   g0468(.A1(new_n665), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT26), .ZN(new_n670));
  INV_X1    g0470(.A(new_n631), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n662), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n587), .A2(new_n661), .ZN(new_n673));
  NOR3_X1   g0473(.A1(new_n642), .A2(new_n581), .A3(new_n631), .ZN(new_n674));
  OAI211_X1 g0474(.A(new_n672), .B(new_n673), .C1(new_n670), .C2(new_n674), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n669), .A2(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n653), .B1(new_n435), .B2(new_n676), .ZN(G369));
  NAND3_X1  g0477(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n678), .A2(KEYINPUT27), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(KEYINPUT27), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n679), .A2(G213), .A3(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(G343), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n512), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g0485(.A(new_n525), .B(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(new_n539), .ZN(new_n687));
  INV_X1    g0487(.A(G330), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n496), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n683), .B1(new_n467), .B2(new_n477), .ZN(new_n691));
  OR2_X1    g0491(.A1(new_n691), .A2(KEYINPUT98), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n536), .B1(KEYINPUT98), .B2(new_n691), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n690), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n496), .A2(new_n683), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n689), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n693), .A2(new_n692), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(new_n496), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n526), .A2(new_n683), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n695), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n697), .A2(new_n701), .ZN(G399));
  INV_X1    g0502(.A(new_n210), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(G41), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(G1), .ZN(new_n706));
  OR2_X1    g0506(.A1(new_n564), .A2(G116), .ZN(new_n707));
  OAI22_X1  g0507(.A1(new_n706), .A2(new_n707), .B1(new_n216), .B2(new_n705), .ZN(new_n708));
  XNOR2_X1  g0508(.A(new_n708), .B(KEYINPUT99), .ZN(new_n709));
  XNOR2_X1  g0509(.A(new_n709), .B(KEYINPUT28), .ZN(new_n710));
  OAI211_X1 g0510(.A(new_n541), .B(new_n684), .C1(new_n641), .C2(new_n645), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n605), .A2(new_n607), .ZN(new_n712));
  NOR3_X1   g0512(.A1(new_n712), .A2(G179), .A3(new_n551), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n713), .A2(new_n493), .A3(new_n519), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n712), .A2(new_n523), .A3(new_n551), .A4(new_n531), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT30), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n714), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n715), .A2(new_n716), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n683), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  XNOR2_X1  g0520(.A(new_n720), .B(KEYINPUT31), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n688), .B1(new_n711), .B2(new_n721), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n673), .A2(KEYINPUT26), .A3(new_n671), .A4(new_n656), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n723), .B1(new_n674), .B2(KEYINPUT26), .ZN(new_n724));
  NOR3_X1   g0524(.A1(new_n666), .A2(new_n657), .A3(new_n663), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n666), .B1(new_n725), .B2(new_n527), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n683), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT101), .ZN(new_n728));
  AND3_X1   g0528(.A1(new_n727), .A2(new_n728), .A3(KEYINPUT29), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n728), .B1(new_n727), .B2(KEYINPUT29), .ZN(new_n730));
  OR2_X1    g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n684), .B1(new_n669), .B2(new_n675), .ZN(new_n732));
  XNOR2_X1  g0532(.A(KEYINPUT100), .B(KEYINPUT29), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n722), .B1(new_n731), .B2(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n710), .B1(new_n735), .B2(G1), .ZN(G364));
  NOR2_X1   g0536(.A1(new_n254), .A2(G20), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n206), .B1(new_n737), .B2(G45), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n705), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n689), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n687), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n741), .B1(G330), .B2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(G13), .A2(G33), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(G20), .ZN(new_n746));
  AND2_X1   g0546(.A1(new_n687), .A2(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n213), .B1(G20), .B2(new_n421), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(G179), .A2(G200), .ZN(new_n750));
  XNOR2_X1  g0550(.A(new_n750), .B(KEYINPUT103), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n207), .B1(new_n751), .B2(G190), .ZN(new_n752));
  OR2_X1    g0552(.A1(new_n752), .A2(KEYINPUT104), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(KEYINPUT104), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G97), .ZN(new_n757));
  NOR4_X1   g0557(.A1(new_n207), .A2(new_n302), .A3(new_n356), .A4(G179), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR4_X1   g0559(.A1(new_n207), .A2(new_n356), .A3(G179), .A4(G190), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  OAI22_X1  g0561(.A1(new_n759), .A2(new_n440), .B1(new_n761), .B2(new_n203), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n207), .A2(G190), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n763), .A2(G179), .A3(new_n356), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n207), .A2(new_n306), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n765), .A2(G190), .A3(new_n356), .ZN(new_n766));
  OAI221_X1 g0566(.A(new_n312), .B1(new_n764), .B2(new_n330), .C1(new_n766), .C2(new_n388), .ZN(new_n767));
  NOR3_X1   g0567(.A1(new_n207), .A2(new_n306), .A3(new_n356), .ZN(new_n768));
  OR2_X1    g0568(.A1(new_n768), .A2(KEYINPUT102), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(KEYINPUT102), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n769), .A2(G190), .A3(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  AOI211_X1 g0572(.A(new_n762), .B(new_n767), .C1(new_n772), .C2(G50), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n751), .A2(new_n763), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(G159), .ZN(new_n776));
  OR2_X1    g0576(.A1(new_n776), .A2(KEYINPUT32), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n769), .A2(new_n302), .A3(new_n770), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  AOI22_X1  g0579(.A1(KEYINPUT32), .A2(new_n776), .B1(new_n779), .B2(G68), .ZN(new_n780));
  NAND4_X1  g0580(.A1(new_n757), .A2(new_n773), .A3(new_n777), .A4(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(G322), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n291), .B1(new_n766), .B2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(G283), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n759), .A2(new_n516), .B1(new_n761), .B2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n764), .ZN(new_n786));
  AOI211_X1 g0586(.A(new_n783), .B(new_n785), .C1(G311), .C2(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n775), .A2(G329), .ZN(new_n788));
  XNOR2_X1  g0588(.A(KEYINPUT33), .B(G317), .ZN(new_n789));
  AOI22_X1  g0589(.A1(G326), .A2(new_n772), .B1(new_n779), .B2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n752), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(G294), .ZN(new_n792));
  NAND4_X1  g0592(.A1(new_n787), .A2(new_n788), .A3(new_n790), .A4(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n749), .B1(new_n781), .B2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n703), .A2(new_n291), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G355), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n796), .B1(G116), .B2(new_n210), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n247), .A2(G45), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n210), .A2(new_n377), .ZN(new_n799));
  INV_X1    g0599(.A(G45), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n799), .B1(new_n800), .B2(new_n217), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n797), .B1(new_n798), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n746), .A2(new_n748), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n740), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  OR3_X1    g0605(.A1(new_n747), .A2(new_n794), .A3(new_n805), .ZN(new_n806));
  AND2_X1   g0606(.A1(new_n743), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(G396));
  NAND2_X1  g0608(.A1(new_n332), .A2(new_n683), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n337), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n323), .A2(new_n332), .A3(new_n683), .ZN(new_n811));
  AND2_X1   g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n732), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n337), .A2(new_n684), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n815), .B1(new_n669), .B2(new_n675), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n722), .B1(new_n813), .B2(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n817), .A2(new_n740), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n813), .A2(new_n722), .A3(new_n816), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n748), .A2(new_n744), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n740), .B1(G77), .B2(new_n822), .ZN(new_n823));
  OAI22_X1  g0623(.A1(new_n759), .A2(new_n203), .B1(new_n761), .B2(new_n440), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n291), .B1(new_n764), .B2(new_n499), .C1(new_n766), .C2(new_n490), .ZN(new_n825));
  AOI211_X1 g0625(.A(new_n824), .B(new_n825), .C1(G311), .C2(new_n775), .ZN(new_n826));
  AOI22_X1  g0626(.A1(G283), .A2(new_n779), .B1(new_n772), .B2(G303), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n757), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n766), .ZN(new_n829));
  AOI22_X1  g0629(.A1(G143), .A2(new_n829), .B1(new_n786), .B2(G159), .ZN(new_n830));
  INV_X1    g0630(.A(G137), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n830), .B1(new_n771), .B2(new_n831), .C1(new_n340), .C2(new_n778), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT34), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n377), .B1(new_n775), .B2(G132), .ZN(new_n835));
  OR2_X1    g0635(.A1(new_n835), .A2(KEYINPUT105), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(KEYINPUT105), .ZN(new_n837));
  OAI22_X1  g0637(.A1(new_n759), .A2(new_n272), .B1(new_n761), .B2(new_n266), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n838), .B1(new_n791), .B2(G58), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n834), .A2(new_n836), .A3(new_n837), .A4(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n832), .A2(new_n833), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n828), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n823), .B1(new_n842), .B2(new_n748), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n810), .A2(new_n811), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n843), .B1(new_n844), .B2(new_n745), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n820), .A2(new_n845), .ZN(G384));
  NOR2_X1   g0646(.A1(new_n215), .A2(new_n499), .ZN(new_n847));
  INV_X1    g0647(.A(new_n625), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT35), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n847), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n850), .B1(new_n849), .B2(new_n848), .ZN(new_n851));
  XNOR2_X1  g0651(.A(new_n851), .B(KEYINPUT36), .ZN(new_n852));
  OR3_X1    g0652(.A1(new_n389), .A2(new_n216), .A3(new_n330), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n272), .A2(G68), .ZN(new_n854));
  AOI211_X1 g0654(.A(new_n206), .B(G13), .C1(new_n853), .C2(new_n854), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n407), .A2(new_n408), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n387), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n858), .A2(new_n409), .A3(new_n253), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n681), .B1(new_n859), .B2(new_n386), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n433), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n405), .A2(new_n412), .ZN(new_n862));
  INV_X1    g0662(.A(new_n422), .ZN(new_n863));
  AOI22_X1  g0663(.A1(new_n863), .A2(new_n681), .B1(new_n859), .B2(new_n386), .ZN(new_n864));
  OAI21_X1  g0664(.A(KEYINPUT37), .B1(new_n862), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n681), .B1(new_n410), .B2(new_n386), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(KEYINPUT37), .B1(new_n418), .B2(new_n422), .ZN(new_n868));
  NAND4_X1  g0668(.A1(new_n867), .A2(new_n868), .A3(new_n405), .A4(new_n412), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n865), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n861), .A2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT38), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n861), .A2(KEYINPUT38), .A3(new_n870), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n279), .A2(new_n683), .ZN(new_n876));
  AND3_X1   g0676(.A1(new_n304), .A2(new_n309), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n876), .B1(new_n304), .B2(new_n309), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n670), .B1(new_n592), .B2(new_n671), .ZN(new_n881));
  NOR4_X1   g0681(.A1(new_n666), .A2(KEYINPUT26), .A3(new_n631), .A4(new_n657), .ZN(new_n882));
  NOR3_X1   g0682(.A1(new_n881), .A2(new_n882), .A3(new_n666), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n673), .A2(new_n656), .A3(new_n664), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(KEYINPUT97), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n662), .A2(new_n654), .A3(new_n664), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n885), .A2(new_n527), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n814), .B1(new_n883), .B2(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n333), .A2(new_n683), .ZN(new_n889));
  OAI211_X1 g0689(.A(new_n875), .B(new_n880), .C1(new_n888), .C2(new_n889), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n429), .A2(new_n423), .A3(new_n681), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n890), .A2(KEYINPUT106), .A3(new_n891), .ZN(new_n892));
  OR2_X1    g0692(.A1(new_n309), .A2(new_n683), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n417), .A2(new_n432), .A3(new_n651), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(new_n866), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n427), .A2(new_n404), .ZN(new_n897));
  OAI21_X1  g0697(.A(KEYINPUT37), .B1(new_n897), .B2(new_n866), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n869), .ZN(new_n899));
  AOI21_X1  g0699(.A(KEYINPUT38), .B1(new_n896), .B2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT39), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n901), .A2(new_n902), .A3(new_n874), .ZN(new_n903));
  AOI221_X4 g0703(.A(new_n872), .B1(new_n869), .B2(new_n865), .C1(new_n433), .C2(new_n860), .ZN(new_n904));
  AOI21_X1  g0704(.A(KEYINPUT38), .B1(new_n861), .B2(new_n870), .ZN(new_n905));
  OAI21_X1  g0705(.A(KEYINPUT39), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT107), .ZN(new_n907));
  AND3_X1   g0707(.A1(new_n903), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n907), .B1(new_n903), .B2(new_n906), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n894), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  AND2_X1   g0710(.A1(new_n892), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(KEYINPUT106), .B1(new_n890), .B2(new_n891), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n435), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n915), .B(new_n734), .C1(new_n729), .C2(new_n730), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(new_n653), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n914), .B(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n711), .A2(new_n721), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n844), .B1(new_n877), .B2(new_n878), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n919), .A2(new_n921), .A3(new_n875), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT40), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n920), .B1(new_n711), .B2(new_n721), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n923), .B1(new_n901), .B2(new_n874), .ZN(new_n925));
  AOI22_X1  g0725(.A1(new_n922), .A2(new_n923), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AND3_X1   g0726(.A1(new_n926), .A2(new_n915), .A3(new_n919), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n926), .B1(new_n915), .B2(new_n919), .ZN(new_n928));
  OR3_X1    g0728(.A1(new_n927), .A2(new_n928), .A3(new_n688), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n918), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n930), .B1(new_n206), .B2(new_n737), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n918), .A2(new_n929), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n856), .B1(new_n931), .B2(new_n932), .ZN(G367));
  INV_X1    g0733(.A(new_n662), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n558), .B1(new_n579), .B2(new_n575), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(new_n683), .ZN(new_n936));
  MUX2_X1   g0736(.A(new_n673), .B(new_n934), .S(new_n936), .Z(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n746), .ZN(new_n938));
  AND3_X1   g0738(.A1(new_n237), .A2(new_n210), .A3(new_n377), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n803), .B1(new_n210), .B2(new_n325), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n740), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n756), .A2(G68), .ZN(new_n942));
  OAI22_X1  g0742(.A1(new_n759), .A2(new_n388), .B1(new_n761), .B2(new_n330), .ZN(new_n943));
  OAI221_X1 g0743(.A(new_n312), .B1(new_n764), .B2(new_n272), .C1(new_n766), .C2(new_n340), .ZN(new_n944));
  AOI211_X1 g0744(.A(new_n943), .B(new_n944), .C1(G137), .C2(new_n775), .ZN(new_n945));
  AOI22_X1  g0745(.A1(G143), .A2(new_n772), .B1(new_n779), .B2(G159), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n942), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT46), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n759), .B2(new_n499), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n758), .A2(KEYINPUT46), .A3(G116), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n949), .B(new_n950), .C1(new_n778), .C2(new_n490), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n951), .A2(KEYINPUT110), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n761), .A2(new_n506), .ZN(new_n953));
  OAI221_X1 g0753(.A(new_n377), .B1(new_n764), .B2(new_n784), .C1(new_n766), .C2(new_n516), .ZN(new_n954));
  AOI211_X1 g0754(.A(new_n953), .B(new_n954), .C1(G317), .C2(new_n775), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n951), .A2(KEYINPUT110), .ZN(new_n956));
  AOI22_X1  g0756(.A1(new_n772), .A2(G311), .B1(new_n791), .B2(G107), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n952), .A2(new_n955), .A3(new_n956), .A4(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n947), .A2(new_n958), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n959), .B(KEYINPUT111), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(KEYINPUT47), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n941), .B1(new_n961), .B2(new_n748), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n938), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n684), .B1(new_n636), .B2(new_n629), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n640), .A2(KEYINPUT108), .A3(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT108), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n644), .B2(new_n964), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n631), .A2(new_n684), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n696), .A2(new_n700), .A3(new_n972), .ZN(new_n973));
  OR2_X1    g0773(.A1(new_n973), .A2(KEYINPUT42), .ZN(new_n974));
  INV_X1    g0774(.A(new_n969), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n631), .B1(new_n975), .B2(new_n496), .ZN(new_n976));
  AOI22_X1  g0776(.A1(new_n973), .A2(KEYINPUT42), .B1(new_n684), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT43), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n937), .A2(new_n979), .ZN(new_n980));
  OR2_X1    g0780(.A1(new_n937), .A2(new_n979), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n978), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n974), .A2(new_n977), .A3(new_n979), .A4(new_n937), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n697), .A2(new_n971), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n985), .B1(new_n982), .B2(new_n983), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  XOR2_X1   g0790(.A(new_n738), .B(KEYINPUT109), .Z(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT45), .ZN(new_n993));
  INV_X1    g0793(.A(new_n700), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n694), .A2(new_n994), .B1(new_n496), .B2(new_n683), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n993), .B1(new_n995), .B2(new_n971), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n701), .A2(new_n972), .A3(KEYINPUT45), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT44), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n701), .B2(new_n972), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n995), .A2(new_n971), .A3(KEYINPUT44), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n697), .B1(new_n998), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n998), .A2(new_n1002), .A3(new_n697), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n696), .B(new_n994), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(new_n689), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n735), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n704), .B(KEYINPUT41), .Z(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n992), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n963), .B1(new_n990), .B2(new_n1012), .ZN(G387));
  OAI21_X1  g0813(.A(new_n377), .B1(new_n761), .B2(new_n499), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(G317), .A2(new_n829), .B1(new_n786), .B2(G303), .ZN(new_n1015));
  INV_X1    g0815(.A(G311), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n1015), .B1(new_n771), .B2(new_n782), .C1(new_n1016), .C2(new_n778), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT48), .ZN(new_n1018));
  OR2_X1    g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n791), .A2(G283), .B1(G294), .B2(new_n758), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1019), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  XOR2_X1   g0822(.A(new_n1022), .B(KEYINPUT49), .Z(new_n1023));
  AOI211_X1 g0823(.A(new_n1014), .B(new_n1023), .C1(G326), .C2(new_n775), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n756), .A2(new_n326), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n758), .A2(G77), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1026), .B1(new_n202), .B2(new_n761), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n377), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1028), .B1(new_n272), .B2(new_n766), .C1(new_n266), .C2(new_n764), .ZN(new_n1029));
  AOI211_X1 g0829(.A(new_n1027), .B(new_n1029), .C1(G150), .C2(new_n775), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(G159), .A2(new_n772), .B1(new_n779), .B2(new_n342), .ZN(new_n1031));
  AND3_X1   g0831(.A1(new_n1025), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n748), .B1(new_n1024), .B2(new_n1032), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n795), .A2(new_n707), .B1(new_n203), .B2(new_n703), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n242), .A2(G45), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n1035), .B(KEYINPUT112), .Z(new_n1036));
  AOI211_X1 g0836(.A(G45), .B(new_n707), .C1(G68), .C2(G77), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n328), .A2(G50), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT50), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n799), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT113), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1034), .B1(new_n1036), .B2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n739), .B1(new_n1042), .B2(new_n803), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1033), .A2(new_n1043), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n1044), .B(KEYINPUT114), .Z(new_n1045));
  INV_X1    g0845(.A(new_n696), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1045), .B1(new_n1046), .B2(new_n746), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n1008), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1047), .B1(new_n1048), .B2(new_n992), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n705), .B1(new_n735), .B2(new_n1048), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n735), .B2(new_n1048), .ZN(new_n1051));
  AND2_X1   g0851(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n1052), .ZN(G393));
  INV_X1    g0853(.A(new_n1005), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n1054), .A2(new_n1003), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n971), .A2(new_n746), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n803), .B1(new_n210), .B2(new_n506), .C1(new_n250), .C2(new_n799), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n740), .A2(new_n1057), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n772), .A2(G317), .B1(G311), .B2(new_n829), .ZN(new_n1059));
  XOR2_X1   g0859(.A(new_n1059), .B(KEYINPUT52), .Z(new_n1060));
  AOI21_X1  g0860(.A(new_n312), .B1(new_n786), .B2(G294), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n1061), .B1(new_n203), .B2(new_n761), .C1(new_n784), .C2(new_n759), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(G322), .B2(new_n775), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n779), .A2(G303), .B1(new_n791), .B2(G116), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1060), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(G159), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n771), .A2(new_n340), .B1(new_n1066), .B2(new_n766), .ZN(new_n1067));
  XOR2_X1   g0867(.A(new_n1067), .B(KEYINPUT51), .Z(new_n1068));
  OAI22_X1  g0868(.A1(new_n778), .A2(new_n272), .B1(new_n328), .B2(new_n764), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT115), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n756), .A2(G77), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n1028), .B1(new_n761), .B2(new_n440), .C1(new_n759), .C2(new_n266), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1072), .B1(G143), .B2(new_n775), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1070), .A2(new_n1071), .A3(new_n1073), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1065), .B1(new_n1068), .B2(new_n1074), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT116), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1058), .B1(new_n1076), .B2(new_n748), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n1055), .A2(new_n992), .B1(new_n1056), .B2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n735), .A2(new_n1055), .A3(new_n1048), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n704), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1055), .B1(new_n735), .B2(new_n1048), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1078), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(KEYINPUT117), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT117), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n1084), .B(new_n1078), .C1(new_n1080), .C2(new_n1081), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1083), .A2(new_n1085), .ZN(G390));
  AOI21_X1  g0886(.A(new_n894), .B1(new_n901), .B2(new_n874), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n889), .B1(new_n727), .B2(new_n844), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1087), .B1(new_n1088), .B2(new_n879), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n889), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n816), .A2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n894), .B1(new_n1091), .B2(new_n880), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n902), .B1(new_n873), .B2(new_n874), .ZN(new_n1093));
  NOR3_X1   g0893(.A1(new_n904), .A2(new_n900), .A3(KEYINPUT39), .ZN(new_n1094));
  OAI21_X1  g0894(.A(KEYINPUT107), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n903), .A2(new_n906), .A3(new_n907), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1089), .B1(new_n1092), .B2(new_n1097), .ZN(new_n1098));
  AND3_X1   g0898(.A1(new_n722), .A2(new_n844), .A3(new_n880), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n879), .B1(new_n816), .B2(new_n1090), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n1095), .B(new_n1096), .C1(new_n1101), .C2(new_n894), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n722), .A2(new_n844), .A3(new_n880), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1102), .A2(new_n1103), .A3(new_n1089), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n915), .A2(new_n722), .ZN(new_n1105));
  AND3_X1   g0905(.A1(new_n916), .A2(new_n1105), .A3(new_n653), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n880), .B1(new_n722), .B2(new_n844), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1091), .B1(new_n1099), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n722), .A2(new_n844), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(new_n879), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1110), .A2(new_n1103), .A3(new_n1088), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1108), .A2(new_n1111), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n1100), .A2(new_n1104), .A3(new_n1106), .A4(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1100), .A2(new_n1104), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1106), .A2(new_n1112), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n705), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1100), .A2(new_n992), .A3(new_n1104), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n739), .B1(new_n328), .B2(new_n821), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(KEYINPUT54), .B(G143), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n764), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(G132), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n312), .B1(new_n766), .B2(new_n1121), .ZN(new_n1122));
  AOI211_X1 g0922(.A(new_n1120), .B(new_n1122), .C1(G50), .C2(new_n760), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n772), .A2(G128), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1123), .B(new_n1124), .C1(new_n831), .C2(new_n778), .ZN(new_n1125));
  XOR2_X1   g0925(.A(KEYINPUT118), .B(KEYINPUT53), .Z(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  NOR3_X1   g0927(.A1(new_n759), .A2(new_n1127), .A3(new_n340), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1127), .B1(new_n759), .B2(new_n340), .ZN(new_n1129));
  INV_X1    g0929(.A(G125), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1129), .B1(new_n774), .B2(new_n1130), .ZN(new_n1131));
  NOR3_X1   g0931(.A1(new_n1125), .A2(new_n1128), .A3(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n756), .A2(G159), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n312), .B1(new_n786), .B2(new_n505), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n758), .A2(G87), .B1(new_n760), .B2(G68), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n1134), .B(new_n1135), .C1(new_n499), .C2(new_n766), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n203), .A2(new_n778), .B1(new_n771), .B2(new_n784), .ZN(new_n1137));
  AOI211_X1 g0937(.A(new_n1136), .B(new_n1137), .C1(G294), .C2(new_n775), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n1132), .A2(new_n1133), .B1(new_n1138), .B2(new_n1071), .ZN(new_n1139));
  OAI221_X1 g0939(.A(new_n1118), .B1(new_n749), .B2(new_n1139), .C1(new_n1097), .C2(new_n745), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1117), .A2(new_n1140), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n1113), .A2(new_n1116), .B1(new_n1141), .B2(KEYINPUT119), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT119), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1117), .A2(new_n1143), .A3(new_n1140), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT120), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1141), .A2(KEYINPUT119), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1104), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1103), .B1(new_n1102), .B2(new_n1089), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1115), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1151), .A2(new_n704), .A3(new_n1113), .ZN(new_n1152));
  AND4_X1   g0952(.A1(KEYINPUT120), .A2(new_n1148), .A3(new_n1152), .A4(new_n1144), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1147), .A2(new_n1154), .ZN(G378));
  NAND2_X1  g0955(.A1(new_n361), .A2(new_n365), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n347), .A2(new_n681), .ZN(new_n1157));
  XOR2_X1   g0957(.A(new_n1157), .B(KEYINPUT55), .Z(new_n1158));
  XNOR2_X1  g0958(.A(new_n1156), .B(new_n1158), .ZN(new_n1159));
  XOR2_X1   g0959(.A(KEYINPUT122), .B(KEYINPUT56), .Z(new_n1160));
  XNOR2_X1  g0960(.A(new_n1159), .B(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n926), .A2(G330), .A3(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n922), .A2(new_n923), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n924), .A2(new_n925), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1163), .A2(G330), .A3(new_n1164), .ZN(new_n1165));
  XOR2_X1   g0965(.A(new_n1159), .B(new_n1160), .Z(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n911), .A2(new_n913), .A3(new_n1162), .A4(new_n1167), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1161), .B1(new_n926), .B2(G330), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n892), .A2(new_n910), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n1169), .A2(new_n1170), .B1(new_n1171), .B2(new_n912), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1168), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(new_n992), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n740), .B1(G50), .B2(new_n822), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(G33), .A2(G41), .ZN(new_n1176));
  AOI211_X1 g0976(.A(G50), .B(new_n1176), .C1(new_n377), .C2(new_n479), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n778), .A2(new_n202), .B1(new_n325), .B2(new_n764), .ZN(new_n1178));
  XOR2_X1   g0978(.A(new_n1178), .B(KEYINPUT121), .Z(new_n1179));
  OAI211_X1 g0979(.A(new_n479), .B(new_n377), .C1(new_n774), .C2(new_n784), .ZN(new_n1180));
  OAI221_X1 g0980(.A(new_n1026), .B1(new_n203), .B2(new_n766), .C1(new_n388), .C2(new_n761), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n1180), .B(new_n1181), .C1(G116), .C2(new_n772), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1179), .A2(new_n942), .A3(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT58), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1177), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n771), .A2(new_n1130), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(G128), .A2(new_n829), .B1(new_n786), .B2(G137), .ZN(new_n1187));
  OAI221_X1 g0987(.A(new_n1187), .B1(new_n759), .B2(new_n1119), .C1(new_n778), .C2(new_n1121), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n1186), .B(new_n1188), .C1(G150), .C2(new_n756), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1190), .A2(KEYINPUT59), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1176), .B1(new_n761), .B2(new_n1066), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(G124), .B2(new_n775), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT59), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1193), .B1(new_n1189), .B2(new_n1194), .ZN(new_n1195));
  OAI221_X1 g0995(.A(new_n1185), .B1(new_n1184), .B2(new_n1183), .C1(new_n1191), .C2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1175), .B1(new_n1196), .B2(new_n748), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1197), .B1(new_n1161), .B2(new_n745), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1174), .A2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n1113), .A2(new_n1106), .B1(new_n1168), .B2(new_n1172), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n704), .B1(new_n1201), .B2(KEYINPUT57), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1113), .A2(new_n1106), .ZN(new_n1203));
  AND3_X1   g1003(.A1(new_n1203), .A2(KEYINPUT57), .A3(new_n1173), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1200), .B1(new_n1202), .B2(new_n1204), .ZN(G375));
  NAND2_X1  g1005(.A1(new_n879), .A2(new_n744), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n759), .A2(new_n202), .B1(new_n761), .B2(new_n330), .ZN(new_n1207));
  OAI221_X1 g1007(.A(new_n291), .B1(new_n764), .B2(new_n203), .C1(new_n766), .C2(new_n784), .ZN(new_n1208));
  AOI211_X1 g1008(.A(new_n1207), .B(new_n1208), .C1(G303), .C2(new_n775), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(G116), .A2(new_n779), .B1(new_n772), .B2(G294), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1025), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n759), .A2(new_n1066), .B1(new_n761), .B2(new_n388), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n1028), .B1(new_n831), .B2(new_n766), .C1(new_n340), .C2(new_n764), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n1212), .B(new_n1213), .C1(G128), .C2(new_n775), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1119), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(G132), .A2(new_n772), .B1(new_n779), .B2(new_n1215), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n1214), .B(new_n1216), .C1(new_n272), .C2(new_n755), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n749), .B1(new_n1211), .B2(new_n1217), .ZN(new_n1218));
  AOI211_X1 g1018(.A(new_n739), .B(new_n1218), .C1(new_n266), .C2(new_n821), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n1112), .A2(new_n992), .B1(new_n1206), .B2(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n916), .A2(new_n1105), .A3(new_n653), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1221), .A2(new_n1108), .A3(new_n1111), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1115), .A2(new_n1222), .ZN(new_n1223));
  XOR2_X1   g1023(.A(new_n1010), .B(KEYINPUT123), .Z(new_n1224));
  OAI21_X1  g1024(.A(new_n1220), .B1(new_n1223), .B2(new_n1224), .ZN(G381));
  NAND2_X1  g1025(.A1(new_n1203), .A2(new_n1173), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT57), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1201), .A2(KEYINPUT57), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1228), .A2(new_n704), .A3(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1141), .B1(new_n1116), .B2(new_n1113), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1230), .A2(new_n1200), .A3(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1012), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(new_n989), .ZN(new_n1234));
  NAND4_X1  g1034(.A1(new_n1083), .A2(new_n1234), .A3(new_n963), .A4(new_n1085), .ZN(new_n1235));
  AND3_X1   g1035(.A1(new_n1049), .A2(new_n807), .A3(new_n1051), .ZN(new_n1236));
  INV_X1    g1036(.A(G384), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  OR4_X1    g1038(.A1(G381), .A2(new_n1232), .A3(new_n1235), .A4(new_n1238), .ZN(G407));
  OAI211_X1 g1039(.A(G407), .B(G213), .C1(G343), .C2(new_n1232), .ZN(G409));
  INV_X1    g1040(.A(new_n1085), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n735), .A2(new_n1048), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(new_n1006), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1243), .A2(new_n704), .A3(new_n1079), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1084), .B1(new_n1244), .B2(new_n1078), .ZN(new_n1245));
  OAI21_X1  g1045(.A(G387), .B1(new_n1241), .B2(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n807), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1236), .A2(new_n1247), .ZN(new_n1248));
  AND3_X1   g1048(.A1(new_n1246), .A2(new_n1235), .A3(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1248), .B1(new_n1246), .B2(new_n1235), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  XOR2_X1   g1051(.A(KEYINPUT127), .B(KEYINPUT61), .Z(new_n1252));
  NAND2_X1  g1052(.A1(new_n682), .A2(G213), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1254), .A2(G2897), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT60), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1222), .A2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(new_n704), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1257), .B1(new_n1115), .B2(new_n1222), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1220), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(new_n1237), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT124), .ZN(new_n1263));
  OAI211_X1 g1063(.A(G384), .B(new_n1220), .C1(new_n1259), .C2(new_n1260), .ZN(new_n1264));
  AND3_X1   g1064(.A1(new_n1262), .A2(new_n1263), .A3(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1263), .B1(new_n1262), .B2(new_n1264), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1256), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1223), .A2(KEYINPUT60), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n705), .B1(new_n1222), .B2(new_n1257), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(G384), .B1(new_n1270), .B2(new_n1220), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1264), .ZN(new_n1272));
  OAI21_X1  g1072(.A(KEYINPUT124), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(new_n1255), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1267), .A2(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(KEYINPUT120), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1276));
  OAI211_X1 g1076(.A(new_n1200), .B(new_n1230), .C1(new_n1276), .C2(new_n1153), .ZN(new_n1277));
  OR2_X1    g1077(.A1(new_n1226), .A2(new_n1224), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1278), .A2(new_n1200), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(new_n1231), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1254), .B1(new_n1277), .B2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1262), .A2(new_n1264), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  AOI21_X1  g1083(.A(G375), .B1(new_n1147), .B2(new_n1154), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1231), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1285), .B1(new_n1278), .B2(new_n1200), .ZN(new_n1286));
  OAI211_X1 g1086(.A(new_n1253), .B(new_n1283), .C1(new_n1284), .C2(new_n1286), .ZN(new_n1287));
  OAI221_X1 g1087(.A(new_n1252), .B1(new_n1275), .B2(new_n1281), .C1(new_n1287), .C2(KEYINPUT62), .ZN(new_n1288));
  AND2_X1   g1088(.A1(new_n1287), .A2(KEYINPUT62), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1251), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT126), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT63), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1282), .A2(new_n1292), .ZN(new_n1293));
  OAI211_X1 g1093(.A(new_n1293), .B(new_n1253), .C1(new_n1284), .C2(new_n1286), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1250), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1246), .A2(new_n1235), .A3(new_n1248), .ZN(new_n1296));
  AOI21_X1  g1096(.A(KEYINPUT61), .B1(new_n1295), .B2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1294), .A2(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(KEYINPUT63), .B1(new_n1281), .B2(new_n1283), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT125), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1262), .A2(new_n1263), .A3(new_n1264), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1255), .B1(new_n1273), .B2(new_n1302), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(new_n1266), .A2(new_n1256), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1301), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1253), .B1(new_n1284), .B2(new_n1286), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1267), .A2(KEYINPUT125), .A3(new_n1274), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1305), .A2(new_n1306), .A3(new_n1307), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1291), .B1(new_n1300), .B2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT61), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1310), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1311), .B1(new_n1281), .B2(new_n1293), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1287), .A2(new_n1292), .ZN(new_n1313));
  AND4_X1   g1113(.A1(new_n1291), .A2(new_n1308), .A3(new_n1312), .A4(new_n1313), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1290), .B1(new_n1309), .B2(new_n1314), .ZN(G405));
  AOI21_X1  g1115(.A(new_n1284), .B1(G375), .B2(new_n1231), .ZN(new_n1316));
  OR2_X1    g1116(.A1(new_n1316), .A2(new_n1282), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1316), .A2(new_n1282), .ZN(new_n1318));
  AND3_X1   g1118(.A1(new_n1317), .A2(new_n1251), .A3(new_n1318), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1251), .B1(new_n1317), .B2(new_n1318), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(new_n1319), .A2(new_n1320), .ZN(G402));
endmodule


