//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 0 0 0 0 1 0 0 1 1 0 1 0 0 1 1 0 0 1 1 1 0 0 0 0 0 0 1 0 1 1 0 1 1 1 1 1 1 1 1 0 1 0 0 0 1 0 0 0 0 0 0 0 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:13 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n661,
    new_n662, new_n663, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974;
  INV_X1    g000(.A(KEYINPUT82), .ZN(new_n187));
  INV_X1    g001(.A(G217), .ZN(new_n188));
  INV_X1    g002(.A(G902), .ZN(new_n189));
  AOI21_X1  g003(.A(new_n188), .B1(G234), .B2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G128), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n192), .A2(G119), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT69), .B(G128), .ZN(new_n194));
  AOI21_X1  g008(.A(new_n193), .B1(new_n194), .B2(G119), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT23), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT23), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n197), .A2(new_n192), .A3(G119), .ZN(new_n198));
  AND2_X1   g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G110), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT76), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G140), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G125), .ZN(new_n204));
  OR2_X1    g018(.A1(new_n204), .A2(KEYINPUT16), .ZN(new_n205));
  INV_X1    g019(.A(G125), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G140), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n204), .A2(new_n207), .A3(KEYINPUT16), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n205), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n205), .A2(G146), .A3(new_n208), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n199), .A2(KEYINPUT76), .A3(G110), .ZN(new_n214));
  XOR2_X1   g028(.A(KEYINPUT24), .B(G110), .Z(new_n215));
  NAND2_X1  g029(.A1(new_n195), .A2(new_n215), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n202), .A2(new_n213), .A3(new_n214), .A4(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n204), .A2(new_n207), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n218), .A2(G146), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  AOI21_X1  g034(.A(G110), .B1(new_n196), .B2(new_n198), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n195), .A2(new_n215), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n212), .B(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT77), .ZN(new_n224));
  OR2_X1    g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n223), .A2(new_n224), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n217), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G953), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n228), .A2(G221), .A3(G234), .ZN(new_n229));
  XNOR2_X1  g043(.A(new_n229), .B(KEYINPUT22), .ZN(new_n230));
  XNOR2_X1  g044(.A(new_n230), .B(G137), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n227), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT78), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n227), .A2(new_n234), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n217), .A2(new_n225), .A3(KEYINPUT78), .A4(new_n226), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n233), .B1(new_n237), .B2(new_n232), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(new_n189), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT25), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n238), .A2(KEYINPUT25), .A3(new_n189), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n191), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n190), .A2(G902), .ZN(new_n244));
  XNOR2_X1  g058(.A(KEYINPUT80), .B(KEYINPUT81), .ZN(new_n245));
  XNOR2_X1  g059(.A(new_n244), .B(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  OR2_X1    g061(.A1(new_n238), .A2(KEYINPUT79), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n238), .A2(KEYINPUT79), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n247), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n187), .B1(new_n243), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n242), .ZN(new_n252));
  AOI21_X1  g066(.A(KEYINPUT25), .B1(new_n238), .B2(new_n189), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n190), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n249), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n238), .A2(KEYINPUT79), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n246), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n254), .A2(KEYINPUT82), .A3(new_n257), .ZN(new_n258));
  AND2_X1   g072(.A1(new_n251), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(G237), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n260), .A2(new_n228), .A3(G210), .ZN(new_n261));
  XOR2_X1   g075(.A(new_n261), .B(KEYINPUT27), .Z(new_n262));
  XNOR2_X1  g076(.A(new_n262), .B(KEYINPUT26), .ZN(new_n263));
  XOR2_X1   g077(.A(new_n263), .B(G101), .Z(new_n264));
  NAND3_X1  g078(.A1(new_n210), .A2(KEYINPUT65), .A3(G143), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n192), .A2(KEYINPUT1), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT65), .ZN(new_n267));
  INV_X1    g081(.A(G143), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n267), .B1(new_n268), .B2(G146), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n268), .A2(G146), .ZN(new_n270));
  OAI211_X1 g084(.A(new_n265), .B(new_n266), .C1(new_n269), .C2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT68), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n210), .A2(G143), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n210), .A2(G143), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n274), .B1(new_n275), .B2(new_n267), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n276), .A2(KEYINPUT68), .A3(new_n265), .A4(new_n266), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n273), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n194), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n274), .A2(KEYINPUT1), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n268), .A2(G146), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n274), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n278), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(G137), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(G134), .ZN(new_n287));
  INV_X1    g101(.A(G134), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(G137), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(G131), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT11), .ZN(new_n292));
  OAI22_X1  g106(.A1(KEYINPUT66), .A2(new_n292), .B1(new_n288), .B2(G137), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT66), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n294), .A2(new_n286), .A3(KEYINPUT11), .A4(G134), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n292), .A2(KEYINPUT66), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n293), .A2(new_n295), .A3(new_n296), .A4(new_n289), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n291), .B1(new_n297), .B2(G131), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n285), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(KEYINPUT0), .A2(G128), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  OAI211_X1 g116(.A(new_n265), .B(new_n302), .C1(new_n269), .C2(new_n270), .ZN(new_n303));
  OR2_X1    g117(.A1(KEYINPUT0), .A2(G128), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n283), .A2(new_n301), .A3(new_n304), .ZN(new_n305));
  AND2_X1   g119(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  AND2_X1   g120(.A1(new_n297), .A2(G131), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n297), .A2(G131), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n306), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  AND2_X1   g123(.A1(new_n300), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(G116), .ZN(new_n311));
  OR3_X1    g125(.A1(new_n311), .A2(KEYINPUT70), .A3(G119), .ZN(new_n312));
  AOI21_X1  g126(.A(KEYINPUT70), .B1(new_n311), .B2(G119), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n311), .A2(G119), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n312), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  XNOR2_X1  g129(.A(KEYINPUT2), .B(G113), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n315), .B(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n310), .A2(new_n318), .ZN(new_n319));
  XNOR2_X1  g133(.A(new_n319), .B(KEYINPUT28), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT67), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n309), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n297), .B(G131), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n323), .A2(KEYINPUT67), .A3(new_n306), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n300), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(new_n317), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n264), .B1(new_n320), .B2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  AOI22_X1  g142(.A1(new_n273), .A2(new_n277), .B1(new_n283), .B2(new_n281), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n309), .B(KEYINPUT30), .C1(new_n329), .C2(new_n298), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT71), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n300), .A2(KEYINPUT71), .A3(KEYINPUT30), .A4(new_n309), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  XNOR2_X1  g148(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n325), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n334), .A2(new_n317), .A3(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT72), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  AOI22_X1  g153(.A1(new_n332), .A2(new_n333), .B1(new_n325), .B2(new_n335), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n340), .A2(KEYINPUT72), .A3(new_n317), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n264), .A2(new_n319), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(KEYINPUT31), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT31), .ZN(new_n346));
  AOI211_X1 g160(.A(new_n346), .B(new_n343), .C1(new_n339), .C2(new_n341), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n328), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(KEYINPUT73), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT73), .ZN(new_n350));
  OAI211_X1 g164(.A(new_n350), .B(new_n328), .C1(new_n345), .C2(new_n347), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  NOR2_X1   g166(.A1(G472), .A2(G902), .ZN(new_n353));
  XNOR2_X1  g167(.A(new_n353), .B(KEYINPUT74), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  AOI21_X1  g169(.A(KEYINPUT32), .B1(new_n352), .B2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT32), .ZN(new_n357));
  AOI211_X1 g171(.A(new_n357), .B(new_n354), .C1(new_n349), .C2(new_n351), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(new_n319), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n360), .B1(new_n339), .B2(new_n341), .ZN(new_n361));
  OR2_X1    g175(.A1(new_n361), .A2(new_n264), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT29), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT75), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n320), .A2(new_n364), .A3(new_n326), .A4(new_n264), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n320), .A2(new_n326), .A3(new_n264), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(KEYINPUT75), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n362), .A2(new_n363), .A3(new_n365), .A4(new_n367), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n310), .A2(new_n318), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n320), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n264), .A2(KEYINPUT29), .ZN(new_n372));
  OAI211_X1 g186(.A(new_n368), .B(new_n189), .C1(new_n371), .C2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(G472), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n259), .B1(new_n359), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(G104), .ZN(new_n376));
  OAI21_X1  g190(.A(KEYINPUT3), .B1(new_n376), .B2(G107), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT3), .ZN(new_n378));
  INV_X1    g192(.A(G107), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n378), .A2(new_n379), .A3(G104), .ZN(new_n380));
  OAI211_X1 g194(.A(new_n377), .B(new_n380), .C1(G104), .C2(new_n379), .ZN(new_n381));
  OR2_X1    g195(.A1(new_n381), .A2(G101), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n376), .A2(G107), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n379), .A2(G104), .ZN(new_n384));
  OAI21_X1  g198(.A(G101), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  AND2_X1   g199(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  OR2_X1    g200(.A1(new_n315), .A2(new_n316), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT5), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n314), .A2(new_n388), .ZN(new_n389));
  OAI211_X1 g203(.A(G113), .B(new_n389), .C1(new_n315), .C2(new_n388), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n386), .A2(new_n387), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n381), .A2(G101), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n382), .A2(KEYINPUT4), .A3(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT4), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n381), .A2(new_n394), .A3(G101), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n393), .A2(new_n317), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n391), .A2(new_n396), .ZN(new_n397));
  XOR2_X1   g211(.A(G110), .B(G122), .Z(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n398), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n391), .A2(new_n396), .A3(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n399), .A2(KEYINPUT6), .A3(new_n401), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n306), .A2(new_n206), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n403), .B1(new_n206), .B2(new_n329), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n228), .A2(G224), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n404), .B(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT6), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n397), .A2(new_n407), .A3(new_n398), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n402), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n404), .A2(KEYINPUT7), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n404), .A2(new_n405), .ZN(new_n411));
  XOR2_X1   g225(.A(KEYINPUT84), .B(KEYINPUT8), .Z(new_n412));
  XNOR2_X1  g226(.A(new_n398), .B(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n390), .A2(new_n387), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n382), .A2(new_n385), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n413), .B1(new_n391), .B2(new_n416), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n411), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n404), .A2(KEYINPUT7), .A3(new_n405), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n418), .A2(new_n419), .A3(new_n401), .ZN(new_n420));
  OAI211_X1 g234(.A(new_n409), .B(new_n189), .C1(new_n410), .C2(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(G210), .B1(G237), .B2(G902), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  OR2_X1    g237(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n421), .A2(new_n423), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(G214), .B1(G237), .B2(G902), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n260), .A2(new_n228), .A3(G214), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n429), .B(G143), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT18), .ZN(new_n431));
  INV_X1    g245(.A(G131), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n430), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n430), .A2(new_n432), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(KEYINPUT18), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT85), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n218), .B(new_n436), .ZN(new_n437));
  AND2_X1   g251(.A1(new_n437), .A2(G146), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n433), .B(new_n435), .C1(new_n438), .C2(new_n219), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n437), .A2(KEYINPUT19), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n440), .B1(KEYINPUT19), .B2(new_n218), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n441), .A2(G146), .ZN(new_n442));
  AND2_X1   g256(.A1(new_n430), .A2(new_n432), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n212), .B1(new_n443), .B2(new_n434), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n439), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  XOR2_X1   g259(.A(G113), .B(G122), .Z(new_n446));
  XNOR2_X1  g260(.A(new_n446), .B(KEYINPUT86), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n447), .B(new_n376), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  OR3_X1    g263(.A1(new_n443), .A2(new_n434), .A3(KEYINPUT17), .ZN(new_n450));
  OR2_X1    g264(.A1(new_n213), .A2(KEYINPUT87), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n434), .A2(KEYINPUT17), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n213), .A2(KEYINPUT87), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n450), .A2(new_n451), .A3(new_n452), .A4(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n448), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n454), .A2(new_n439), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n449), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(G475), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n457), .A2(new_n458), .A3(new_n189), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(KEYINPUT20), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT88), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n459), .A2(KEYINPUT88), .A3(KEYINPUT20), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT20), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n457), .A2(new_n464), .A3(new_n458), .A4(new_n189), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(KEYINPUT89), .ZN(new_n466));
  AOI21_X1  g280(.A(G475), .B1(new_n449), .B2(new_n456), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT89), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n467), .A2(new_n468), .A3(new_n464), .A4(new_n189), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n462), .A2(new_n463), .A3(new_n466), .A4(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n454), .A2(new_n439), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(new_n448), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(new_n456), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n458), .B1(new_n473), .B2(new_n189), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n470), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(G234), .A2(G237), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n477), .A2(G952), .A3(new_n228), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  XOR2_X1   g293(.A(KEYINPUT21), .B(G898), .Z(new_n480));
  XNOR2_X1  g294(.A(new_n480), .B(KEYINPUT92), .ZN(new_n481));
  AND3_X1   g295(.A1(new_n477), .A2(G902), .A3(G953), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n479), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(G122), .ZN(new_n484));
  OAI21_X1  g298(.A(KEYINPUT14), .B1(new_n484), .B2(G116), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n485), .B1(new_n311), .B2(G122), .ZN(new_n486));
  NOR3_X1   g300(.A1(new_n484), .A2(KEYINPUT14), .A3(G116), .ZN(new_n487));
  OAI21_X1  g301(.A(G107), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT91), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n488), .B(new_n489), .ZN(new_n490));
  XNOR2_X1  g304(.A(G116), .B(G122), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(new_n379), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT90), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n493), .B1(new_n279), .B2(new_n268), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n194), .A2(KEYINPUT90), .A3(G143), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n192), .A2(G143), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n288), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  AOI211_X1 g313(.A(G134), .B(new_n497), .C1(new_n494), .C2(new_n495), .ZN(new_n500));
  OAI211_X1 g314(.A(new_n490), .B(new_n492), .C1(new_n499), .C2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n496), .A2(new_n288), .A3(new_n498), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n491), .B(new_n379), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n497), .B(KEYINPUT13), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n504), .B1(new_n494), .B2(new_n495), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n502), .B(new_n503), .C1(new_n288), .C2(new_n505), .ZN(new_n506));
  XOR2_X1   g320(.A(KEYINPUT9), .B(G234), .Z(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  NOR3_X1   g322(.A1(new_n508), .A2(new_n188), .A3(G953), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  AND3_X1   g324(.A1(new_n501), .A2(new_n506), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n510), .B1(new_n501), .B2(new_n506), .ZN(new_n512));
  NOR3_X1   g326(.A1(new_n511), .A2(new_n512), .A3(G902), .ZN(new_n513));
  INV_X1    g327(.A(G478), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n514), .A2(KEYINPUT15), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n513), .B(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  NOR4_X1   g331(.A1(new_n428), .A2(new_n476), .A3(new_n483), .A4(new_n517), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n285), .A2(new_n386), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n276), .A2(new_n265), .ZN(new_n520));
  INV_X1    g334(.A(new_n280), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n520), .B1(new_n192), .B2(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n415), .B1(new_n278), .B2(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n323), .B1(new_n519), .B2(new_n523), .ZN(new_n524));
  XOR2_X1   g338(.A(new_n524), .B(KEYINPUT12), .Z(new_n525));
  OR2_X1    g339(.A1(new_n523), .A2(KEYINPUT10), .ZN(new_n526));
  INV_X1    g340(.A(new_n323), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n393), .A2(new_n306), .A3(new_n395), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n285), .A2(new_n386), .A3(KEYINPUT10), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n526), .A2(new_n527), .A3(new_n528), .A4(new_n529), .ZN(new_n530));
  XOR2_X1   g344(.A(G110), .B(G140), .Z(new_n531));
  XNOR2_X1  g345(.A(new_n531), .B(KEYINPUT83), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n228), .A2(G227), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n532), .B(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  AND2_X1   g349(.A1(new_n530), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n525), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n526), .A2(new_n528), .A3(new_n529), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(new_n323), .ZN(new_n539));
  AND2_X1   g353(.A1(new_n539), .A2(new_n530), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n537), .B1(new_n540), .B2(new_n535), .ZN(new_n541));
  INV_X1    g355(.A(G469), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n541), .A2(new_n542), .A3(new_n189), .ZN(new_n543));
  NAND2_X1  g357(.A1(G469), .A2(G902), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n536), .A2(new_n539), .ZN(new_n545));
  AND2_X1   g359(.A1(new_n525), .A2(new_n530), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n545), .B1(new_n546), .B2(new_n535), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n543), .B(new_n544), .C1(new_n542), .C2(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(G221), .B1(new_n508), .B2(G902), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  AND2_X1   g365(.A1(new_n518), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n375), .A2(new_n552), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n553), .B(G101), .ZN(G3));
  AOI21_X1  g368(.A(new_n354), .B1(new_n349), .B2(new_n351), .ZN(new_n555));
  AOI21_X1  g369(.A(KEYINPUT72), .B1(new_n340), .B2(new_n317), .ZN(new_n556));
  AND4_X1   g370(.A1(KEYINPUT72), .A2(new_n334), .A3(new_n317), .A4(new_n336), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n344), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(new_n346), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n342), .A2(KEYINPUT31), .A3(new_n344), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n350), .B1(new_n561), .B2(new_n328), .ZN(new_n562));
  AOI211_X1 g376(.A(KEYINPUT73), .B(new_n327), .C1(new_n559), .C2(new_n560), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n189), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n555), .B1(new_n564), .B2(G472), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n251), .A2(new_n258), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n565), .A2(new_n566), .A3(new_n551), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT93), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n428), .A2(new_n483), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n565), .A2(new_n566), .A3(KEYINPUT93), .A4(new_n551), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n511), .A2(new_n512), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT94), .ZN(new_n574));
  OR2_X1    g388(.A1(new_n509), .A2(KEYINPUT95), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n573), .A2(new_n574), .A3(KEYINPUT33), .A4(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n501), .A2(new_n506), .ZN(new_n577));
  OR2_X1    g391(.A1(new_n577), .A2(new_n575), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n509), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n501), .A2(new_n506), .A3(new_n510), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n579), .A2(new_n574), .A3(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT33), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n576), .A2(new_n578), .A3(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n584), .A2(G478), .A3(new_n189), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT97), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT96), .ZN(new_n587));
  OR3_X1    g401(.A1(new_n513), .A2(new_n587), .A3(G478), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n587), .B1(new_n513), .B2(G478), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  AND3_X1   g404(.A1(new_n585), .A2(new_n586), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n586), .B1(new_n585), .B2(new_n590), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AOI211_X1 g407(.A(new_n461), .B(new_n464), .C1(new_n467), .C2(new_n189), .ZN(new_n594));
  AOI21_X1  g408(.A(KEYINPUT88), .B1(new_n459), .B2(KEYINPUT20), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AND2_X1   g410(.A1(new_n466), .A2(new_n469), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n474), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n593), .A2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n572), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g415(.A(KEYINPUT34), .B(G104), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n601), .B(new_n602), .ZN(G6));
  AOI21_X1  g417(.A(new_n474), .B1(new_n596), .B2(new_n465), .ZN(new_n604));
  AND2_X1   g418(.A1(new_n604), .A2(new_n517), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n572), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(KEYINPUT35), .B(G107), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n607), .B(new_n608), .ZN(G9));
  NOR2_X1   g423(.A1(new_n232), .A2(KEYINPUT36), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(KEYINPUT98), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n237), .B(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n246), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n254), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n552), .A2(new_n565), .A3(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(KEYINPUT99), .ZN(new_n616));
  XNOR2_X1  g430(.A(KEYINPUT37), .B(G110), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G12));
  INV_X1    g432(.A(new_n614), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n619), .B1(new_n359), .B2(new_n374), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT102), .ZN(new_n621));
  XOR2_X1   g435(.A(new_n478), .B(KEYINPUT101), .Z(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(G900), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n477), .A2(new_n624), .A3(G902), .A4(G953), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(KEYINPUT100), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n604), .A2(new_n621), .A3(new_n517), .A4(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n462), .A2(new_n463), .A3(new_n465), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n629), .A2(new_n517), .A3(new_n475), .A4(new_n627), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(KEYINPUT102), .ZN(new_n631));
  INV_X1    g445(.A(new_n428), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n628), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  OR2_X1    g447(.A1(new_n633), .A2(KEYINPUT103), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(KEYINPUT103), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n620), .A2(new_n551), .A3(new_n634), .A4(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(KEYINPUT104), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(G128), .ZN(G30));
  XOR2_X1   g452(.A(new_n627), .B(KEYINPUT39), .Z(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n551), .A2(new_n640), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n619), .B1(new_n641), .B2(KEYINPUT40), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n642), .B1(KEYINPUT40), .B2(new_n641), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT38), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n426), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n424), .A2(KEYINPUT38), .A3(new_n425), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n427), .ZN(new_n648));
  NOR4_X1   g462(.A1(new_n647), .A2(new_n648), .A3(new_n516), .A4(new_n598), .ZN(new_n649));
  INV_X1    g463(.A(G472), .ZN(new_n650));
  INV_X1    g464(.A(new_n264), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n361), .A2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n360), .A2(new_n264), .ZN(new_n654));
  AOI21_X1  g468(.A(G902), .B1(new_n654), .B2(new_n370), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n650), .B1(new_n653), .B2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n359), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n643), .A2(new_n649), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G143), .ZN(G45));
  OAI211_X1 g474(.A(new_n476), .B(new_n627), .C1(new_n591), .C2(new_n592), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n620), .A2(new_n632), .A3(new_n551), .A4(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G146), .ZN(G48));
  INV_X1    g478(.A(KEYINPUT106), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n585), .A2(new_n590), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(KEYINPUT97), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n585), .A2(new_n586), .A3(new_n590), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n570), .A2(new_n669), .A3(new_n476), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n541), .A2(new_n189), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(G469), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n673), .A2(new_n549), .A3(new_n543), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT105), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n673), .A2(KEYINPUT105), .A3(new_n549), .A4(new_n543), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n375), .A2(new_n665), .A3(new_n671), .A4(new_n678), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n355), .B1(new_n562), .B2(new_n563), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(new_n357), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n555), .A2(KEYINPUT32), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n681), .A2(new_n682), .A3(new_n374), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n683), .A2(new_n566), .A3(new_n671), .A4(new_n678), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(KEYINPUT106), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n679), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(KEYINPUT41), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G113), .ZN(G15));
  NAND4_X1  g502(.A1(new_n683), .A2(new_n566), .A3(new_n570), .A4(new_n678), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n689), .A2(new_n606), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(new_n311), .ZN(G18));
  INV_X1    g505(.A(new_n674), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n683), .A2(new_n518), .A3(new_n614), .A4(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G119), .ZN(G21));
  AOI21_X1  g508(.A(new_n516), .B1(new_n470), .B2(new_n475), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n695), .A2(new_n427), .A3(new_n426), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT107), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n695), .A2(KEYINPUT107), .A3(new_n427), .A4(new_n426), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n243), .A2(new_n250), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n371), .A2(new_n651), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n354), .B1(new_n561), .B2(new_n702), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n703), .B1(new_n564), .B2(G472), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n483), .B1(new_n676), .B2(new_n677), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n700), .A2(new_n701), .A3(new_n704), .A4(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G122), .ZN(G24));
  NOR2_X1   g521(.A1(new_n674), .A2(new_n428), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n704), .A2(new_n614), .A3(new_n662), .A4(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT108), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(new_n703), .ZN(new_n712));
  AOI21_X1  g526(.A(G902), .B1(new_n349), .B2(new_n351), .ZN(new_n713));
  OAI211_X1 g527(.A(new_n614), .B(new_n712), .C1(new_n713), .C2(new_n650), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n715), .A2(KEYINPUT108), .A3(new_n662), .A4(new_n708), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n711), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G125), .ZN(G27));
  NOR3_X1   g532(.A1(new_n550), .A2(new_n648), .A3(new_n426), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n683), .A2(new_n566), .A3(new_n662), .A4(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(KEYINPUT109), .A2(KEYINPUT42), .ZN(new_n721));
  OR2_X1    g535(.A1(KEYINPUT109), .A2(KEYINPUT42), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n720), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT110), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n720), .A2(KEYINPUT110), .A3(new_n721), .A4(new_n722), .ZN(new_n726));
  AND2_X1   g540(.A1(new_n683), .A2(new_n701), .ZN(new_n727));
  AND3_X1   g541(.A1(new_n727), .A2(KEYINPUT42), .A3(new_n551), .ZN(new_n728));
  NOR3_X1   g542(.A1(new_n661), .A2(new_n648), .A3(new_n426), .ZN(new_n729));
  AOI22_X1  g543(.A1(new_n725), .A2(new_n726), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(new_n432), .ZN(G33));
  AND2_X1   g545(.A1(new_n375), .A2(new_n719), .ZN(new_n732));
  AND2_X1   g546(.A1(new_n628), .A2(new_n631), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G134), .ZN(G36));
  NOR2_X1   g549(.A1(new_n565), .A2(new_n619), .ZN(new_n736));
  AOI21_X1  g550(.A(KEYINPUT43), .B1(new_n669), .B2(new_n598), .ZN(new_n737));
  OAI211_X1 g551(.A(new_n598), .B(KEYINPUT43), .C1(new_n591), .C2(new_n592), .ZN(new_n738));
  INV_X1    g552(.A(new_n738), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n736), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(KEYINPUT44), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n426), .A2(new_n648), .ZN(new_n742));
  INV_X1    g556(.A(new_n549), .ZN(new_n743));
  OAI211_X1 g557(.A(new_n545), .B(KEYINPUT45), .C1(new_n546), .C2(new_n535), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT45), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n535), .B1(new_n525), .B2(new_n530), .ZN(new_n746));
  AND2_X1   g560(.A1(new_n536), .A2(new_n539), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n745), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n744), .A2(new_n748), .A3(G469), .ZN(new_n749));
  AOI21_X1  g563(.A(KEYINPUT46), .B1(new_n749), .B2(new_n544), .ZN(new_n750));
  INV_X1    g564(.A(new_n543), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n749), .A2(KEYINPUT46), .A3(new_n544), .ZN(new_n753));
  AOI211_X1 g567(.A(new_n743), .B(new_n639), .C1(new_n752), .C2(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n741), .A2(new_n742), .A3(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G137), .ZN(G39));
  INV_X1    g570(.A(KEYINPUT47), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n752), .A2(new_n753), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n757), .B1(new_n758), .B2(new_n549), .ZN(new_n759));
  AOI211_X1 g573(.A(KEYINPUT47), .B(new_n743), .C1(new_n752), .C2(new_n753), .ZN(new_n760));
  NOR3_X1   g574(.A1(new_n759), .A2(new_n760), .A3(new_n566), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n761), .A2(new_n359), .A3(new_n374), .A4(new_n729), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G140), .ZN(G42));
  INV_X1    g577(.A(KEYINPUT119), .ZN(new_n764));
  NOR2_X1   g578(.A1(G952), .A2(G953), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT53), .ZN(new_n766));
  XOR2_X1   g580(.A(new_n627), .B(KEYINPUT113), .Z(new_n767));
  NOR2_X1   g581(.A1(new_n614), .A2(new_n767), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n658), .A2(new_n551), .A3(new_n700), .A4(new_n768), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n636), .A2(new_n663), .A3(new_n717), .A4(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT52), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  AND4_X1   g586(.A1(new_n683), .A2(new_n635), .A3(new_n551), .A4(new_n614), .ZN(new_n773));
  AOI22_X1  g587(.A1(new_n773), .A2(new_n634), .B1(new_n711), .B2(new_n716), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n774), .A2(KEYINPUT52), .A3(new_n663), .A4(new_n769), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n772), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n683), .A2(new_n516), .A3(new_n604), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n704), .A2(new_n599), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n779), .A2(new_n614), .A3(new_n627), .A4(new_n719), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n734), .A2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT112), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n734), .A2(new_n780), .A3(KEYINPUT112), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n776), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n725), .A2(new_n726), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n728), .A2(new_n729), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n600), .B1(new_n516), .B2(new_n476), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n569), .A2(new_n570), .A3(new_n571), .A4(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n790), .A2(new_n553), .A3(new_n615), .ZN(new_n791));
  INV_X1    g605(.A(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n684), .B(new_n665), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n693), .B(new_n706), .C1(new_n689), .C2(new_n606), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n793), .A2(KEYINPUT111), .A3(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT111), .ZN(new_n796));
  INV_X1    g610(.A(new_n794), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n796), .B1(new_n797), .B2(new_n686), .ZN(new_n798));
  OAI211_X1 g612(.A(new_n788), .B(new_n792), .C1(new_n795), .C2(new_n798), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n766), .B1(new_n785), .B2(new_n799), .ZN(new_n800));
  NOR4_X1   g614(.A1(new_n730), .A2(new_n766), .A3(new_n793), .A4(new_n794), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n783), .A2(new_n784), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n801), .A2(new_n802), .A3(new_n792), .A4(new_n776), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT54), .ZN(new_n804));
  AND3_X1   g618(.A1(new_n800), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  AND3_X1   g619(.A1(new_n776), .A2(new_n783), .A3(new_n784), .ZN(new_n806));
  OAI21_X1  g620(.A(KEYINPUT111), .B1(new_n793), .B2(new_n794), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n797), .A2(new_n686), .A3(new_n796), .ZN(new_n808));
  AOI221_X4 g622(.A(new_n791), .B1(new_n786), .B2(new_n787), .C1(new_n807), .C2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n806), .A2(new_n809), .A3(KEYINPUT53), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n804), .B1(new_n810), .B2(new_n800), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n805), .A2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT43), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n813), .B1(new_n593), .B2(new_n476), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n623), .B1(new_n814), .B2(new_n738), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n427), .B1(new_n645), .B2(new_n646), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n816), .A2(new_n692), .A3(KEYINPUT114), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n815), .A2(new_n701), .A3(new_n817), .A4(new_n704), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n816), .A2(new_n692), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n819), .A2(KEYINPUT114), .ZN(new_n820));
  OAI21_X1  g634(.A(KEYINPUT115), .B1(new_n818), .B2(new_n820), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n622), .B1(new_n737), .B2(new_n739), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n704), .A2(new_n701), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT115), .ZN(new_n825));
  INV_X1    g639(.A(new_n820), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n824), .A2(new_n825), .A3(new_n826), .A4(new_n817), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT50), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n821), .A2(new_n827), .A3(KEYINPUT116), .A4(new_n828), .ZN(new_n829));
  NOR4_X1   g643(.A1(new_n822), .A2(new_n823), .A3(new_n648), .A4(new_n426), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n673), .A2(new_n543), .ZN(new_n831));
  OAI22_X1  g645(.A1(new_n759), .A2(new_n760), .B1(new_n549), .B2(new_n831), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n674), .A2(new_n648), .A3(new_n426), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n815), .A2(new_n833), .ZN(new_n834));
  AOI22_X1  g648(.A1(new_n830), .A2(new_n832), .B1(new_n715), .B2(new_n834), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n829), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n830), .A2(new_n832), .ZN(new_n837));
  AOI21_X1  g651(.A(KEYINPUT51), .B1(new_n837), .B2(KEYINPUT117), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n821), .A2(new_n827), .A3(new_n828), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n818), .A2(new_n820), .ZN(new_n840));
  AOI21_X1  g654(.A(KEYINPUT116), .B1(new_n840), .B2(KEYINPUT50), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n566), .A2(new_n833), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n658), .A2(new_n843), .A3(new_n478), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n844), .A2(new_n598), .A3(new_n593), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n836), .A2(new_n838), .A3(new_n842), .A4(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(new_n838), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n839), .A2(new_n841), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n829), .A2(new_n845), .A3(new_n835), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n847), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n846), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n834), .A2(new_n727), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n852), .B(KEYINPUT48), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n228), .A2(G952), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n854), .B1(new_n844), .B2(new_n599), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n824), .A2(new_n708), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n853), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(KEYINPUT118), .B1(new_n851), .B2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT118), .ZN(new_n860));
  AOI211_X1 g674(.A(new_n860), .B(new_n857), .C1(new_n846), .C2(new_n850), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n765), .B1(new_n812), .B2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(new_n658), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n593), .A2(new_n476), .ZN(new_n865));
  AND4_X1   g679(.A1(new_n701), .A2(new_n865), .A3(new_n427), .A4(new_n647), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n549), .B1(new_n831), .B2(KEYINPUT49), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n867), .B1(KEYINPUT49), .B2(new_n831), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n864), .A2(new_n866), .A3(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(new_n869), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n764), .B1(new_n863), .B2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(new_n800), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n785), .A2(new_n799), .A3(new_n766), .ZN(new_n873));
  OAI21_X1  g687(.A(KEYINPUT54), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n800), .A2(new_n803), .A3(new_n804), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n862), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(new_n765), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n878), .A2(KEYINPUT119), .A3(new_n869), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n871), .A2(new_n879), .ZN(G75));
  AOI21_X1  g694(.A(new_n189), .B1(new_n800), .B2(new_n803), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(G210), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n402), .A2(new_n408), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n883), .B(new_n406), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n884), .B(KEYINPUT55), .ZN(new_n885));
  XNOR2_X1  g699(.A(KEYINPUT120), .B(KEYINPUT56), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n882), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT56), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n885), .B1(new_n882), .B2(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n228), .A2(G952), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n887), .A2(new_n889), .A3(new_n890), .ZN(G51));
  XOR2_X1   g705(.A(new_n544), .B(KEYINPUT57), .Z(new_n892));
  AOI21_X1  g706(.A(new_n804), .B1(new_n800), .B2(new_n803), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n892), .B1(new_n805), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(new_n541), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n800), .A2(new_n803), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(G902), .ZN(new_n897));
  OR2_X1    g711(.A1(new_n897), .A2(new_n749), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n890), .B1(new_n895), .B2(new_n898), .ZN(G54));
  NAND2_X1  g713(.A1(KEYINPUT58), .A2(G475), .ZN(new_n900));
  OAI211_X1 g714(.A(new_n456), .B(new_n449), .C1(new_n897), .C2(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(new_n890), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n881), .A2(KEYINPUT58), .A3(G475), .A4(new_n457), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT121), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n901), .A2(KEYINPUT121), .A3(new_n902), .A4(new_n903), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(G60));
  NAND2_X1  g722(.A1(G478), .A2(G902), .ZN(new_n909));
  XOR2_X1   g723(.A(new_n909), .B(KEYINPUT59), .Z(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  OAI211_X1 g725(.A(new_n584), .B(new_n911), .C1(new_n805), .C2(new_n893), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n812), .A2(new_n910), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n902), .B(new_n912), .C1(new_n913), .C2(new_n584), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(G63));
  NAND2_X1  g729(.A1(G217), .A2(G902), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(KEYINPUT60), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n917), .B1(new_n800), .B2(new_n803), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n248), .A2(new_n249), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n902), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT61), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n918), .A2(new_n612), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n921), .A2(KEYINPUT122), .A3(new_n922), .A4(new_n923), .ZN(new_n924));
  OR2_X1    g738(.A1(new_n922), .A2(KEYINPUT122), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n922), .A2(KEYINPUT122), .ZN(new_n926));
  INV_X1    g740(.A(new_n923), .ZN(new_n927));
  OAI211_X1 g741(.A(new_n925), .B(new_n926), .C1(new_n927), .C2(new_n920), .ZN(new_n928));
  AND2_X1   g742(.A1(new_n924), .A2(new_n928), .ZN(G66));
  OAI21_X1  g743(.A(new_n792), .B1(new_n795), .B2(new_n798), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT123), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(new_n228), .ZN(new_n932));
  INV_X1    g746(.A(G224), .ZN(new_n933));
  OAI21_X1  g747(.A(G953), .B1(new_n481), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n883), .B1(G898), .B2(new_n228), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n935), .B(new_n936), .ZN(G69));
  INV_X1    g751(.A(G227), .ZN(new_n938));
  OAI21_X1  g752(.A(G953), .B1(new_n938), .B2(new_n624), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n939), .A2(KEYINPUT126), .ZN(new_n940));
  AND2_X1   g754(.A1(new_n774), .A2(new_n663), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(new_n659), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n942), .B(KEYINPUT62), .Z(new_n943));
  AND3_X1   g757(.A1(new_n732), .A2(new_n640), .A3(new_n789), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT124), .ZN(new_n945));
  OR2_X1    g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  AND2_X1   g760(.A1(new_n946), .A2(new_n755), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n944), .A2(new_n945), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n943), .A2(new_n947), .A3(new_n762), .A4(new_n948), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n340), .B(new_n441), .Z(new_n950));
  INV_X1    g764(.A(new_n950), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n949), .A2(new_n228), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n741), .A2(new_n742), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n727), .A2(new_n700), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  AOI22_X1  g769(.A1(new_n955), .A2(new_n754), .B1(new_n733), .B2(new_n732), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n956), .A2(new_n788), .A3(new_n762), .A4(new_n941), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(new_n228), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n624), .A2(G953), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(KEYINPUT125), .ZN(new_n960));
  INV_X1    g774(.A(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n958), .A2(new_n950), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n940), .B1(new_n952), .B2(new_n962), .ZN(new_n963));
  AND2_X1   g777(.A1(new_n939), .A2(KEYINPUT126), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n963), .B(new_n964), .ZN(G72));
  NAND2_X1  g779(.A1(G472), .A2(G902), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT63), .Z(new_n967));
  OAI21_X1  g781(.A(new_n967), .B1(new_n931), .B2(new_n957), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n968), .A2(new_n342), .A3(new_n654), .ZN(new_n969));
  INV_X1    g783(.A(new_n558), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n362), .B(KEYINPUT127), .ZN(new_n971));
  OAI221_X1 g785(.A(new_n967), .B1(new_n970), .B2(new_n971), .C1(new_n872), .C2(new_n873), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n969), .A2(new_n902), .A3(new_n972), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n967), .B1(new_n949), .B2(new_n931), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n973), .B1(new_n652), .B2(new_n974), .ZN(G57));
endmodule


