//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 0 0 1 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 0 0 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:41 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1336, new_n1337, new_n1338;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  OAI21_X1  g0011(.A(G50), .B1(G58), .B2(G68), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n206), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n217));
  INV_X1    g0017(.A(G244), .ZN(new_n218));
  INV_X1    g0018(.A(G87), .ZN(new_n219));
  INV_X1    g0019(.A(G250), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n217), .B1(new_n202), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n222));
  INV_X1    g0022(.A(G58), .ZN(new_n223));
  INV_X1    g0023(.A(G232), .ZN(new_n224));
  INV_X1    g0024(.A(G68), .ZN(new_n225));
  INV_X1    g0025(.A(G238), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n222), .B1(new_n223), .B2(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n208), .B1(new_n221), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n211), .B(new_n216), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XOR2_X1   g0030(.A(G226), .B(G232), .Z(new_n231));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n235), .B(new_n238), .Z(G358));
  XNOR2_X1  g0039(.A(G87), .B(G97), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT65), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G107), .ZN(new_n242));
  INV_X1    g0042(.A(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G68), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G351));
  NAND2_X1  g0048(.A1(G33), .A2(G41), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(KEYINPUT66), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT66), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n251), .A2(G33), .A3(G41), .ZN(new_n252));
  AND2_X1   g0052(.A1(G1), .A2(G13), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n250), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G41), .ZN(new_n255));
  INV_X1    g0055(.A(G45), .ZN(new_n256));
  AOI21_X1  g0056(.A(G1), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n254), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G238), .ZN(new_n261));
  AND2_X1   g0061(.A1(KEYINPUT3), .A2(G33), .ZN(new_n262));
  NOR2_X1   g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  OAI211_X1 g0063(.A(G232), .B(G1698), .C1(new_n262), .C2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(G33), .A2(G97), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G226), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n267), .A2(G1698), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT71), .ZN(new_n269));
  OAI211_X1 g0069(.A(new_n268), .B(new_n269), .C1(new_n263), .C2(new_n262), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n268), .B1(new_n262), .B2(new_n263), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(KEYINPUT71), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n266), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n253), .A2(new_n249), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT68), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n253), .A2(KEYINPUT68), .A3(new_n249), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n261), .B1(new_n273), .B2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G274), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n214), .B1(KEYINPUT66), .B2(new_n249), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n281), .B1(new_n282), .B2(new_n252), .ZN(new_n283));
  AOI21_X1  g0083(.A(KEYINPUT67), .B1(new_n283), .B2(new_n257), .ZN(new_n284));
  NAND4_X1  g0084(.A1(new_n254), .A2(KEYINPUT67), .A3(G274), .A4(new_n257), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  OAI21_X1  g0087(.A(KEYINPUT13), .B1(new_n280), .B2(new_n287), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n259), .A2(new_n226), .ZN(new_n289));
  INV_X1    g0089(.A(new_n265), .ZN(new_n290));
  INV_X1    g0090(.A(G1698), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT3), .ZN(new_n292));
  INV_X1    g0092(.A(G33), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(KEYINPUT3), .A2(G33), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n291), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n290), .B1(new_n296), .B2(G232), .ZN(new_n297));
  INV_X1    g0097(.A(new_n270), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n294), .A2(new_n295), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n269), .B1(new_n299), .B2(new_n268), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n297), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n289), .B1(new_n301), .B2(new_n278), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n254), .A2(G274), .A3(new_n257), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT67), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(new_n285), .ZN(new_n306));
  XNOR2_X1  g0106(.A(KEYINPUT72), .B(KEYINPUT13), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n302), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n288), .A2(G179), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(KEYINPUT74), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT74), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n288), .A2(new_n308), .A3(new_n311), .A4(G179), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n308), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n307), .B1(new_n302), .B2(new_n306), .ZN(new_n315));
  OAI21_X1  g0115(.A(G169), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(KEYINPUT14), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT14), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n318), .B(G169), .C1(new_n314), .C2(new_n315), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n313), .A2(new_n317), .A3(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(new_n214), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n206), .A2(G33), .ZN(new_n324));
  OAI22_X1  g0124(.A1(new_n324), .A2(new_n202), .B1(new_n206), .B2(G68), .ZN(new_n325));
  OR2_X1    g0125(.A1(new_n325), .A2(KEYINPUT73), .ZN(new_n326));
  NOR2_X1   g0126(.A1(G20), .A2(G33), .ZN(new_n327));
  AOI22_X1  g0127(.A1(new_n325), .A2(KEYINPUT73), .B1(G50), .B2(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n323), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(KEYINPUT11), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n331), .A2(G68), .ZN(new_n332));
  XNOR2_X1  g0132(.A(new_n332), .B(KEYINPUT12), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n322), .B1(new_n205), .B2(G20), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n333), .B1(G68), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n330), .A2(new_n335), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n329), .A2(KEYINPUT11), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  AND2_X1   g0139(.A1(new_n320), .A2(new_n339), .ZN(new_n340));
  OR2_X1    g0140(.A1(G223), .A2(G1698), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n267), .A2(G1698), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n341), .B(new_n342), .C1(new_n262), .C2(new_n263), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n343), .B1(new_n293), .B2(new_n219), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT76), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n343), .B(KEYINPUT76), .C1(new_n293), .C2(new_n219), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n346), .A2(new_n347), .A3(new_n278), .ZN(new_n348));
  AND3_X1   g0148(.A1(new_n254), .A2(G232), .A3(new_n258), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n349), .B1(new_n305), .B2(new_n285), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT77), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n348), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  AOI211_X1 g0152(.A(KEYINPUT77), .B(new_n349), .C1(new_n305), .C2(new_n285), .ZN(new_n353));
  OAI21_X1  g0153(.A(G169), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(KEYINPUT77), .B1(new_n287), .B2(new_n349), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n350), .A2(new_n351), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n355), .A2(G179), .A3(new_n356), .A4(new_n348), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n323), .A2(new_n331), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT69), .ZN(new_n360));
  XNOR2_X1  g0160(.A(new_n359), .B(new_n360), .ZN(new_n361));
  XNOR2_X1  g0161(.A(KEYINPUT8), .B(G58), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n205), .A2(G20), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n331), .ZN(new_n367));
  AOI22_X1  g0167(.A1(new_n361), .A2(new_n366), .B1(new_n367), .B2(new_n362), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT75), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n294), .A2(new_n206), .A3(new_n295), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT7), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n294), .A2(KEYINPUT7), .A3(new_n206), .A4(new_n295), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n369), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(KEYINPUT75), .B1(new_n370), .B2(new_n371), .ZN(new_n375));
  OAI21_X1  g0175(.A(G68), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n223), .A2(new_n225), .ZN(new_n377));
  NOR2_X1   g0177(.A1(G58), .A2(G68), .ZN(new_n378));
  OAI21_X1  g0178(.A(G20), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n327), .A2(G159), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(KEYINPUT16), .B1(new_n376), .B2(new_n382), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n262), .A2(new_n263), .ZN(new_n384));
  AOI21_X1  g0184(.A(KEYINPUT7), .B1(new_n384), .B2(new_n206), .ZN(new_n385));
  INV_X1    g0185(.A(new_n373), .ZN(new_n386));
  OAI21_X1  g0186(.A(G68), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n387), .A2(KEYINPUT16), .A3(new_n382), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(new_n322), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n368), .B1(new_n383), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n358), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(KEYINPUT18), .ZN(new_n392));
  XNOR2_X1  g0192(.A(new_n359), .B(KEYINPUT69), .ZN(new_n393));
  OAI22_X1  g0193(.A1(new_n393), .A2(new_n365), .B1(new_n331), .B2(new_n363), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT16), .ZN(new_n395));
  OAI21_X1  g0195(.A(KEYINPUT75), .B1(new_n385), .B2(new_n386), .ZN(new_n396));
  INV_X1    g0196(.A(new_n375), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n225), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n395), .B1(new_n398), .B2(new_n381), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n225), .B1(new_n372), .B2(new_n373), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n400), .A2(new_n381), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n323), .B1(new_n401), .B2(KEYINPUT16), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n394), .B1(new_n399), .B2(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n403), .B1(new_n354), .B2(new_n357), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT18), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(G200), .B1(new_n352), .B2(new_n353), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n355), .A2(G190), .A3(new_n356), .A4(new_n348), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n403), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  AND2_X1   g0209(.A1(new_n409), .A2(KEYINPUT17), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n409), .A2(KEYINPUT17), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n392), .B(new_n406), .C1(new_n410), .C2(new_n411), .ZN(new_n412));
  XNOR2_X1  g0212(.A(KEYINPUT15), .B(G87), .ZN(new_n413));
  OAI22_X1  g0213(.A1(new_n413), .A2(new_n324), .B1(new_n206), .B2(new_n202), .ZN(new_n414));
  XOR2_X1   g0214(.A(new_n362), .B(KEYINPUT70), .Z(new_n415));
  AOI21_X1  g0215(.A(new_n414), .B1(new_n415), .B2(new_n327), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n416), .A2(new_n323), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n334), .A2(G77), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(G77), .B2(new_n331), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(G238), .A2(G1698), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n299), .B(new_n421), .C1(new_n224), .C2(G1698), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n278), .B(new_n422), .C1(G107), .C2(new_n299), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n306), .B(new_n423), .C1(new_n218), .C2(new_n259), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(G200), .ZN(new_n425));
  INV_X1    g0225(.A(G190), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n420), .B(new_n425), .C1(new_n426), .C2(new_n424), .ZN(new_n427));
  INV_X1    g0227(.A(G169), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n424), .A2(new_n428), .ZN(new_n429));
  OAI221_X1 g0229(.A(new_n429), .B1(G179), .B2(new_n424), .C1(new_n417), .C2(new_n419), .ZN(new_n430));
  AND2_X1   g0230(.A1(new_n427), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n291), .A2(G222), .ZN(new_n432));
  NAND2_X1  g0232(.A1(G223), .A2(G1698), .ZN(new_n433));
  AND3_X1   g0233(.A1(new_n299), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n434), .B1(new_n202), .B2(new_n384), .ZN(new_n435));
  AOI22_X1  g0235(.A1(new_n435), .A2(new_n278), .B1(G226), .B2(new_n260), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(new_n306), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(G179), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n361), .A2(G50), .A3(new_n364), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n327), .A2(G150), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n442), .B1(new_n362), .B2(new_n324), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n201), .A2(new_n206), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n322), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(G50), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n367), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n441), .A2(new_n449), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n440), .B(new_n450), .C1(G169), .C2(new_n438), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n364), .A2(G50), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n393), .A2(new_n452), .ZN(new_n453));
  OAI21_X1  g0253(.A(KEYINPUT9), .B1(new_n453), .B2(new_n448), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT9), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n441), .A2(new_n455), .A3(new_n449), .ZN(new_n456));
  AOI22_X1  g0256(.A1(new_n454), .A2(new_n456), .B1(new_n437), .B2(G200), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT10), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n438), .A2(G190), .ZN(new_n459));
  AND3_X1   g0259(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n458), .B1(new_n457), .B2(new_n459), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n431), .B(new_n451), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n288), .A2(G190), .A3(new_n308), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(new_n338), .ZN(new_n464));
  INV_X1    g0264(.A(G200), .ZN(new_n465));
  INV_X1    g0265(.A(new_n315), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n465), .B1(new_n466), .B2(new_n308), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  NOR4_X1   g0268(.A1(new_n340), .A2(new_n412), .A3(new_n462), .A4(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n205), .A2(G33), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n331), .A2(new_n470), .A3(new_n214), .A4(new_n321), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(G97), .ZN(new_n472));
  INV_X1    g0272(.A(G97), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n331), .A2(new_n473), .ZN(new_n474));
  AND3_X1   g0274(.A1(new_n472), .A2(KEYINPUT78), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g0275(.A(KEYINPUT78), .B1(new_n472), .B2(new_n474), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g0277(.A(G107), .B1(new_n374), .B2(new_n375), .ZN(new_n478));
  INV_X1    g0278(.A(G107), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n479), .A2(KEYINPUT6), .A3(G97), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n473), .A2(new_n479), .ZN(new_n481));
  NOR2_X1   g0281(.A1(G97), .A2(G107), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n480), .B1(new_n483), .B2(KEYINPUT6), .ZN(new_n484));
  AOI22_X1  g0284(.A1(new_n484), .A2(G20), .B1(G77), .B2(new_n327), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n478), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n477), .B1(new_n486), .B2(new_n322), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n255), .A2(KEYINPUT5), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n205), .A2(G45), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n255), .A2(KEYINPUT5), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n254), .A2(new_n490), .A3(G274), .A4(new_n491), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n256), .A2(G1), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT5), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(G41), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n493), .A2(new_n491), .A3(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n254), .A2(new_n496), .A3(G257), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n492), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n220), .B1(new_n294), .B2(new_n295), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT4), .ZN(new_n500));
  OAI21_X1  g0300(.A(G1698), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n500), .B1(new_n384), .B2(new_n218), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n500), .A2(G1698), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n503), .B(G244), .C1(new_n263), .C2(new_n262), .ZN(new_n504));
  NAND2_X1  g0304(.A1(G33), .A2(G283), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n501), .A2(new_n502), .A3(new_n504), .A4(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n498), .B1(new_n506), .B2(new_n278), .ZN(new_n507));
  OAI21_X1  g0307(.A(KEYINPUT79), .B1(new_n507), .B2(new_n465), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(G190), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n218), .B1(new_n294), .B2(new_n295), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n504), .B(new_n505), .C1(new_n510), .C2(KEYINPUT4), .ZN(new_n511));
  OAI21_X1  g0311(.A(G250), .B1(new_n262), .B2(new_n263), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n291), .B1(new_n512), .B2(KEYINPUT4), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n278), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  AND2_X1   g0314(.A1(new_n492), .A2(new_n497), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT79), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n516), .A2(new_n517), .A3(G200), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n487), .A2(new_n508), .A3(new_n509), .A4(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n514), .A2(new_n439), .A3(new_n515), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n323), .B1(new_n478), .B2(new_n485), .ZN(new_n521));
  OAI221_X1 g0321(.A(new_n520), .B1(G169), .B2(new_n507), .C1(new_n521), .C2(new_n477), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n367), .A2(new_n479), .ZN(new_n523));
  OR2_X1    g0323(.A1(new_n523), .A2(KEYINPUT25), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(KEYINPUT25), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n524), .B(new_n525), .C1(new_n479), .C2(new_n471), .ZN(new_n526));
  AND2_X1   g0326(.A1(KEYINPUT82), .A2(KEYINPUT22), .ZN(new_n527));
  NOR2_X1   g0327(.A1(KEYINPUT82), .A2(KEYINPUT22), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n299), .A2(new_n529), .A3(new_n206), .A4(G87), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n206), .B(G87), .C1(new_n262), .C2(new_n263), .ZN(new_n531));
  OR2_X1    g0331(.A1(new_n527), .A2(new_n528), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  OAI211_X1 g0333(.A(KEYINPUT83), .B(KEYINPUT23), .C1(new_n206), .C2(G107), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n206), .A2(G33), .A3(G116), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT23), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n536), .A2(new_n479), .A3(G20), .ZN(new_n537));
  AND3_X1   g0337(.A1(new_n534), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  OAI21_X1  g0338(.A(KEYINPUT23), .B1(new_n206), .B2(G107), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT83), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n530), .A2(new_n533), .A3(new_n538), .A4(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(KEYINPUT24), .ZN(new_n543));
  AND4_X1   g0343(.A1(new_n541), .A2(new_n534), .A3(new_n535), .A4(new_n537), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT24), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n544), .A2(new_n545), .A3(new_n533), .A4(new_n530), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n526), .B1(new_n547), .B2(new_n322), .ZN(new_n548));
  OAI211_X1 g0348(.A(G250), .B(new_n291), .C1(new_n262), .C2(new_n263), .ZN(new_n549));
  OAI211_X1 g0349(.A(G257), .B(G1698), .C1(new_n262), .C2(new_n263), .ZN(new_n550));
  NAND2_X1  g0350(.A1(G33), .A2(G294), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n278), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n254), .A2(new_n496), .A3(G264), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n553), .A2(new_n492), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(G200), .ZN(new_n556));
  AND2_X1   g0356(.A1(new_n254), .A2(new_n496), .ZN(new_n557));
  AOI22_X1  g0357(.A1(G264), .A2(new_n557), .B1(new_n552), .B2(new_n278), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n558), .A2(G190), .A3(new_n492), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n548), .A2(new_n556), .A3(new_n559), .ZN(new_n560));
  AND3_X1   g0360(.A1(new_n519), .A2(new_n522), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(KEYINPUT84), .B1(new_n555), .B2(G169), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n555), .A2(new_n439), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AND3_X1   g0364(.A1(new_n555), .A2(KEYINPUT84), .A3(G169), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n548), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n413), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n568), .A2(new_n331), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n219), .A2(KEYINPUT81), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT81), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(G87), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n570), .A2(new_n572), .A3(new_n482), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT19), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n574), .B1(new_n265), .B2(new_n206), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n299), .A2(new_n206), .A3(G68), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n574), .B1(new_n324), .B2(new_n473), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n569), .B1(new_n579), .B2(new_n322), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n580), .B1(new_n413), .B2(new_n471), .ZN(new_n581));
  OAI211_X1 g0381(.A(G244), .B(G1698), .C1(new_n262), .C2(new_n263), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT80), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n293), .A2(new_n243), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n226), .A2(G1698), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n585), .B1(new_n299), .B2(new_n586), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n299), .A2(KEYINPUT80), .A3(G244), .A4(G1698), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n584), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n278), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n489), .A2(new_n220), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n493), .A2(new_n281), .ZN(new_n592));
  AND3_X1   g0392(.A1(new_n254), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n428), .B1(new_n590), .B2(new_n594), .ZN(new_n595));
  AOI211_X1 g0395(.A(new_n439), .B(new_n593), .C1(new_n589), .C2(new_n278), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n581), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n590), .A2(G190), .A3(new_n594), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n471), .A2(new_n219), .ZN(new_n599));
  AOI211_X1 g0399(.A(new_n569), .B(new_n599), .C1(new_n579), .C2(new_n322), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n593), .B1(new_n589), .B2(new_n278), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n598), .B(new_n600), .C1(new_n465), .C2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n597), .A2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(G303), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n294), .A2(new_n604), .A3(new_n295), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n291), .A2(G257), .ZN(new_n606));
  NAND2_X1  g0406(.A1(G264), .A2(G1698), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n606), .B(new_n607), .C1(new_n262), .C2(new_n263), .ZN(new_n608));
  AND4_X1   g0408(.A1(KEYINPUT68), .A2(new_n249), .A3(G1), .A4(G13), .ZN(new_n609));
  AOI21_X1  g0409(.A(KEYINPUT68), .B1(new_n253), .B2(new_n249), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n605), .B(new_n608), .C1(new_n609), .C2(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n254), .A2(new_n496), .A3(G270), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n611), .A2(new_n492), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(G200), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n505), .B(new_n206), .C1(G33), .C2(new_n473), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n243), .A2(G20), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n615), .A2(new_n322), .A3(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT20), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n615), .A2(KEYINPUT20), .A3(new_n322), .A4(new_n616), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n471), .A2(G116), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n331), .A2(new_n243), .ZN(new_n622));
  AOI22_X1  g0422(.A1(new_n619), .A2(new_n620), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n614), .B(new_n623), .C1(new_n426), .C2(new_n613), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT21), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n613), .A2(G169), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n625), .B1(new_n626), .B2(new_n623), .ZN(new_n627));
  INV_X1    g0427(.A(new_n613), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n619), .A2(new_n620), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n621), .A2(new_n622), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n628), .A2(new_n631), .A3(G179), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n631), .A2(KEYINPUT21), .A3(G169), .A4(new_n613), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n624), .A2(new_n627), .A3(new_n632), .A4(new_n633), .ZN(new_n634));
  NOR3_X1   g0434(.A1(new_n567), .A2(new_n603), .A3(new_n634), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n469), .A2(new_n561), .A3(new_n635), .ZN(G372));
  INV_X1    g0436(.A(new_n451), .ZN(new_n637));
  XNOR2_X1  g0437(.A(new_n409), .B(KEYINPUT17), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n468), .A2(new_n430), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n638), .B1(new_n340), .B2(new_n639), .ZN(new_n640));
  AND3_X1   g0440(.A1(new_n358), .A2(new_n405), .A3(new_n390), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n405), .B1(new_n358), .B2(new_n390), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  OR2_X1    g0444(.A1(new_n460), .A2(new_n461), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n637), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n469), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n520), .B1(new_n507), .B2(G169), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n487), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n516), .A2(new_n426), .ZN(new_n650));
  NOR3_X1   g0450(.A1(new_n650), .A2(new_n521), .A3(new_n477), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n508), .A2(new_n518), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n649), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n602), .ZN(new_n654));
  INV_X1    g0454(.A(new_n581), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n590), .A2(G179), .A3(new_n594), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n656), .B1(new_n428), .B2(new_n601), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT85), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n655), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  OAI211_X1 g0459(.A(new_n656), .B(KEYINPUT85), .C1(new_n428), .C2(new_n601), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n654), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n627), .A2(new_n632), .A3(new_n633), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NOR3_X1   g0463(.A1(new_n565), .A2(new_n562), .A3(new_n563), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n663), .B1(new_n664), .B2(new_n548), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n653), .A2(new_n661), .A3(new_n665), .A4(new_n560), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n658), .B1(new_n595), .B2(new_n596), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n667), .A2(new_n660), .A3(new_n581), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n668), .A2(new_n649), .A3(new_n602), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT86), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT26), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n670), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n670), .A2(new_n672), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n522), .A2(new_n603), .ZN(new_n675));
  AOI22_X1  g0475(.A1(new_n674), .A2(KEYINPUT86), .B1(KEYINPUT26), .B2(new_n675), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n669), .B1(new_n673), .B2(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n646), .B1(new_n647), .B2(new_n677), .ZN(G369));
  NAND2_X1  g0478(.A1(new_n564), .A2(new_n566), .ZN(new_n679));
  INV_X1    g0479(.A(new_n548), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n560), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n205), .A2(new_n206), .A3(G13), .ZN(new_n683));
  OR2_X1    g0483(.A1(new_n683), .A2(KEYINPUT27), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(KEYINPUT27), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n684), .A2(new_n685), .A3(G213), .ZN(new_n686));
  INV_X1    g0486(.A(G343), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n548), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n681), .B1(new_n682), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n567), .A2(new_n689), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n689), .A2(new_n623), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n662), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n695), .B1(new_n634), .B2(new_n694), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(G330), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n693), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n681), .A2(new_n688), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n662), .A2(new_n689), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(KEYINPUT87), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT87), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n662), .A2(new_n703), .A3(new_n689), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n700), .B1(new_n691), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n699), .A2(new_n706), .ZN(G399));
  INV_X1    g0507(.A(new_n209), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n708), .A2(G41), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(G1), .ZN(new_n711));
  OR2_X1    g0511(.A1(new_n573), .A2(G116), .ZN(new_n712));
  OAI22_X1  g0512(.A1(new_n711), .A2(new_n712), .B1(new_n212), .B2(new_n710), .ZN(new_n713));
  XOR2_X1   g0513(.A(new_n713), .B(KEYINPUT28), .Z(new_n714));
  NAND4_X1  g0514(.A1(new_n668), .A2(KEYINPUT26), .A3(new_n649), .A4(new_n602), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n672), .B1(new_n522), .B2(new_n603), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n666), .A2(new_n668), .A3(new_n717), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n718), .A2(KEYINPUT29), .A3(new_n689), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT91), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n718), .A2(KEYINPUT91), .A3(KEYINPUT29), .A4(new_n689), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n674), .A2(KEYINPUT86), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n675), .A2(KEYINPUT26), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n723), .A2(new_n673), .A3(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n519), .A2(new_n560), .A3(new_n522), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n668), .A2(new_n602), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  AOI22_X1  g0528(.A1(new_n728), .A2(new_n665), .B1(new_n660), .B2(new_n659), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n688), .B1(new_n725), .B2(new_n729), .ZN(new_n730));
  OAI211_X1 g0530(.A(new_n721), .B(new_n722), .C1(KEYINPUT29), .C2(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n635), .A2(new_n561), .A3(new_n689), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(KEYINPUT90), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n611), .A2(new_n492), .A3(new_n612), .A4(G179), .ZN(new_n734));
  XNOR2_X1  g0534(.A(new_n734), .B(KEYINPUT89), .ZN(new_n735));
  AND3_X1   g0535(.A1(new_n601), .A2(KEYINPUT88), .A3(new_n558), .ZN(new_n736));
  AOI21_X1  g0536(.A(KEYINPUT88), .B1(new_n601), .B2(new_n558), .ZN(new_n737));
  OAI211_X1 g0537(.A(new_n735), .B(new_n507), .C1(new_n736), .C2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT30), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  OR2_X1    g0540(.A1(new_n734), .A2(KEYINPUT89), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n734), .A2(KEYINPUT89), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n516), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  OAI211_X1 g0543(.A(new_n743), .B(KEYINPUT30), .C1(new_n737), .C2(new_n736), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n628), .A2(G179), .ZN(new_n745));
  INV_X1    g0545(.A(new_n601), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n745), .A2(new_n746), .A3(new_n516), .A4(new_n555), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n740), .A2(new_n744), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(new_n688), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT31), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT90), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n635), .A2(new_n561), .A3(new_n752), .A4(new_n689), .ZN(new_n753));
  INV_X1    g0553(.A(new_n747), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n754), .B1(new_n738), .B2(new_n739), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n689), .B1(new_n755), .B2(new_n744), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(KEYINPUT31), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n733), .A2(new_n751), .A3(new_n753), .A4(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(G330), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n731), .A2(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n714), .B1(new_n760), .B2(new_n205), .ZN(new_n761));
  XNOR2_X1  g0561(.A(new_n761), .B(KEYINPUT92), .ZN(G364));
  NOR2_X1   g0562(.A1(G13), .A2(G33), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(G20), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n214), .B1(G20), .B2(new_n428), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g0567(.A(new_n767), .B(KEYINPUT94), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n708), .A2(new_n299), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n247), .A2(G45), .ZN(new_n771));
  XOR2_X1   g0571(.A(new_n771), .B(KEYINPUT93), .Z(new_n772));
  AOI211_X1 g0572(.A(new_n770), .B(new_n772), .C1(new_n256), .C2(new_n213), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n708), .A2(new_n384), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G355), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n775), .B1(G116), .B2(new_n209), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n768), .B1(new_n773), .B2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(G13), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(G20), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n205), .B1(new_n779), .B2(G45), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n709), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n777), .A2(new_n782), .ZN(new_n783));
  NOR3_X1   g0583(.A1(new_n426), .A2(G179), .A3(G200), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(new_n206), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(new_n473), .ZN(new_n786));
  NAND2_X1  g0586(.A1(G20), .A2(G179), .ZN(new_n787));
  NOR3_X1   g0587(.A1(new_n787), .A2(G190), .A3(G200), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NOR3_X1   g0589(.A1(new_n787), .A2(new_n426), .A3(G200), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  OAI221_X1 g0591(.A(new_n299), .B1(new_n789), .B2(new_n202), .C1(new_n223), .C2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n787), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n793), .A2(G190), .A3(G200), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  AOI211_X1 g0595(.A(new_n786), .B(new_n792), .C1(G50), .C2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n206), .A2(G190), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n797), .A2(new_n439), .A3(new_n465), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(G159), .ZN(new_n800));
  XNOR2_X1  g0600(.A(new_n800), .B(KEYINPUT32), .ZN(new_n801));
  NOR3_X1   g0601(.A1(new_n787), .A2(new_n465), .A3(G190), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n801), .B1(G68), .B2(new_n802), .ZN(new_n803));
  OR3_X1    g0603(.A1(new_n465), .A2(KEYINPUT95), .A3(G179), .ZN(new_n804));
  OAI21_X1  g0604(.A(KEYINPUT95), .B1(new_n465), .B2(G179), .ZN(new_n805));
  NAND4_X1  g0605(.A1(new_n804), .A2(G20), .A3(G190), .A4(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n806), .B1(new_n570), .B2(new_n572), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n804), .A2(new_n805), .A3(new_n797), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n807), .B1(G107), .B2(new_n809), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n796), .A2(new_n803), .A3(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(KEYINPUT33), .A2(G317), .ZN(new_n812));
  AND2_X1   g0612(.A1(KEYINPUT33), .A2(G317), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n802), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(G326), .ZN(new_n815));
  INV_X1    g0615(.A(G294), .ZN(new_n816));
  OAI221_X1 g0616(.A(new_n814), .B1(new_n815), .B2(new_n794), .C1(new_n816), .C2(new_n785), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n799), .A2(G329), .B1(new_n790), .B2(G322), .ZN(new_n818));
  INV_X1    g0618(.A(G311), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n818), .B1(new_n819), .B2(new_n789), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n817), .B(new_n820), .C1(G283), .C2(new_n809), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n806), .B(KEYINPUT96), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n299), .B1(new_n822), .B2(G303), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(KEYINPUT97), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n823), .A2(KEYINPUT97), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n811), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n783), .B1(new_n766), .B2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n765), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n828), .B1(new_n696), .B2(new_n829), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n830), .B(KEYINPUT98), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n696), .A2(G330), .ZN(new_n832));
  INV_X1    g0632(.A(new_n782), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n697), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n831), .B1(new_n832), .B2(new_n834), .ZN(G396));
  NAND2_X1  g0635(.A1(new_n725), .A2(new_n729), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n836), .A2(new_n431), .A3(new_n689), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n427), .B1(new_n420), .B2(new_n689), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(new_n430), .ZN(new_n839));
  OR2_X1    g0639(.A1(new_n430), .A2(new_n688), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n837), .B1(new_n730), .B2(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n782), .B1(new_n843), .B2(new_n759), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n844), .B1(new_n759), .B2(new_n843), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n384), .B1(new_n791), .B2(new_n816), .ZN(new_n846));
  OAI22_X1  g0646(.A1(new_n789), .A2(new_n243), .B1(new_n798), .B2(new_n819), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n846), .B(new_n847), .C1(G87), .C2(new_n809), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n794), .A2(new_n604), .ZN(new_n849));
  XNOR2_X1  g0649(.A(KEYINPUT99), .B(G283), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  AOI211_X1 g0651(.A(new_n849), .B(new_n786), .C1(new_n802), .C2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n822), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n848), .B(new_n852), .C1(new_n853), .C2(new_n479), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n785), .A2(new_n223), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n384), .B(new_n855), .C1(G132), .C2(new_n799), .ZN(new_n856));
  AOI22_X1  g0656(.A1(G143), .A2(new_n790), .B1(new_n788), .B2(G159), .ZN(new_n857));
  INV_X1    g0657(.A(G137), .ZN(new_n858));
  INV_X1    g0658(.A(G150), .ZN(new_n859));
  INV_X1    g0659(.A(new_n802), .ZN(new_n860));
  OAI221_X1 g0660(.A(new_n857), .B1(new_n858), .B2(new_n794), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT34), .ZN(new_n862));
  OAI221_X1 g0662(.A(new_n856), .B1(new_n225), .B2(new_n808), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n861), .A2(new_n862), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n864), .B1(new_n853), .B2(new_n446), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n854), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(new_n766), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n766), .A2(new_n763), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n833), .B1(new_n202), .B2(new_n868), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n867), .B(new_n869), .C1(new_n842), .C2(new_n764), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n845), .A2(new_n870), .ZN(G384));
  NAND2_X1  g0671(.A1(new_n320), .A2(new_n339), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n872), .A2(new_n688), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT38), .ZN(new_n874));
  INV_X1    g0674(.A(new_n686), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n390), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n876), .B1(new_n643), .B2(new_n638), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n409), .A2(new_n876), .ZN(new_n878));
  OAI21_X1  g0678(.A(KEYINPUT37), .B1(new_n878), .B2(new_n404), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT37), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n391), .A2(new_n880), .A3(new_n409), .A4(new_n876), .ZN(new_n881));
  AND2_X1   g0681(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n874), .B1(new_n877), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n395), .B1(new_n400), .B2(new_n381), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n402), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n368), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n875), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n412), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n409), .A2(new_n887), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n354), .A2(new_n357), .B1(new_n368), .B2(new_n885), .ZN(new_n891));
  OAI21_X1  g0691(.A(KEYINPUT37), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n881), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n889), .A2(KEYINPUT38), .A3(new_n893), .ZN(new_n894));
  XNOR2_X1  g0694(.A(KEYINPUT100), .B(KEYINPUT39), .ZN(new_n895));
  AND3_X1   g0695(.A1(new_n883), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT39), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n887), .B1(new_n643), .B2(new_n638), .ZN(new_n898));
  AND2_X1   g0698(.A1(new_n892), .A2(new_n881), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n874), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n897), .B1(new_n900), .B2(new_n894), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n873), .B1(new_n896), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n837), .A2(new_n840), .ZN(new_n903));
  INV_X1    g0703(.A(new_n468), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n339), .A2(new_n688), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n872), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n339), .B(new_n688), .C1(new_n320), .C2(new_n468), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(KEYINPUT38), .B1(new_n889), .B2(new_n893), .ZN(new_n909));
  AOI221_X4 g0709(.A(new_n874), .B1(new_n892), .B2(new_n881), .C1(new_n412), .C2(new_n888), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n903), .B(new_n908), .C1(new_n909), .C2(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n643), .A2(new_n875), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n902), .A2(new_n911), .A3(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT101), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(KEYINPUT39), .B1(new_n910), .B2(new_n909), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n883), .A2(new_n894), .A3(new_n895), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n912), .B1(new_n919), .B2(new_n873), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n920), .A2(KEYINPUT101), .A3(new_n911), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n916), .A2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT29), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n677), .B2(new_n688), .ZN(new_n924));
  NAND4_X1  g0724(.A1(new_n924), .A2(new_n469), .A3(new_n722), .A4(new_n721), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n646), .ZN(new_n926));
  XOR2_X1   g0726(.A(new_n926), .B(KEYINPUT102), .Z(new_n927));
  XNOR2_X1  g0727(.A(new_n922), .B(new_n927), .ZN(new_n928));
  AOI22_X1  g0728(.A1(new_n732), .A2(KEYINPUT90), .B1(new_n756), .B2(KEYINPUT31), .ZN(new_n929));
  OAI21_X1  g0729(.A(KEYINPUT103), .B1(new_n756), .B2(KEYINPUT31), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT103), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n749), .A2(new_n931), .A3(new_n750), .ZN(new_n932));
  NAND4_X1  g0732(.A1(new_n929), .A2(new_n753), .A3(new_n930), .A4(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n841), .B1(new_n906), .B2(new_n907), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n933), .B(new_n934), .C1(new_n910), .C2(new_n909), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT40), .ZN(new_n936));
  AND2_X1   g0736(.A1(new_n933), .A2(new_n934), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n936), .B1(new_n883), .B2(new_n894), .ZN(new_n938));
  AOI22_X1  g0738(.A1(new_n935), .A2(new_n936), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n469), .A2(new_n933), .ZN(new_n941));
  OAI21_X1  g0741(.A(G330), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n942), .B1(new_n941), .B2(new_n940), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n928), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n928), .A2(new_n943), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n945), .B1(new_n205), .B2(new_n779), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n944), .B1(new_n946), .B2(KEYINPUT104), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(KEYINPUT104), .B2(new_n946), .ZN(new_n948));
  OR2_X1    g0748(.A1(new_n484), .A2(KEYINPUT35), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n484), .A2(KEYINPUT35), .ZN(new_n950));
  NAND4_X1  g0750(.A1(new_n949), .A2(G116), .A3(new_n215), .A4(new_n950), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT36), .ZN(new_n952));
  NOR3_X1   g0752(.A1(new_n377), .A2(new_n212), .A3(new_n202), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n225), .A2(G50), .ZN(new_n954));
  OAI211_X1 g0754(.A(G1), .B(new_n778), .C1(new_n953), .C2(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n948), .A2(new_n952), .A3(new_n955), .ZN(G367));
  OAI21_X1  g0756(.A(new_n767), .B1(new_n209), .B2(new_n413), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n957), .B1(new_n769), .B2(new_n238), .ZN(new_n958));
  INV_X1    g0758(.A(G159), .ZN(new_n959));
  INV_X1    g0759(.A(G143), .ZN(new_n960));
  OAI22_X1  g0760(.A1(new_n860), .A2(new_n959), .B1(new_n794), .B2(new_n960), .ZN(new_n961));
  OAI22_X1  g0761(.A1(new_n791), .A2(new_n859), .B1(new_n789), .B2(new_n446), .ZN(new_n962));
  AOI211_X1 g0762(.A(new_n384), .B(new_n962), .C1(G137), .C2(new_n799), .ZN(new_n963));
  OAI221_X1 g0763(.A(new_n963), .B1(new_n223), .B2(new_n806), .C1(new_n202), .C2(new_n808), .ZN(new_n964));
  INV_X1    g0764(.A(new_n785), .ZN(new_n965));
  AOI211_X1 g0765(.A(new_n961), .B(new_n964), .C1(G68), .C2(new_n965), .ZN(new_n966));
  AOI22_X1  g0766(.A1(new_n965), .A2(G107), .B1(new_n795), .B2(G311), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n816), .B2(new_n860), .ZN(new_n968));
  INV_X1    g0768(.A(new_n806), .ZN(new_n969));
  AOI21_X1  g0769(.A(KEYINPUT46), .B1(new_n969), .B2(G116), .ZN(new_n970));
  AOI22_X1  g0770(.A1(new_n799), .A2(G317), .B1(new_n851), .B2(new_n788), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n299), .B1(G303), .B2(new_n790), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n808), .A2(new_n473), .ZN(new_n974));
  NOR4_X1   g0774(.A1(new_n968), .A2(new_n970), .A3(new_n973), .A4(new_n974), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n822), .A2(KEYINPUT46), .A3(G116), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT110), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n966), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n978), .B(KEYINPUT47), .Z(new_n979));
  AOI211_X1 g0779(.A(new_n833), .B(new_n958), .C1(new_n979), .C2(new_n766), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n600), .A2(new_n689), .ZN(new_n981));
  MUX2_X1   g0781(.A(new_n727), .B(new_n668), .S(new_n981), .Z(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(new_n765), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n980), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n688), .B1(new_n521), .B2(new_n477), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n519), .A2(new_n522), .A3(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n649), .A2(new_n688), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n704), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n703), .B1(new_n662), .B2(new_n689), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n690), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n567), .B1(new_n992), .B2(new_n560), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n692), .B(new_n988), .C1(new_n991), .C2(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT45), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n706), .A2(KEYINPUT45), .A3(new_n988), .ZN(new_n997));
  AND2_X1   g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(KEYINPUT44), .B1(new_n706), .B2(new_n988), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n692), .B1(new_n991), .B2(new_n993), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT44), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n988), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n1000), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n999), .A2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n698), .B1(new_n998), .B2(new_n1004), .ZN(new_n1005));
  AND2_X1   g0805(.A1(new_n999), .A2(new_n1003), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n996), .A2(new_n997), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1006), .A2(new_n699), .A3(new_n1007), .ZN(new_n1008));
  AND2_X1   g0808(.A1(new_n1005), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n693), .A2(new_n991), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n691), .A2(new_n705), .A3(new_n692), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n697), .A2(KEYINPUT107), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1012), .B(new_n1013), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n760), .B1(new_n1009), .B2(new_n1014), .ZN(new_n1015));
  XOR2_X1   g0815(.A(KEYINPUT106), .B(KEYINPUT41), .Z(new_n1016));
  XOR2_X1   g0816(.A(new_n709), .B(new_n1016), .Z(new_n1017));
  OAI21_X1  g0817(.A(KEYINPUT108), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1005), .A2(new_n1008), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1014), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n759), .B(new_n731), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT108), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1017), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1021), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n781), .B1(new_n1018), .B2(new_n1024), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n1011), .A2(new_n1002), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT42), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n522), .B1(new_n986), .B2(new_n681), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1028), .A2(new_n689), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  XOR2_X1   g0830(.A(KEYINPUT105), .B(KEYINPUT43), .Z(new_n1031));
  NAND2_X1  g0831(.A1(new_n982), .A2(new_n1031), .ZN(new_n1032));
  OR2_X1    g0832(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n1030), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT43), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1032), .B1(new_n1035), .B2(new_n982), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1033), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n699), .A2(new_n1002), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1033), .B(new_n1038), .C1(new_n1034), .C2(new_n1036), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NOR3_X1   g0842(.A1(new_n1025), .A2(KEYINPUT109), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT109), .ZN(new_n1044));
  NOR3_X1   g0844(.A1(new_n1015), .A2(KEYINPUT108), .A3(new_n1017), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1022), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n780), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n1042), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1044), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n984), .B1(new_n1043), .B2(new_n1049), .ZN(G387));
  AOI22_X1  g0850(.A1(G303), .A2(new_n788), .B1(new_n790), .B2(G317), .ZN(new_n1051));
  INV_X1    g0851(.A(G322), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n1051), .B1(new_n819), .B2(new_n860), .C1(new_n1052), .C2(new_n794), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT48), .ZN(new_n1054));
  OR2_X1    g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n969), .A2(G294), .B1(new_n965), .B2(new_n851), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1055), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT49), .Z(new_n1059));
  OAI221_X1 g0859(.A(new_n384), .B1(new_n798), .B2(new_n815), .C1(new_n808), .C2(new_n243), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT111), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n785), .A2(new_n413), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(G159), .B2(new_n795), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(new_n362), .B2(new_n860), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n806), .A2(new_n202), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(G50), .A2(new_n790), .B1(new_n788), .B2(G68), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1067), .B(new_n299), .C1(new_n859), .C2(new_n798), .ZN(new_n1068));
  NOR4_X1   g0868(.A1(new_n1065), .A2(new_n974), .A3(new_n1066), .A4(new_n1068), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n766), .B1(new_n1062), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n693), .A2(new_n765), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n774), .A2(new_n712), .B1(new_n479), .B2(new_n708), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n415), .A2(new_n446), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT50), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n256), .B1(new_n225), .B2(new_n202), .ZN(new_n1075));
  NOR3_X1   g0875(.A1(new_n1074), .A2(new_n712), .A3(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n769), .B1(new_n235), .B2(new_n256), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1072), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n833), .B1(new_n1078), .B2(new_n768), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1070), .A2(new_n1071), .A3(new_n1079), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1080), .B(KEYINPUT112), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(new_n781), .B2(new_n1014), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n731), .A2(new_n1014), .A3(new_n759), .ZN(new_n1083));
  XOR2_X1   g0883(.A(new_n709), .B(KEYINPUT113), .Z(new_n1084));
  NAND2_X1  g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1014), .B1(new_n731), .B2(new_n759), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1082), .B1(new_n1085), .B2(new_n1086), .ZN(G393));
  INV_X1    g0887(.A(KEYINPUT114), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1005), .A2(new_n1008), .A3(new_n1088), .ZN(new_n1089));
  NAND4_X1  g0889(.A1(new_n1006), .A2(KEYINPUT114), .A3(new_n699), .A4(new_n1007), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1091), .A2(new_n781), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1002), .A2(new_n765), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n244), .A2(new_n770), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n767), .B1(new_n473), .B2(new_n209), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n782), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  OAI221_X1 g0896(.A(new_n299), .B1(new_n798), .B2(new_n960), .C1(new_n860), .C2(new_n446), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(G77), .B2(new_n965), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n791), .A2(new_n959), .B1(new_n794), .B2(new_n859), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT51), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n415), .A2(new_n788), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(G68), .A2(new_n969), .B1(new_n809), .B2(G87), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n1098), .A2(new_n1100), .A3(new_n1101), .A4(new_n1102), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n806), .A2(new_n850), .B1(new_n808), .B2(new_n479), .ZN(new_n1104));
  OAI221_X1 g0904(.A(new_n384), .B1(new_n798), .B2(new_n1052), .C1(new_n789), .C2(new_n816), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n785), .A2(new_n243), .B1(new_n860), .B2(new_n604), .ZN(new_n1106));
  OR3_X1    g0906(.A1(new_n1104), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n795), .A2(G317), .B1(G311), .B2(new_n790), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1108), .B(KEYINPUT52), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1103), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1096), .B1(new_n766), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1093), .A2(new_n1111), .ZN(new_n1112));
  AND3_X1   g0912(.A1(new_n1089), .A2(new_n1083), .A3(new_n1090), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1084), .B1(new_n1083), .B2(new_n1019), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n1092), .B(new_n1112), .C1(new_n1113), .C2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(KEYINPUT115), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n1091), .A2(new_n781), .B1(new_n1093), .B2(new_n1111), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT115), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1117), .B(new_n1118), .C1(new_n1113), .C2(new_n1114), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1116), .A2(new_n1119), .ZN(G390));
  INV_X1    g0920(.A(new_n1084), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n873), .B1(new_n883), .B2(new_n894), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n908), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n840), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n688), .B1(new_n729), .B2(new_n717), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1124), .B1(new_n1125), .B2(new_n839), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1122), .B1(new_n1123), .B2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n873), .B1(new_n903), .B2(new_n908), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1127), .B1(new_n1128), .B2(new_n919), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n933), .A2(new_n934), .A3(G330), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n908), .A2(new_n758), .A3(G330), .A4(new_n842), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1127), .B(new_n1133), .C1(new_n1128), .C2(new_n919), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n469), .A2(new_n933), .A3(G330), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n646), .B(new_n1136), .C1(new_n731), .C2(new_n647), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n758), .A2(G330), .A3(new_n842), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(new_n1123), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1139), .A2(new_n1130), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n903), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n733), .A2(new_n753), .A3(new_n757), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n932), .A2(new_n930), .ZN(new_n1143));
  OAI211_X1 g0943(.A(G330), .B(new_n842), .C1(new_n1142), .C2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n1123), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1145), .A2(new_n1126), .A3(new_n1133), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1137), .B1(new_n1141), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1121), .B1(new_n1135), .B2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1132), .A2(new_n1147), .A3(new_n1134), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1135), .A2(new_n780), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n917), .A2(new_n763), .A3(new_n918), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n868), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n782), .B1(new_n363), .B2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n384), .B1(new_n798), .B2(new_n816), .ZN(new_n1156));
  INV_X1    g0956(.A(G283), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n860), .A2(new_n479), .B1(new_n794), .B2(new_n1157), .ZN(new_n1158));
  AOI211_X1 g0958(.A(new_n1156), .B(new_n1158), .C1(G97), .C2(new_n788), .ZN(new_n1159));
  OAI221_X1 g0959(.A(new_n1159), .B1(new_n225), .B2(new_n808), .C1(new_n853), .C2(new_n219), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n785), .A2(new_n202), .B1(new_n791), .B2(new_n243), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1161), .B(KEYINPUT116), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n969), .A2(G150), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(new_n1163), .B(KEYINPUT53), .ZN(new_n1164));
  INV_X1    g0964(.A(G128), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n785), .A2(new_n959), .B1(new_n794), .B2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1166), .B1(G137), .B2(new_n802), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n809), .A2(G50), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n384), .B1(new_n799), .B2(G125), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(KEYINPUT54), .B(G143), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(new_n1171), .A2(new_n788), .B1(new_n790), .B2(G132), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n1167), .A2(new_n1168), .A3(new_n1169), .A4(new_n1172), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n1160), .A2(new_n1162), .B1(new_n1164), .B2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1155), .B1(new_n1174), .B2(new_n766), .ZN(new_n1175));
  AND2_X1   g0975(.A1(new_n1153), .A2(new_n1175), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1152), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1151), .A2(new_n1177), .ZN(G378));
  AOI21_X1  g0978(.A(KEYINPUT101), .B1(new_n920), .B2(new_n911), .ZN(new_n1179));
  AND4_X1   g0979(.A1(KEYINPUT101), .A2(new_n902), .A3(new_n911), .A4(new_n913), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(KEYINPUT120), .B(KEYINPUT56), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n645), .A2(KEYINPUT119), .A3(new_n451), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n450), .A2(new_n875), .ZN(new_n1184));
  XOR2_X1   g0984(.A(new_n1184), .B(KEYINPUT55), .Z(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n451), .B1(new_n460), .B2(new_n461), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT119), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1183), .A2(new_n1186), .A3(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1186), .B1(new_n1183), .B2(new_n1189), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1182), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1189), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1185), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1196), .A2(new_n1181), .A3(new_n1190), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1193), .A2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n935), .A2(new_n936), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n937), .A2(new_n938), .ZN(new_n1200));
  AND4_X1   g1000(.A1(G330), .A2(new_n1198), .A3(new_n1199), .A4(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1198), .B1(new_n939), .B2(G330), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n1179), .A2(new_n1180), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1199), .A2(G330), .A3(new_n1200), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1198), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n939), .A2(G330), .A3(new_n1198), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n916), .A2(new_n921), .A3(new_n1206), .A4(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1203), .A2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1198), .A2(new_n763), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n782), .B1(G50), .B2(new_n1154), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n255), .B(new_n384), .C1(new_n806), .C2(new_n202), .ZN(new_n1212));
  OR2_X1    g1012(.A1(new_n1212), .A2(KEYINPUT117), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(KEYINPUT117), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n808), .A2(new_n223), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(G283), .B2(new_n799), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1213), .A2(new_n1214), .A3(new_n1216), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(new_n1217), .B(KEYINPUT118), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n479), .A2(new_n791), .B1(new_n789), .B2(new_n413), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(G68), .B2(new_n965), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n795), .A2(G116), .B1(G97), .B2(new_n802), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1218), .A2(new_n1220), .A3(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT58), .ZN(new_n1223));
  OR2_X1    g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1225));
  AOI21_X1  g1025(.A(G50), .B1(new_n295), .B2(new_n255), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n791), .A2(new_n1165), .B1(new_n789), .B2(new_n858), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(G132), .B2(new_n802), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n965), .A2(G150), .B1(new_n795), .B2(G125), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n1228), .B(new_n1229), .C1(new_n806), .C2(new_n1170), .ZN(new_n1230));
  OR2_X1    g1030(.A1(new_n1230), .A2(KEYINPUT59), .ZN(new_n1231));
  AOI211_X1 g1031(.A(G33), .B(G41), .C1(new_n799), .C2(G124), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1232), .B1(new_n959), .B2(new_n808), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1233), .B1(new_n1230), .B2(KEYINPUT59), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1226), .B1(new_n1231), .B2(new_n1234), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1224), .A2(new_n1225), .A3(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1211), .B1(new_n1236), .B2(new_n766), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n1209), .A2(new_n781), .B1(new_n1210), .B2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1137), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(new_n1203), .A2(new_n1208), .B1(new_n1239), .B2(new_n1150), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1084), .B1(new_n1240), .B2(KEYINPUT57), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1150), .A2(new_n1239), .ZN(new_n1242));
  AND3_X1   g1042(.A1(new_n1209), .A2(KEYINPUT57), .A3(new_n1242), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1238), .B1(new_n1241), .B2(new_n1243), .ZN(G375));
  NAND3_X1  g1044(.A1(new_n1141), .A2(new_n1137), .A3(new_n1146), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(new_n1017), .B(KEYINPUT121), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1148), .A2(new_n1245), .A3(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1141), .A2(new_n1146), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1123), .A2(new_n763), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n782), .B1(G68), .B2(new_n1154), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n384), .B1(new_n789), .B2(new_n479), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n791), .A2(new_n1157), .B1(new_n798), .B2(new_n604), .ZN(new_n1252));
  AOI211_X1 g1052(.A(new_n1251), .B(new_n1252), .C1(G77), .C2(new_n809), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n794), .A2(new_n816), .ZN(new_n1254));
  AOI211_X1 g1054(.A(new_n1254), .B(new_n1063), .C1(G116), .C2(new_n802), .ZN(new_n1255));
  OAI211_X1 g1055(.A(new_n1253), .B(new_n1255), .C1(new_n853), .C2(new_n473), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(new_n822), .A2(G159), .B1(G128), .B2(new_n799), .ZN(new_n1257));
  XNOR2_X1  g1057(.A(new_n1257), .B(KEYINPUT122), .ZN(new_n1258));
  OAI221_X1 g1058(.A(new_n299), .B1(new_n789), .B2(new_n859), .C1(new_n858), .C2(new_n791), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1259), .A2(new_n1215), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(new_n795), .A2(G132), .B1(new_n1171), .B2(new_n802), .ZN(new_n1261));
  OAI211_X1 g1061(.A(new_n1260), .B(new_n1261), .C1(new_n446), .C2(new_n785), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1256), .B1(new_n1258), .B2(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1250), .B1(new_n1263), .B2(new_n766), .ZN(new_n1264));
  AOI22_X1  g1064(.A1(new_n1248), .A2(new_n781), .B1(new_n1249), .B2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1247), .A2(new_n1265), .ZN(G381));
  OR2_X1    g1066(.A1(G375), .A2(G378), .ZN(new_n1267));
  OAI21_X1  g1067(.A(KEYINPUT109), .B1(new_n1025), .B2(new_n1042), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1047), .A2(new_n1044), .A3(new_n1048), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(G390), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1270), .A2(new_n984), .A3(new_n1271), .ZN(new_n1272));
  OR2_X1    g1072(.A1(G393), .A2(G396), .ZN(new_n1273));
  OR2_X1    g1073(.A1(new_n1273), .A2(G384), .ZN(new_n1274));
  OR4_X1    g1074(.A1(G381), .A2(new_n1267), .A3(new_n1272), .A4(new_n1274), .ZN(G407));
  OAI211_X1 g1075(.A(G407), .B(G213), .C1(G343), .C2(new_n1267), .ZN(G409));
  INV_X1    g1076(.A(KEYINPUT61), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n687), .A2(G213), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  OAI211_X1 g1079(.A(G378), .B(new_n1238), .C1(new_n1241), .C2(new_n1243), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1209), .A2(new_n1242), .A3(new_n1246), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1238), .A2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(G378), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1279), .B1(new_n1280), .B2(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1121), .B1(new_n1248), .B2(new_n1239), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT60), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1245), .A2(new_n1287), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1141), .A2(new_n1137), .A3(KEYINPUT60), .A4(new_n1146), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1286), .A2(new_n1288), .A3(new_n1289), .ZN(new_n1290));
  AND3_X1   g1090(.A1(new_n1290), .A2(G384), .A3(new_n1265), .ZN(new_n1291));
  AOI21_X1  g1091(.A(G384), .B1(new_n1290), .B2(new_n1265), .ZN(new_n1292));
  OAI211_X1 g1092(.A(G2897), .B(new_n1279), .C1(new_n1291), .C2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT124), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1295));
  INV_X1    g1095(.A(G2897), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1278), .B1(KEYINPUT123), .B2(new_n1296), .ZN(new_n1297));
  OR2_X1    g1097(.A1(new_n1296), .A2(KEYINPUT123), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1294), .B1(new_n1295), .B2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1299), .ZN(new_n1301));
  NOR4_X1   g1101(.A1(new_n1291), .A2(new_n1292), .A3(KEYINPUT124), .A4(new_n1301), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1293), .B1(new_n1300), .B2(new_n1302), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1277), .B1(new_n1285), .B2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(KEYINPUT127), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT127), .ZN(new_n1306));
  OAI211_X1 g1106(.A(new_n1306), .B(new_n1277), .C1(new_n1285), .C2(new_n1303), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1285), .A2(new_n1295), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1308), .A2(KEYINPUT62), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT62), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1285), .A2(new_n1310), .A3(new_n1295), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1305), .A2(new_n1307), .A3(new_n1309), .A4(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1273), .ZN(new_n1313));
  AND2_X1   g1113(.A1(G393), .A2(G396), .ZN(new_n1314));
  OR3_X1    g1114(.A1(new_n1313), .A2(KEYINPUT125), .A3(new_n1314), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1271), .B1(new_n1270), .B2(new_n984), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n984), .ZN(new_n1317));
  AOI211_X1 g1117(.A(new_n1317), .B(G390), .C1(new_n1268), .C2(new_n1269), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1315), .B1(new_n1316), .B2(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(G387), .A2(G390), .ZN(new_n1320));
  OAI21_X1  g1120(.A(KEYINPUT125), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1315), .A2(new_n1321), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1320), .A2(new_n1272), .A3(new_n1322), .ZN(new_n1323));
  AND2_X1   g1123(.A1(new_n1319), .A2(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1312), .A2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1319), .A2(new_n1323), .ZN(new_n1326));
  OAI211_X1 g1126(.A(new_n1326), .B(new_n1277), .C1(new_n1285), .C2(new_n1303), .ZN(new_n1327));
  AND3_X1   g1127(.A1(new_n1285), .A2(KEYINPUT63), .A3(new_n1295), .ZN(new_n1328));
  AOI21_X1  g1128(.A(KEYINPUT63), .B1(new_n1285), .B2(new_n1295), .ZN(new_n1329));
  NOR4_X1   g1129(.A1(new_n1327), .A2(new_n1328), .A3(KEYINPUT126), .A4(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT126), .ZN(new_n1331));
  NOR2_X1   g1131(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1332));
  NOR2_X1   g1132(.A1(new_n1304), .A2(new_n1324), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1331), .B1(new_n1332), .B2(new_n1333), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1325), .B1(new_n1330), .B2(new_n1334), .ZN(G405));
  NAND2_X1  g1135(.A1(G375), .A2(new_n1283), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1336), .A2(new_n1280), .ZN(new_n1337));
  XNOR2_X1  g1137(.A(new_n1337), .B(new_n1295), .ZN(new_n1338));
  XNOR2_X1  g1138(.A(new_n1338), .B(new_n1324), .ZN(G402));
endmodule


