//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 1 1 0 0 0 0 1 1 1 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 0 0 1 0 1 1 1 1 0 0 0 0 0 0 0 0 1 0 0 1 0 0 1 1 1 0 0 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:42 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n547, new_n549, new_n550, new_n551,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n565, new_n566, new_n567, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n576, new_n577, new_n578,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n591, new_n592, new_n593, new_n596, new_n597,
    new_n599, new_n600, new_n601, new_n602, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n790, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT65), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT66), .ZN(new_n437));
  INV_X1    g012(.A(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n437), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n454), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n454), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  AOI22_X1  g037(.A1(new_n462), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  OR2_X1    g040(.A1(new_n465), .A2(KEYINPUT68), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(KEYINPUT3), .B1(new_n467), .B2(KEYINPUT69), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT69), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n469), .A2(new_n470), .A3(G2104), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n468), .A2(new_n471), .A3(G137), .ZN(new_n472));
  NAND2_X1  g047(.A1(G101), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(G2105), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  OAI21_X1  g049(.A(KEYINPUT68), .B1(new_n465), .B2(new_n474), .ZN(new_n475));
  AND2_X1   g050(.A1(new_n466), .A2(new_n475), .ZN(G160));
  NAND2_X1  g051(.A1(new_n468), .A2(new_n471), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n477), .A2(new_n464), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n477), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n479), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  NAND3_X1  g060(.A1(new_n468), .A2(new_n471), .A3(G126), .ZN(new_n486));
  NAND2_X1  g061(.A1(G114), .A2(G2104), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n464), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n467), .A2(G2105), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G102), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  AND2_X1   g067(.A1(KEYINPUT4), .A2(G138), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n462), .A2(G138), .A3(new_n464), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  AOI22_X1  g070(.A1(new_n480), .A2(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n492), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G164));
  XOR2_X1   g073(.A(KEYINPUT6), .B(G651), .Z(new_n499));
  INV_X1    g074(.A(G543), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT5), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT5), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  OAI21_X1  g079(.A(KEYINPUT70), .B1(new_n499), .B2(new_n504), .ZN(new_n505));
  AND2_X1   g080(.A1(new_n501), .A2(new_n503), .ZN(new_n506));
  XNOR2_X1  g081(.A(KEYINPUT6), .B(G651), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT70), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  AND2_X1   g084(.A1(new_n505), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G88), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n499), .A2(new_n500), .ZN(new_n512));
  NAND2_X1  g087(.A1(G75), .A2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G62), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n513), .B1(new_n504), .B2(new_n514), .ZN(new_n515));
  AOI22_X1  g090(.A1(G50), .A2(new_n512), .B1(new_n515), .B2(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n511), .A2(new_n516), .ZN(G303));
  INV_X1    g092(.A(G303), .ZN(G166));
  NAND2_X1  g093(.A1(new_n510), .A2(G89), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n499), .A2(KEYINPUT71), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT71), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n507), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n520), .A2(G543), .A3(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G51), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n526), .B(KEYINPUT7), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n506), .A2(G63), .A3(G651), .ZN(new_n528));
  NAND4_X1  g103(.A1(new_n519), .A2(new_n525), .A3(new_n527), .A4(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(G168));
  NAND2_X1  g105(.A1(new_n510), .A2(G90), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n524), .A2(G52), .ZN(new_n532));
  INV_X1    g107(.A(G651), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n506), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n534));
  OAI211_X1 g109(.A(new_n531), .B(new_n532), .C1(new_n533), .C2(new_n534), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n535), .B(KEYINPUT72), .ZN(G171));
  NAND2_X1  g111(.A1(new_n505), .A2(new_n509), .ZN(new_n537));
  INV_X1    g112(.A(G81), .ZN(new_n538));
  INV_X1    g113(.A(G43), .ZN(new_n539));
  OAI22_X1  g114(.A1(new_n537), .A2(new_n538), .B1(new_n523), .B2(new_n539), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT73), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n506), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n542), .A2(new_n533), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G860), .ZN(G153));
  AND3_X1   g121(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G36), .ZN(G176));
  XOR2_X1   g123(.A(KEYINPUT74), .B(KEYINPUT8), .Z(new_n549));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n549), .B(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n547), .A2(new_n551), .ZN(G188));
  INV_X1    g127(.A(KEYINPUT9), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n553), .A2(KEYINPUT75), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n524), .A2(G53), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n510), .A2(G91), .ZN(new_n556));
  INV_X1    g131(.A(G53), .ZN(new_n557));
  OAI22_X1  g132(.A1(new_n523), .A2(new_n557), .B1(KEYINPUT75), .B2(new_n553), .ZN(new_n558));
  AND3_X1   g133(.A1(new_n555), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n506), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n560));
  OR2_X1    g135(.A1(new_n560), .A2(new_n533), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n559), .A2(new_n561), .ZN(G299));
  INV_X1    g137(.A(G171), .ZN(G301));
  XNOR2_X1  g138(.A(new_n529), .B(KEYINPUT76), .ZN(G286));
  NAND2_X1  g139(.A1(new_n510), .A2(G87), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n524), .A2(G49), .ZN(new_n566));
  OAI21_X1  g141(.A(G651), .B1(new_n506), .B2(G74), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(G288));
  NAND2_X1  g143(.A1(new_n510), .A2(G86), .ZN(new_n569));
  NAND2_X1  g144(.A1(G73), .A2(G543), .ZN(new_n570));
  INV_X1    g145(.A(G61), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n504), .B2(new_n571), .ZN(new_n572));
  AOI22_X1  g147(.A1(G48), .A2(new_n512), .B1(new_n572), .B2(G651), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n569), .A2(new_n573), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n574), .B(KEYINPUT77), .ZN(G305));
  NAND2_X1  g150(.A1(new_n510), .A2(G85), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n506), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n577));
  XOR2_X1   g152(.A(KEYINPUT78), .B(G47), .Z(new_n578));
  OAI221_X1 g153(.A(new_n576), .B1(new_n533), .B2(new_n577), .C1(new_n523), .C2(new_n578), .ZN(G290));
  NAND2_X1  g154(.A1(new_n510), .A2(G92), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n580), .B(KEYINPUT10), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n506), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n582), .A2(new_n533), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n524), .A2(G54), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(G868), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n588), .B1(new_n587), .B2(G171), .ZN(G284));
  OAI21_X1  g164(.A(new_n588), .B1(new_n587), .B2(G171), .ZN(G321));
  NAND2_X1  g165(.A1(G286), .A2(G868), .ZN(new_n591));
  XOR2_X1   g166(.A(new_n591), .B(KEYINPUT79), .Z(new_n592));
  INV_X1    g167(.A(G299), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(G868), .B2(new_n593), .ZN(G297));
  OAI21_X1  g169(.A(new_n592), .B1(G868), .B2(new_n593), .ZN(G280));
  INV_X1    g170(.A(new_n586), .ZN(new_n596));
  INV_X1    g171(.A(G559), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n597), .B2(G860), .ZN(G148));
  NAND2_X1  g173(.A1(new_n596), .A2(new_n597), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n599), .A2(G868), .ZN(new_n600));
  OR2_X1    g175(.A1(new_n600), .A2(KEYINPUT80), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(KEYINPUT80), .ZN(new_n602));
  OAI211_X1 g177(.A(new_n601), .B(new_n602), .C1(G868), .C2(new_n545), .ZN(G323));
  XNOR2_X1  g178(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g179(.A1(new_n462), .A2(new_n489), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n605), .B(KEYINPUT12), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(G2100), .ZN(new_n607));
  XNOR2_X1  g182(.A(KEYINPUT81), .B(KEYINPUT13), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n607), .B(new_n608), .ZN(new_n609));
  AOI22_X1  g184(.A1(G123), .A2(new_n478), .B1(new_n480), .B2(G135), .ZN(new_n610));
  OAI21_X1  g185(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT82), .ZN(new_n612));
  OR2_X1    g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n611), .A2(new_n612), .ZN(new_n614));
  OAI211_X1 g189(.A(new_n613), .B(new_n614), .C1(G111), .C2(new_n464), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n610), .A2(new_n615), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(G2096), .Z(new_n617));
  NAND2_X1  g192(.A1(new_n609), .A2(new_n617), .ZN(G156));
  XNOR2_X1  g193(.A(G2451), .B(G2454), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT16), .ZN(new_n620));
  XOR2_X1   g195(.A(G2443), .B(G2446), .Z(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XNOR2_X1  g197(.A(G1341), .B(G1348), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XNOR2_X1  g199(.A(G2427), .B(G2438), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(G2430), .ZN(new_n626));
  XOR2_X1   g201(.A(KEYINPUT15), .B(G2435), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(KEYINPUT14), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n624), .B(new_n629), .ZN(new_n630));
  AND2_X1   g205(.A1(new_n630), .A2(G14), .ZN(G401));
  XOR2_X1   g206(.A(G2084), .B(G2090), .Z(new_n632));
  INV_X1    g207(.A(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(G2067), .B(G2678), .Z(new_n634));
  NOR2_X1   g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g210(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n633), .A2(new_n634), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n636), .A2(new_n637), .A3(KEYINPUT17), .ZN(new_n638));
  INV_X1    g213(.A(KEYINPUT18), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2072), .B(G2078), .ZN(new_n641));
  OAI211_X1 g216(.A(new_n640), .B(new_n641), .C1(new_n639), .C2(new_n635), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n642), .B1(new_n641), .B2(new_n640), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2096), .B(G2100), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(G227));
  XNOR2_X1  g220(.A(G1971), .B(G1976), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT19), .ZN(new_n647));
  XOR2_X1   g222(.A(G1956), .B(G2474), .Z(new_n648));
  XOR2_X1   g223(.A(G1961), .B(G1966), .Z(new_n649));
  NAND2_X1  g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(new_n647), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n648), .A2(new_n649), .ZN(new_n653));
  AOI22_X1  g228(.A1(new_n651), .A2(KEYINPUT20), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n653), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n655), .A2(new_n647), .A3(new_n650), .ZN(new_n656));
  OAI211_X1 g231(.A(new_n654), .B(new_n656), .C1(KEYINPUT20), .C2(new_n651), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1986), .B(G1996), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G1981), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(G1991), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n659), .B(new_n662), .ZN(G229));
  XNOR2_X1  g238(.A(KEYINPUT31), .B(G11), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT91), .ZN(new_n665));
  INV_X1    g240(.A(G28), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n666), .A2(KEYINPUT30), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(KEYINPUT30), .ZN(new_n668));
  INV_X1    g243(.A(G29), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  OAI211_X1 g245(.A(new_n665), .B(new_n670), .C1(new_n616), .C2(new_n669), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(KEYINPUT92), .Z(new_n672));
  INV_X1    g247(.A(KEYINPUT24), .ZN(new_n673));
  AND2_X1   g248(.A1(new_n673), .A2(G34), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n673), .A2(G34), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n669), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n676), .B1(G160), .B2(new_n669), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n677), .A2(G2084), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT95), .ZN(new_n679));
  OR2_X1    g254(.A1(G29), .A2(G32), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n478), .A2(G129), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT88), .ZN(new_n682));
  NAND3_X1  g257(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(KEYINPUT26), .Z(new_n684));
  AOI22_X1  g259(.A1(new_n480), .A2(G141), .B1(G105), .B2(new_n489), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n682), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n680), .B1(new_n686), .B2(new_n669), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT27), .B(G1996), .ZN(new_n688));
  NOR2_X1   g263(.A1(G5), .A2(G16), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n689), .B1(G171), .B2(G16), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT93), .ZN(new_n691));
  OAI221_X1 g266(.A(new_n679), .B1(new_n687), .B2(new_n688), .C1(new_n691), .C2(G1961), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n692), .B(KEYINPUT96), .Z(new_n693));
  NAND2_X1  g268(.A1(new_n691), .A2(G1961), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n694), .B(KEYINPUT94), .Z(new_n695));
  INV_X1    g270(.A(G16), .ZN(new_n696));
  OAI21_X1  g271(.A(KEYINPUT23), .B1(new_n593), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n696), .A2(G20), .ZN(new_n698));
  MUX2_X1   g273(.A(KEYINPUT23), .B(new_n697), .S(new_n698), .Z(new_n699));
  OR2_X1    g274(.A1(new_n699), .A2(G1956), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n687), .A2(new_n688), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT89), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n699), .A2(G1956), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n696), .A2(G4), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(new_n596), .B2(new_n696), .ZN(new_n705));
  OR2_X1    g280(.A1(new_n705), .A2(G1348), .ZN(new_n706));
  NAND4_X1  g281(.A1(new_n700), .A2(new_n702), .A3(new_n703), .A4(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n696), .A2(G19), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(new_n545), .B2(new_n696), .ZN(new_n709));
  INV_X1    g284(.A(KEYINPUT28), .ZN(new_n710));
  INV_X1    g285(.A(G26), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n710), .B1(new_n711), .B2(G29), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n711), .A2(G29), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n478), .A2(G128), .ZN(new_n714));
  INV_X1    g289(.A(KEYINPUT87), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  OR2_X1    g291(.A1(G104), .A2(G2105), .ZN(new_n717));
  OAI211_X1 g292(.A(new_n717), .B(G2104), .C1(G116), .C2(new_n464), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n480), .A2(G140), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n716), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n713), .B1(new_n720), .B2(G29), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n712), .B1(new_n721), .B2(new_n710), .ZN(new_n722));
  AOI22_X1  g297(.A1(new_n709), .A2(G1341), .B1(G2067), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n669), .A2(G27), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(G164), .B2(new_n669), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT97), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(G2078), .ZN(new_n727));
  OAI211_X1 g302(.A(new_n723), .B(new_n727), .C1(G2067), .C2(new_n722), .ZN(new_n728));
  NOR2_X1   g303(.A1(G168), .A2(new_n696), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(new_n696), .B2(G21), .ZN(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT90), .B(G1966), .ZN(new_n731));
  INV_X1    g306(.A(G2072), .ZN(new_n732));
  AND2_X1   g307(.A1(new_n669), .A2(G33), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n489), .A2(G103), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT25), .Z(new_n735));
  NAND2_X1  g310(.A1(new_n480), .A2(G139), .ZN(new_n736));
  AOI22_X1  g311(.A1(new_n462), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n737));
  OAI211_X1 g312(.A(new_n735), .B(new_n736), .C1(new_n464), .C2(new_n737), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n733), .B1(new_n738), .B2(G29), .ZN(new_n739));
  OAI22_X1  g314(.A1(new_n730), .A2(new_n731), .B1(new_n732), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n669), .A2(G35), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G162), .B2(new_n669), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT29), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n740), .B1(G2090), .B2(new_n743), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n743), .A2(G2090), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(new_n705), .B2(G1348), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n739), .A2(new_n732), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n744), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n730), .A2(new_n731), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n677), .A2(G2084), .ZN(new_n750));
  OAI211_X1 g325(.A(new_n749), .B(new_n750), .C1(G1341), .C2(new_n709), .ZN(new_n751));
  NOR4_X1   g326(.A1(new_n707), .A2(new_n728), .A3(new_n748), .A4(new_n751), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n693), .A2(new_n695), .A3(new_n752), .ZN(new_n753));
  MUX2_X1   g328(.A(G6), .B(G305), .S(G16), .Z(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT84), .ZN(new_n755));
  XOR2_X1   g330(.A(KEYINPUT32), .B(G1981), .Z(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(G166), .A2(new_n696), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(new_n696), .B2(G22), .ZN(new_n759));
  INV_X1    g334(.A(G1971), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT85), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G16), .B2(G23), .ZN(new_n763));
  OR3_X1    g338(.A1(new_n762), .A2(G16), .A3(G23), .ZN(new_n764));
  XOR2_X1   g339(.A(G288), .B(KEYINPUT86), .Z(new_n765));
  OAI211_X1 g340(.A(new_n763), .B(new_n764), .C1(new_n765), .C2(new_n696), .ZN(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT33), .B(G1976), .ZN(new_n767));
  OAI22_X1  g342(.A1(new_n766), .A2(new_n767), .B1(new_n760), .B2(new_n759), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(new_n767), .B2(new_n766), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n757), .A2(new_n761), .A3(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n770), .A2(KEYINPUT34), .ZN(new_n771));
  MUX2_X1   g346(.A(G24), .B(G290), .S(G16), .Z(new_n772));
  OR2_X1    g347(.A1(new_n772), .A2(G1986), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT34), .ZN(new_n774));
  NAND4_X1  g349(.A1(new_n757), .A2(new_n774), .A3(new_n761), .A4(new_n769), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n480), .A2(G131), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT83), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n478), .A2(G119), .ZN(new_n778));
  NOR2_X1   g353(.A1(G95), .A2(G2105), .ZN(new_n779));
  OAI21_X1  g354(.A(G2104), .B1(new_n464), .B2(G107), .ZN(new_n780));
  OAI211_X1 g355(.A(new_n777), .B(new_n778), .C1(new_n779), .C2(new_n780), .ZN(new_n781));
  MUX2_X1   g356(.A(G25), .B(new_n781), .S(G29), .Z(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT35), .B(G1991), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(G1986), .B2(new_n772), .ZN(new_n785));
  NAND4_X1  g360(.A1(new_n771), .A2(new_n773), .A3(new_n775), .A4(new_n785), .ZN(new_n786));
  OR2_X1    g361(.A1(new_n786), .A2(KEYINPUT36), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n786), .A2(KEYINPUT36), .ZN(new_n788));
  AOI211_X1 g363(.A(new_n672), .B(new_n753), .C1(new_n787), .C2(new_n788), .ZN(G311));
  AOI21_X1  g364(.A(new_n753), .B1(new_n787), .B2(new_n788), .ZN(new_n790));
  INV_X1    g365(.A(new_n672), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n790), .A2(new_n791), .ZN(G150));
  AND2_X1   g367(.A1(new_n510), .A2(G93), .ZN(new_n793));
  INV_X1    g368(.A(G55), .ZN(new_n794));
  AOI22_X1  g369(.A1(new_n506), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n795));
  OAI22_X1  g370(.A1(new_n523), .A2(new_n794), .B1(new_n533), .B2(new_n795), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n798), .A2(G860), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT37), .Z(new_n800));
  NOR2_X1   g375(.A1(new_n586), .A2(new_n597), .ZN(new_n801));
  XNOR2_X1  g376(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT39), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n801), .B(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(KEYINPUT99), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n797), .B1(new_n544), .B2(new_n805), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(new_n805), .B2(new_n544), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n545), .A2(KEYINPUT99), .A3(new_n797), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n804), .B(new_n809), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n800), .B1(new_n810), .B2(G860), .ZN(G145));
  NAND2_X1  g386(.A1(new_n478), .A2(G130), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n480), .A2(G142), .ZN(new_n813));
  NOR2_X1   g388(.A1(G106), .A2(G2105), .ZN(new_n814));
  OAI21_X1  g389(.A(G2104), .B1(new_n464), .B2(G118), .ZN(new_n815));
  OAI211_X1 g390(.A(new_n812), .B(new_n813), .C1(new_n814), .C2(new_n815), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n686), .B(new_n816), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT100), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n486), .A2(new_n487), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n820), .A2(G2105), .ZN(new_n821));
  AOI21_X1  g396(.A(KEYINPUT101), .B1(new_n821), .B2(new_n490), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT101), .ZN(new_n823));
  NOR3_X1   g398(.A1(new_n488), .A2(new_n823), .A3(new_n491), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n496), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n720), .B(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(new_n781), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n738), .B(new_n606), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(new_n484), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n829), .A2(new_n484), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n819), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(new_n832), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n834), .A2(new_n818), .A3(new_n830), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  XOR2_X1   g411(.A(G160), .B(new_n616), .Z(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(G37), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n833), .A2(new_n835), .A3(new_n837), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n839), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g418(.A1(new_n596), .A2(new_n593), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n586), .A2(G299), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(KEYINPUT41), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT41), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n844), .A2(new_n848), .A3(new_n845), .ZN(new_n849));
  AND2_X1   g424(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n809), .B(new_n599), .ZN(new_n851));
  MUX2_X1   g426(.A(new_n850), .B(new_n846), .S(new_n851), .Z(new_n852));
  OR2_X1    g427(.A1(new_n852), .A2(KEYINPUT42), .ZN(new_n853));
  XNOR2_X1  g428(.A(G290), .B(G166), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(G305), .ZN(new_n855));
  INV_X1    g430(.A(new_n765), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n855), .B(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n852), .A2(KEYINPUT42), .ZN(new_n859));
  AND3_X1   g434(.A1(new_n853), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n858), .B1(new_n853), .B2(new_n859), .ZN(new_n861));
  OAI21_X1  g436(.A(G868), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n798), .A2(new_n587), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(G295));
  NAND2_X1  g439(.A1(new_n862), .A2(new_n863), .ZN(G331));
  INV_X1    g440(.A(KEYINPUT44), .ZN(new_n866));
  NAND2_X1  g441(.A1(G171), .A2(G286), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT103), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n867), .B(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(G301), .A2(G168), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(new_n809), .ZN(new_n872));
  NAND4_X1  g447(.A1(new_n869), .A2(new_n808), .A3(new_n807), .A4(new_n870), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n846), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n872), .A2(new_n873), .ZN(new_n876));
  OAI211_X1 g451(.A(new_n875), .B(new_n857), .C1(new_n850), .C2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT105), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n847), .A2(new_n849), .A3(new_n878), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n846), .A2(KEYINPUT105), .A3(KEYINPUT41), .ZN(new_n880));
  AND4_X1   g455(.A1(new_n873), .A2(new_n872), .A3(new_n879), .A4(new_n880), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n858), .B1(new_n881), .B2(new_n874), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n877), .A2(new_n882), .A3(new_n840), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(KEYINPUT43), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n857), .A2(KEYINPUT104), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  OAI211_X1 g461(.A(new_n875), .B(new_n886), .C1(new_n850), .C2(new_n876), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n876), .A2(new_n850), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n885), .B1(new_n888), .B2(new_n874), .ZN(new_n889));
  XOR2_X1   g464(.A(KEYINPUT102), .B(KEYINPUT43), .Z(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  NAND4_X1  g466(.A1(new_n887), .A2(new_n889), .A3(new_n840), .A4(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n866), .B1(new_n884), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n887), .A2(new_n889), .A3(new_n840), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(new_n890), .ZN(new_n895));
  NAND4_X1  g470(.A1(new_n877), .A2(new_n882), .A3(new_n840), .A4(new_n891), .ZN(new_n896));
  AND2_X1   g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n893), .B1(new_n866), .B2(new_n897), .ZN(G397));
  NAND3_X1  g473(.A1(new_n821), .A2(KEYINPUT101), .A3(new_n490), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n823), .B1(new_n488), .B2(new_n491), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(G1384), .B1(new_n901), .B2(new_n496), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n902), .A2(KEYINPUT45), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n466), .A2(G40), .A3(new_n475), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NOR3_X1   g481(.A1(new_n906), .A2(G1996), .A3(new_n686), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n906), .B(KEYINPUT106), .ZN(new_n908));
  INV_X1    g483(.A(G2067), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n720), .B(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n686), .A2(G1996), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n907), .B1(new_n908), .B2(new_n912), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n781), .A2(new_n783), .ZN(new_n914));
  AND2_X1   g489(.A1(new_n781), .A2(new_n783), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n908), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n913), .A2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n906), .ZN(new_n918));
  XNOR2_X1  g493(.A(G290), .B(G1986), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n917), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(G40), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n903), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(G1384), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n497), .A2(KEYINPUT45), .A3(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n922), .A2(G160), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(new_n731), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n497), .A2(new_n923), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(KEYINPUT50), .ZN(new_n928));
  XOR2_X1   g503(.A(new_n928), .B(KEYINPUT107), .Z(new_n929));
  INV_X1    g504(.A(KEYINPUT50), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n902), .A2(new_n930), .ZN(new_n931));
  XNOR2_X1  g506(.A(KEYINPUT115), .B(G2084), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n929), .A2(new_n905), .A3(new_n931), .A4(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n926), .A2(new_n933), .A3(KEYINPUT124), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(KEYINPUT124), .B1(new_n926), .B2(new_n933), .ZN(new_n936));
  OAI211_X1 g511(.A(G8), .B(new_n529), .C1(new_n935), .C2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT51), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n926), .A2(new_n933), .ZN(new_n939));
  OAI211_X1 g514(.A(new_n938), .B(G8), .C1(new_n939), .C2(new_n529), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n937), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n936), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n943), .A2(G168), .A3(new_n934), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(G8), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(KEYINPUT51), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n942), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n574), .A2(G1981), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT108), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n950), .B1(new_n574), .B2(G1981), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(new_n574), .ZN(new_n953));
  INV_X1    g528(.A(G1981), .ZN(new_n954));
  NOR3_X1   g529(.A1(new_n953), .A2(new_n950), .A3(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT49), .B1(new_n952), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n905), .A2(new_n902), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(G8), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  OAI21_X1  g534(.A(KEYINPUT109), .B1(new_n952), .B2(new_n955), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n953), .A2(new_n954), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n961), .A2(new_n950), .A3(new_n948), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n949), .A2(new_n951), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT109), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n962), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n960), .A2(new_n965), .ZN(new_n966));
  XOR2_X1   g541(.A(KEYINPUT110), .B(KEYINPUT49), .Z(new_n967));
  AOI21_X1  g542(.A(KEYINPUT111), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT111), .ZN(new_n969));
  INV_X1    g544(.A(new_n967), .ZN(new_n970));
  AOI211_X1 g545(.A(new_n969), .B(new_n970), .C1(new_n960), .C2(new_n965), .ZN(new_n971));
  OAI211_X1 g546(.A(new_n956), .B(new_n959), .C1(new_n968), .C2(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n958), .B1(new_n856), .B2(G1976), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT52), .ZN(new_n974));
  OR2_X1    g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(G288), .ZN(new_n976));
  OAI211_X1 g551(.A(new_n973), .B(new_n974), .C1(G1976), .C2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n972), .A2(new_n975), .A3(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(G8), .ZN(new_n979));
  INV_X1    g554(.A(G2090), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n929), .A2(new_n980), .A3(new_n905), .A4(new_n931), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n902), .A2(KEYINPUT45), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT45), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n927), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n982), .A2(new_n905), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(new_n760), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n979), .B1(new_n981), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(G303), .A2(G8), .ZN(new_n988));
  XOR2_X1   g563(.A(new_n988), .B(KEYINPUT55), .Z(new_n989));
  AND2_X1   g564(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n930), .B1(new_n825), .B2(new_n923), .ZN(new_n991));
  OAI21_X1  g566(.A(KEYINPUT113), .B1(new_n991), .B2(new_n904), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n497), .A2(new_n930), .A3(new_n923), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT114), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n993), .B(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT113), .ZN(new_n996));
  OAI211_X1 g571(.A(new_n905), .B(new_n996), .C1(new_n902), .C2(new_n930), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n992), .A2(new_n995), .A3(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n986), .B1(new_n998), .B2(G2090), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n989), .B1(new_n999), .B2(G8), .ZN(new_n1000));
  NOR3_X1   g575(.A1(new_n978), .A2(new_n990), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT54), .ZN(new_n1002));
  AND3_X1   g577(.A1(new_n982), .A2(new_n905), .A3(new_n984), .ZN(new_n1003));
  INV_X1    g578(.A(G2078), .ZN(new_n1004));
  AOI21_X1  g579(.A(KEYINPUT53), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(G1961), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n929), .A2(new_n905), .A3(new_n931), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1005), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1004), .A2(KEYINPUT53), .ZN(new_n1009));
  OR2_X1    g584(.A1(new_n925), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1008), .A2(G301), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT126), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n465), .A2(new_n474), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n922), .A2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1009), .B1(new_n1015), .B2(KEYINPUT125), .ZN(new_n1016));
  OAI211_X1 g591(.A(new_n1016), .B(new_n982), .C1(KEYINPUT125), .C2(new_n1015), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(new_n1008), .ZN(new_n1018));
  AOI21_X1  g593(.A(KEYINPUT126), .B1(new_n1018), .B2(G171), .ZN(new_n1019));
  AOI211_X1 g594(.A(new_n1002), .B(new_n1013), .C1(new_n1019), .C2(new_n1011), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1018), .A2(G171), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(G171), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1023), .ZN(new_n1024));
  NOR3_X1   g599(.A1(new_n1021), .A2(new_n1024), .A3(KEYINPUT54), .ZN(new_n1025));
  OAI211_X1 g600(.A(new_n947), .B(new_n1001), .C1(new_n1020), .C2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(G1956), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n998), .A2(new_n1027), .ZN(new_n1028));
  XNOR2_X1  g603(.A(KEYINPUT56), .B(G2072), .ZN(new_n1029));
  XNOR2_X1  g604(.A(new_n1029), .B(KEYINPUT117), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1003), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1028), .A2(new_n1031), .ZN(new_n1032));
  XOR2_X1   g607(.A(G299), .B(KEYINPUT57), .Z(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1028), .A2(new_n1033), .A3(new_n1031), .ZN(new_n1036));
  AND2_X1   g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(G1996), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1003), .A2(KEYINPUT119), .A3(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT119), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1040), .B1(new_n985), .B2(G1996), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(new_n957), .ZN(new_n1043));
  XNOR2_X1  g618(.A(KEYINPUT58), .B(G1341), .ZN(new_n1044));
  OAI21_X1  g619(.A(KEYINPUT120), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT120), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1044), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n957), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1042), .A2(new_n1045), .A3(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT121), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT59), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .A4(new_n545), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1045), .A2(new_n1048), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1053), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n545), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1055));
  OAI22_X1  g630(.A1(new_n1054), .A2(new_n1055), .B1(KEYINPUT121), .B2(KEYINPUT59), .ZN(new_n1056));
  AOI22_X1  g631(.A1(new_n1037), .A2(KEYINPUT61), .B1(new_n1052), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT118), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1036), .A2(new_n1058), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1028), .A2(new_n1033), .A3(KEYINPUT118), .A4(new_n1031), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1059), .A2(new_n1035), .A3(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT122), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT61), .ZN(new_n1063));
  AND3_X1   g638(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1062), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1057), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(KEYINPUT123), .ZN(new_n1067));
  INV_X1    g642(.A(G1348), .ZN(new_n1068));
  AOI22_X1  g643(.A1(new_n1007), .A2(new_n1068), .B1(new_n909), .B2(new_n1043), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(KEYINPUT60), .ZN(new_n1070));
  XNOR2_X1  g645(.A(new_n1070), .B(new_n596), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1071), .B1(KEYINPUT60), .B2(new_n1069), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT123), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1057), .B(new_n1073), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1067), .A2(new_n1072), .A3(new_n1074), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1035), .B1(new_n586), .B2(new_n1069), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1076), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1026), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT62), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n942), .A2(new_n946), .A3(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n938), .B1(new_n944), .B2(G8), .ZN(new_n1081));
  OAI21_X1  g656(.A(KEYINPUT62), .B1(new_n1081), .B2(new_n941), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1080), .A2(new_n1082), .A3(new_n1024), .A4(new_n1001), .ZN(new_n1083));
  INV_X1    g658(.A(G286), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n939), .A2(G8), .A3(new_n1084), .ZN(new_n1085));
  NOR4_X1   g660(.A1(new_n978), .A2(new_n1085), .A3(new_n990), .A4(new_n1000), .ZN(new_n1086));
  INV_X1    g661(.A(new_n978), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT116), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n989), .A2(new_n1088), .ZN(new_n1089));
  XNOR2_X1  g664(.A(new_n987), .B(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1087), .A2(new_n1090), .A3(KEYINPUT63), .ZN(new_n1091));
  OAI22_X1  g666(.A1(new_n1086), .A2(KEYINPUT63), .B1(new_n1091), .B2(new_n1085), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1087), .A2(new_n990), .ZN(new_n1093));
  INV_X1    g668(.A(G1976), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n972), .A2(new_n1094), .A3(new_n976), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(new_n961), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(KEYINPUT112), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT112), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1095), .A2(new_n1098), .A3(new_n961), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1097), .A2(new_n959), .A3(new_n1099), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1083), .A2(new_n1092), .A3(new_n1093), .A4(new_n1100), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n920), .B1(new_n1078), .B2(new_n1101), .ZN(new_n1102));
  NOR3_X1   g677(.A1(new_n906), .A2(G1986), .A3(G290), .ZN(new_n1103));
  XOR2_X1   g678(.A(new_n1103), .B(KEYINPUT127), .Z(new_n1104));
  XNOR2_X1  g679(.A(new_n1104), .B(KEYINPUT48), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1105), .A2(new_n913), .A3(new_n916), .ZN(new_n1106));
  AND2_X1   g681(.A1(new_n913), .A2(new_n914), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n720), .A2(G2067), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n908), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n906), .A2(G1996), .ZN(new_n1110));
  XOR2_X1   g685(.A(new_n1110), .B(KEYINPUT46), .Z(new_n1111));
  INV_X1    g686(.A(new_n910), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n908), .B1(new_n686), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1114));
  XNOR2_X1  g689(.A(new_n1114), .B(KEYINPUT47), .ZN(new_n1115));
  AND3_X1   g690(.A1(new_n1106), .A2(new_n1109), .A3(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1102), .A2(new_n1116), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g692(.A1(G401), .A2(G227), .ZN(new_n1119));
  AND2_X1   g693(.A1(new_n842), .A2(new_n1119), .ZN(new_n1120));
  NOR2_X1   g694(.A1(G229), .A2(new_n460), .ZN(new_n1121));
  INV_X1    g695(.A(new_n1121), .ZN(new_n1122));
  AOI21_X1  g696(.A(new_n1122), .B1(new_n895), .B2(new_n896), .ZN(new_n1123));
  AND2_X1   g697(.A1(new_n1120), .A2(new_n1123), .ZN(G308));
  NAND2_X1  g698(.A1(new_n1120), .A2(new_n1123), .ZN(G225));
endmodule


