//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 0 1 1 1 0 1 1 0 1 0 0 0 1 1 1 1 0 0 0 0 0 0 0 1 0 0 1 1 1 1 1 0 1 0 1 0 0 0 1 0 0 1 0 0 1 1 1 0 0 1 1 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:58 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1282, new_n1283, new_n1284, new_n1285,
    new_n1286, new_n1287, new_n1288, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NOR2_X1   g0002(.A1(G58), .A2(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  INV_X1    g0004(.A(new_n204), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(new_n203), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G50), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT65), .Z(new_n209));
  AND2_X1   g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  NAND3_X1  g0010(.A1(new_n209), .A2(G20), .A3(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(KEYINPUT0), .ZN(new_n212));
  INV_X1    g0012(.A(G1), .ZN(new_n213));
  INV_X1    g0013(.A(G20), .ZN(new_n214));
  NOR3_X1   g0014(.A1(new_n213), .A2(new_n214), .A3(G13), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  OAI21_X1  g0016(.A(new_n211), .B1(new_n212), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G116), .A2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G244), .ZN(new_n219));
  INV_X1    g0019(.A(G87), .ZN(new_n220));
  INV_X1    g0020(.A(G250), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n218), .B1(new_n202), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n223));
  INV_X1    g0023(.A(G50), .ZN(new_n224));
  INV_X1    g0024(.A(G226), .ZN(new_n225));
  INV_X1    g0025(.A(G68), .ZN(new_n226));
  INV_X1    g0026(.A(G238), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n223), .B1(new_n224), .B2(new_n225), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  AOI211_X1 g0028(.A(new_n222), .B(new_n228), .C1(G97), .C2(G257), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(G1), .B2(G20), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n230), .B(KEYINPUT1), .Z(new_n231));
  AOI211_X1 g0031(.A(new_n217), .B(new_n231), .C1(new_n212), .C2(new_n216), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT66), .B(G264), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n236), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G58), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  INV_X1    g0048(.A(G1698), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n225), .A2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G232), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G1698), .ZN(new_n252));
  AND2_X1   g0052(.A1(KEYINPUT3), .A2(G33), .ZN(new_n253));
  NOR2_X1   g0053(.A1(KEYINPUT3), .A2(G33), .ZN(new_n254));
  OAI211_X1 g0054(.A(new_n250), .B(new_n252), .C1(new_n253), .C2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(G33), .A2(G97), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(G33), .A2(G41), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n210), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  AND2_X1   g0061(.A1(G33), .A2(G41), .ZN(new_n262));
  NAND2_X1  g0062(.A1(G1), .A2(G13), .ZN(new_n263));
  OAI21_X1  g0063(.A(KEYINPUT67), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT67), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n210), .A2(new_n265), .A3(new_n258), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G41), .ZN(new_n268));
  INV_X1    g0068(.A(G45), .ZN(new_n269));
  AOI21_X1  g0069(.A(G1), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n267), .A2(G238), .A3(new_n271), .ZN(new_n272));
  NOR3_X1   g0072(.A1(new_n262), .A2(KEYINPUT67), .A3(new_n263), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n265), .B1(new_n210), .B2(new_n258), .ZN(new_n274));
  OAI211_X1 g0074(.A(G274), .B(new_n270), .C1(new_n273), .C2(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n261), .A2(new_n272), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(KEYINPUT13), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT76), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT13), .ZN(new_n279));
  NAND4_X1  g0079(.A1(new_n261), .A2(new_n272), .A3(new_n279), .A4(new_n275), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n277), .A2(new_n278), .A3(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n276), .A2(KEYINPUT76), .A3(KEYINPUT13), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G179), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(KEYINPUT79), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n277), .A2(KEYINPUT75), .A3(new_n280), .ZN(new_n286));
  OR3_X1    g0086(.A1(new_n276), .A2(KEYINPUT75), .A3(KEYINPUT13), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n286), .A2(new_n287), .A3(G169), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(KEYINPUT14), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT14), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n286), .A2(new_n287), .A3(new_n290), .A4(G169), .ZN(new_n291));
  INV_X1    g0091(.A(G179), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n292), .B1(new_n281), .B2(new_n282), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT79), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n285), .A2(new_n289), .A3(new_n291), .A4(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G33), .ZN(new_n297));
  OAI21_X1  g0097(.A(KEYINPUT68), .B1(new_n297), .B2(G20), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT68), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n299), .A2(new_n214), .A3(G33), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  OAI22_X1  g0101(.A1(new_n301), .A2(new_n202), .B1(new_n214), .B2(G68), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(KEYINPUT77), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT77), .ZN(new_n304));
  OAI221_X1 g0104(.A(new_n304), .B1(new_n214), .B2(G68), .C1(new_n301), .C2(new_n202), .ZN(new_n305));
  NOR2_X1   g0105(.A1(G20), .A2(G33), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G50), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n303), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(new_n263), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n308), .A2(KEYINPUT11), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n310), .B1(new_n213), .B2(G20), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(G68), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G13), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n315), .A2(G1), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n316), .A2(G20), .A3(new_n226), .ZN(new_n317));
  XOR2_X1   g0117(.A(new_n317), .B(KEYINPUT12), .Z(new_n318));
  AOI21_X1  g0118(.A(KEYINPUT11), .B1(new_n308), .B2(new_n310), .ZN(new_n319));
  NOR3_X1   g0119(.A1(new_n314), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n296), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n283), .A2(G190), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n286), .A2(new_n287), .A3(G200), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n320), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT78), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n320), .A2(new_n323), .A3(KEYINPUT78), .A4(new_n324), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n322), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT82), .ZN(new_n331));
  INV_X1    g0131(.A(G169), .ZN(new_n332));
  OAI211_X1 g0132(.A(G232), .B(new_n271), .C1(new_n273), .C2(new_n274), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n275), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(G223), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(new_n249), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n225), .A2(G1698), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n336), .B(new_n337), .C1(new_n253), .C2(new_n254), .ZN(new_n338));
  NAND2_X1  g0138(.A1(G33), .A2(G87), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n259), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n332), .B1(new_n334), .B2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n340), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n342), .A2(new_n292), .A3(new_n275), .A4(new_n333), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n331), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  AND2_X1   g0144(.A1(new_n343), .A2(new_n331), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n253), .A2(new_n254), .ZN(new_n347));
  XNOR2_X1  g0147(.A(KEYINPUT80), .B(KEYINPUT7), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n347), .A2(new_n348), .A3(new_n214), .ZN(new_n349));
  OR2_X1    g0149(.A1(KEYINPUT3), .A2(G33), .ZN(new_n350));
  NAND2_X1  g0150(.A1(KEYINPUT3), .A2(G33), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n350), .A2(new_n214), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(KEYINPUT7), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n349), .A2(new_n353), .A3(G68), .ZN(new_n354));
  XNOR2_X1  g0154(.A(G58), .B(G68), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n355), .A2(G20), .B1(G159), .B2(new_n306), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n354), .A2(KEYINPUT16), .A3(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT81), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT16), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n352), .A2(new_n348), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n350), .A2(KEYINPUT7), .A3(new_n214), .A4(new_n351), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n226), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n356), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n360), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n354), .A2(KEYINPUT81), .A3(KEYINPUT16), .A4(new_n356), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n359), .A2(new_n310), .A3(new_n365), .A4(new_n366), .ZN(new_n367));
  OR2_X1    g0167(.A1(KEYINPUT8), .A2(G58), .ZN(new_n368));
  NAND2_X1  g0168(.A1(KEYINPUT8), .A2(G58), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n213), .A2(G13), .A3(G20), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n372), .B1(new_n312), .B2(new_n370), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n367), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n346), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(KEYINPUT18), .ZN(new_n376));
  AND2_X1   g0176(.A1(new_n367), .A2(new_n373), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n342), .A2(G190), .A3(new_n275), .A4(new_n333), .ZN(new_n378));
  OAI21_X1  g0178(.A(G200), .B1(new_n334), .B2(new_n340), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n377), .A2(KEYINPUT17), .A3(new_n378), .A4(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT18), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n346), .A2(new_n374), .A3(new_n381), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n367), .A2(new_n373), .A3(new_n378), .A4(new_n379), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT17), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n376), .A2(new_n380), .A3(new_n382), .A4(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n347), .B1(G222), .B2(new_n249), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n387), .B1(new_n335), .B2(new_n249), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n350), .A2(new_n351), .ZN(new_n389));
  OAI211_X1 g0189(.A(new_n388), .B(new_n260), .C1(G77), .C2(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n270), .B1(new_n264), .B2(new_n266), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(G226), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n390), .A2(new_n275), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(new_n332), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n371), .A2(G50), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n312), .A2(G50), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n298), .A2(new_n300), .A3(new_n368), .A4(new_n369), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n306), .A2(G150), .ZN(new_n399));
  AND3_X1   g0199(.A1(new_n398), .A2(KEYINPUT69), .A3(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(KEYINPUT69), .B1(new_n398), .B2(new_n399), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n214), .B1(new_n201), .B2(new_n203), .ZN(new_n402));
  NOR3_X1   g0202(.A1(new_n400), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n310), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n396), .B(new_n397), .C1(new_n403), .C2(new_n404), .ZN(new_n405));
  OAI211_X1 g0205(.A(new_n394), .B(new_n405), .C1(G179), .C2(new_n393), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n371), .A2(G77), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n312), .A2(G77), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n370), .ZN(new_n411));
  INV_X1    g0211(.A(new_n306), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(KEYINPUT70), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT70), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n306), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n411), .A2(new_n413), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(G20), .A2(G77), .ZN(new_n417));
  NOR2_X1   g0217(.A1(KEYINPUT15), .A2(G87), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT71), .ZN(new_n420));
  NAND2_X1  g0220(.A1(KEYINPUT15), .A2(G87), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n419), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n421), .ZN(new_n423));
  OAI21_X1  g0223(.A(KEYINPUT71), .B1(new_n423), .B2(new_n418), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n416), .B(new_n417), .C1(new_n425), .C2(new_n301), .ZN(new_n426));
  AOI211_X1 g0226(.A(new_n408), .B(new_n410), .C1(new_n426), .C2(new_n310), .ZN(new_n427));
  NAND2_X1  g0227(.A1(G238), .A2(G1698), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n389), .B(new_n428), .C1(new_n251), .C2(G1698), .ZN(new_n429));
  INV_X1    g0229(.A(G107), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n347), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n429), .A2(new_n260), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n391), .A2(G244), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n432), .A2(new_n433), .A3(new_n275), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(new_n332), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  OAI21_X1  g0236(.A(KEYINPUT72), .B1(new_n427), .B2(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n408), .B1(new_n426), .B2(new_n310), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n409), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT72), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n439), .A2(new_n440), .A3(new_n435), .ZN(new_n441));
  OR2_X1    g0241(.A1(new_n434), .A2(G179), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n437), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(G190), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n427), .B1(new_n445), .B2(new_n434), .ZN(new_n446));
  AND2_X1   g0246(.A1(new_n434), .A2(G200), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  OR4_X1    g0248(.A1(new_n386), .A2(new_n407), .A3(new_n444), .A4(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n405), .A2(KEYINPUT73), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT9), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n398), .A2(new_n399), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT69), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n402), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n398), .A2(KEYINPUT69), .A3(new_n399), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n395), .B1(new_n457), .B2(new_n310), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT73), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n458), .A2(new_n459), .A3(new_n397), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n450), .A2(new_n451), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n393), .A2(G200), .ZN(new_n462));
  AND2_X1   g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  OR2_X1    g0263(.A1(new_n393), .A2(new_n445), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT74), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n450), .A2(new_n460), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n465), .B1(new_n466), .B2(KEYINPUT9), .ZN(new_n467));
  AOI211_X1 g0267(.A(KEYINPUT74), .B(new_n451), .C1(new_n450), .C2(new_n460), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n463), .B(new_n464), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(KEYINPUT10), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n461), .A2(new_n462), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n405), .A2(KEYINPUT73), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n459), .B1(new_n458), .B2(new_n397), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  OAI21_X1  g0274(.A(KEYINPUT74), .B1(new_n474), .B2(new_n451), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n466), .A2(new_n465), .A3(KEYINPUT9), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n471), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT10), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n477), .A2(new_n478), .A3(new_n464), .ZN(new_n479));
  AOI211_X1 g0279(.A(new_n330), .B(new_n449), .C1(new_n470), .C2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT24), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n214), .B(G87), .C1(new_n253), .C2(new_n254), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(KEYINPUT22), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT22), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n389), .A2(new_n484), .A3(new_n214), .A4(G87), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n214), .A2(G33), .A3(G116), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT23), .ZN(new_n488));
  NOR3_X1   g0288(.A1(new_n488), .A2(new_n214), .A3(G107), .ZN(new_n489));
  AOI21_X1  g0289(.A(KEYINPUT23), .B1(new_n430), .B2(G20), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  AND4_X1   g0292(.A1(new_n481), .A2(new_n486), .A3(new_n487), .A4(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n491), .B1(new_n483), .B2(new_n485), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n481), .B1(new_n494), .B2(new_n487), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n310), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT84), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n497), .B1(new_n297), .B2(G1), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n213), .A2(KEYINPUT84), .A3(G33), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n404), .A2(new_n371), .A3(new_n498), .A4(new_n499), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n500), .A2(new_n430), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n316), .A2(G20), .A3(new_n430), .ZN(new_n503));
  XNOR2_X1  g0303(.A(new_n503), .B(KEYINPUT25), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n496), .A2(new_n502), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n221), .A2(new_n249), .ZN(new_n507));
  INV_X1    g0307(.A(G257), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(G1698), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n507), .B(new_n509), .C1(new_n253), .C2(new_n254), .ZN(new_n510));
  NAND2_X1  g0310(.A1(G33), .A2(G294), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n260), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n269), .A2(G1), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT5), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(G41), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n268), .A2(KEYINPUT5), .ZN(new_n517));
  AND3_X1   g0317(.A1(new_n514), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n267), .A2(G274), .A3(new_n518), .ZN(new_n519));
  XNOR2_X1  g0319(.A(KEYINPUT5), .B(G41), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n514), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n267), .A2(G264), .A3(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n513), .A2(new_n519), .A3(new_n522), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n523), .A2(new_n292), .ZN(new_n524));
  AOI22_X1  g0324(.A1(new_n264), .A2(new_n266), .B1(new_n520), .B2(new_n514), .ZN(new_n525));
  AOI22_X1  g0325(.A1(new_n525), .A2(G264), .B1(new_n512), .B2(new_n260), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n332), .B1(new_n526), .B2(new_n519), .ZN(new_n527));
  OAI21_X1  g0327(.A(KEYINPUT94), .B1(new_n524), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n523), .A2(G169), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT94), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n529), .B(new_n530), .C1(new_n292), .C2(new_n523), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n506), .A2(new_n528), .A3(new_n531), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n513), .A2(new_n519), .A3(new_n522), .A4(new_n445), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(KEYINPUT95), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT95), .ZN(new_n536));
  INV_X1    g0336(.A(G200), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n536), .B1(new_n523), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n535), .B1(new_n534), .B2(new_n538), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n539), .A2(new_n502), .A3(new_n496), .A4(new_n505), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n532), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n267), .A2(G270), .A3(new_n521), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(KEYINPUT91), .ZN(new_n543));
  NAND2_X1  g0343(.A1(G264), .A2(G1698), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n389), .B(new_n544), .C1(new_n508), .C2(G1698), .ZN(new_n545));
  INV_X1    g0345(.A(G303), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n347), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n545), .A2(new_n260), .A3(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT91), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n267), .A2(new_n549), .A3(new_n521), .A4(G270), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n543), .A2(new_n519), .A3(new_n548), .A4(new_n550), .ZN(new_n551));
  AND2_X1   g0351(.A1(new_n551), .A2(G200), .ZN(new_n552));
  INV_X1    g0352(.A(G116), .ZN(new_n553));
  AOI22_X1  g0353(.A1(new_n309), .A2(new_n263), .B1(G20), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(G33), .A2(G283), .ZN(new_n555));
  INV_X1    g0355(.A(G97), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n555), .B(new_n214), .C1(G33), .C2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n554), .A2(KEYINPUT20), .A3(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(KEYINPUT20), .B1(new_n554), .B2(new_n557), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n371), .A2(new_n553), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n563), .B1(new_n500), .B2(G116), .ZN(new_n564));
  OAI21_X1  g0364(.A(KEYINPUT92), .B1(new_n561), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n553), .A2(G20), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n557), .A2(new_n310), .A3(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT20), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n558), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n498), .A2(new_n263), .A3(new_n309), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n371), .A2(new_n499), .ZN(new_n572));
  OAI21_X1  g0372(.A(G116), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n562), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT92), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n570), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n565), .A2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT93), .ZN(new_n578));
  NOR3_X1   g0378(.A1(new_n552), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  AND3_X1   g0379(.A1(new_n570), .A2(new_n574), .A3(new_n575), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n575), .B1(new_n570), .B2(new_n574), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n551), .A2(G200), .ZN(new_n583));
  AOI21_X1  g0383(.A(KEYINPUT93), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n551), .A2(new_n445), .ZN(new_n585));
  NOR3_X1   g0385(.A1(new_n579), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT21), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n551), .A2(G169), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n587), .B1(new_n582), .B2(new_n588), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n577), .A2(KEYINPUT21), .A3(G169), .A4(new_n551), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n551), .A2(new_n292), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n577), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n589), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  NOR3_X1   g0393(.A1(new_n541), .A2(new_n586), .A3(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT4), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n595), .A2(G1698), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n596), .B(G244), .C1(new_n254), .C2(new_n253), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n219), .B1(new_n350), .B2(new_n351), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n597), .B(new_n555), .C1(new_n598), .C2(KEYINPUT4), .ZN(new_n599));
  OAI21_X1  g0399(.A(G250), .B1(new_n253), .B2(new_n254), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n249), .B1(new_n600), .B2(KEYINPUT4), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n260), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(G274), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n603), .B1(new_n264), .B2(new_n266), .ZN(new_n604));
  AOI22_X1  g0404(.A1(G257), .A2(new_n525), .B1(new_n604), .B2(new_n518), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n602), .A2(new_n605), .A3(G190), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT86), .ZN(new_n607));
  XNOR2_X1  g0407(.A(new_n606), .B(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(new_n500), .ZN(new_n609));
  OR3_X1    g0409(.A1(new_n371), .A2(KEYINPUT83), .A3(G97), .ZN(new_n610));
  OAI21_X1  g0410(.A(KEYINPUT83), .B1(new_n371), .B2(G97), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n609), .A2(G97), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n430), .B1(new_n361), .B2(new_n362), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT6), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n556), .A2(new_n430), .ZN(new_n615));
  NOR2_X1   g0415(.A1(G97), .A2(G107), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n614), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n430), .A2(KEYINPUT6), .A3(G97), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n214), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n412), .A2(new_n202), .ZN(new_n620));
  NOR3_X1   g0420(.A1(new_n613), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n612), .B1(new_n621), .B2(new_n404), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n267), .A2(G257), .A3(new_n521), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n519), .A2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT85), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n519), .A2(new_n623), .A3(KEYINPUT85), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n626), .A2(new_n602), .A3(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n622), .B1(G200), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n608), .A2(new_n629), .ZN(new_n630));
  NOR3_X1   g0430(.A1(new_n253), .A2(new_n254), .A3(G20), .ZN(new_n631));
  XOR2_X1   g0431(.A(KEYINPUT80), .B(KEYINPUT7), .Z(new_n632));
  OAI21_X1  g0432(.A(new_n362), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(G107), .ZN(new_n634));
  INV_X1    g0434(.A(new_n620), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n617), .A2(new_n618), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(G20), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n634), .A2(new_n635), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n310), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n602), .A2(new_n605), .ZN(new_n640));
  AOI22_X1  g0440(.A1(new_n639), .A2(new_n612), .B1(new_n640), .B2(new_n332), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n626), .A2(new_n292), .A3(new_n602), .A4(new_n627), .ZN(new_n642));
  AOI21_X1  g0442(.A(KEYINPUT87), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n640), .A2(new_n332), .ZN(new_n644));
  AND4_X1   g0444(.A1(KEYINPUT87), .A2(new_n642), .A3(new_n644), .A4(new_n622), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n630), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT88), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n371), .B1(new_n422), .B2(new_n424), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n298), .A2(new_n300), .A3(G97), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT19), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n389), .A2(new_n214), .A3(G68), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n214), .B1(new_n256), .B2(new_n651), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n220), .A2(new_n556), .A3(new_n430), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n652), .A2(new_n653), .A3(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n649), .B1(new_n657), .B2(new_n310), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT90), .ZN(new_n659));
  INV_X1    g0459(.A(new_n425), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n609), .A2(new_n660), .ZN(new_n661));
  AND3_X1   g0461(.A1(new_n658), .A2(new_n659), .A3(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n659), .B1(new_n658), .B2(new_n661), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  AOI21_X1  g0464(.A(G250), .B1(new_n213), .B2(G45), .ZN(new_n665));
  NOR3_X1   g0465(.A1(new_n269), .A2(G1), .A3(G274), .ZN(new_n666));
  AOI211_X1 g0466(.A(new_n665), .B(new_n666), .C1(new_n264), .C2(new_n266), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n227), .A2(new_n249), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n219), .A2(G1698), .ZN(new_n669));
  OAI211_X1 g0469(.A(new_n668), .B(new_n669), .C1(new_n253), .C2(new_n254), .ZN(new_n670));
  NAND2_X1  g0470(.A1(G33), .A2(G116), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n259), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(KEYINPUT89), .B1(new_n667), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n670), .A2(new_n671), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(new_n260), .ZN(new_n675));
  INV_X1    g0475(.A(new_n665), .ZN(new_n676));
  INV_X1    g0476(.A(new_n666), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n267), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT89), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n675), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  AND3_X1   g0480(.A1(new_n673), .A2(new_n332), .A3(new_n680), .ZN(new_n681));
  AOI21_X1  g0481(.A(G179), .B1(new_n673), .B2(new_n680), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NOR3_X1   g0483(.A1(new_n667), .A2(new_n672), .A3(KEYINPUT89), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n679), .B1(new_n675), .B2(new_n678), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(G200), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n445), .B1(new_n673), .B2(new_n680), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n609), .A2(G87), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n658), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  AOI22_X1  g0491(.A1(new_n664), .A2(new_n683), .B1(new_n687), .B2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n642), .A2(new_n622), .A3(new_n644), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT87), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n641), .A2(KEYINPUT87), .A3(new_n642), .ZN(new_n697));
  AOI22_X1  g0497(.A1(new_n696), .A2(new_n697), .B1(new_n629), .B2(new_n608), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n693), .B1(new_n698), .B2(KEYINPUT88), .ZN(new_n699));
  AND4_X1   g0499(.A1(new_n480), .A2(new_n594), .A3(new_n648), .A4(new_n699), .ZN(G372));
  AOI21_X1  g0500(.A(new_n665), .B1(new_n264), .B2(new_n266), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT96), .ZN(new_n702));
  AND3_X1   g0502(.A1(new_n701), .A2(new_n702), .A3(new_n677), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n702), .B1(new_n701), .B2(new_n677), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n675), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(G200), .ZN(new_n706));
  AND2_X1   g0506(.A1(new_n658), .A2(new_n689), .ZN(new_n707));
  OAI21_X1  g0507(.A(G190), .B1(new_n684), .B2(new_n685), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n706), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n705), .A2(new_n332), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n292), .B1(new_n684), .B2(new_n685), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n658), .A2(new_n661), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n710), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n709), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n486), .A2(new_n487), .A3(new_n492), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(KEYINPUT24), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n494), .A2(new_n481), .A3(new_n487), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n404), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NOR3_X1   g0518(.A1(new_n718), .A2(new_n501), .A3(new_n504), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n714), .B1(new_n719), .B2(new_n539), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n529), .B1(new_n292), .B2(new_n523), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n506), .A2(new_n721), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n722), .A2(new_n589), .A3(new_n590), .A4(new_n592), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n720), .A2(new_n723), .A3(new_n698), .ZN(new_n724));
  INV_X1    g0524(.A(new_n713), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n691), .A2(new_n687), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n712), .A2(KEYINPUT90), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n673), .A2(new_n680), .A3(new_n332), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n658), .A2(new_n659), .A3(new_n661), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n727), .A2(new_n711), .A3(new_n728), .A4(new_n729), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n696), .A2(new_n697), .A3(new_n726), .A4(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n725), .B1(new_n731), .B2(KEYINPUT26), .ZN(new_n732));
  AND2_X1   g0532(.A1(new_n709), .A2(new_n713), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT26), .ZN(new_n734));
  INV_X1    g0534(.A(new_n694), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n733), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n724), .A2(new_n732), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n480), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT97), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n478), .B1(new_n477), .B2(new_n464), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n469), .A2(KEYINPUT10), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n479), .A2(new_n470), .A3(KEYINPUT97), .ZN(new_n743));
  AND2_X1   g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g0544(.A(new_n293), .B(KEYINPUT79), .ZN(new_n745));
  AND2_X1   g0545(.A1(new_n289), .A2(new_n291), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n320), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n747), .B1(new_n329), .B2(new_n444), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n380), .A2(new_n385), .ZN(new_n749));
  OAI211_X1 g0549(.A(new_n376), .B(new_n382), .C1(new_n748), .C2(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n407), .B1(new_n744), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n738), .A2(new_n751), .ZN(G369));
  NOR2_X1   g0552(.A1(new_n586), .A2(new_n593), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n315), .A2(G20), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n316), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(KEYINPUT27), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT98), .ZN(new_n757));
  XNOR2_X1  g0557(.A(new_n756), .B(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n755), .A2(KEYINPUT27), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n758), .A2(G213), .A3(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(G343), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(new_n582), .ZN(new_n764));
  MUX2_X1   g0564(.A(new_n753), .B(new_n593), .S(new_n764), .Z(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(G330), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n719), .A2(new_n763), .ZN(new_n768));
  OAI22_X1  g0568(.A1(new_n541), .A2(new_n768), .B1(new_n532), .B2(new_n763), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n593), .A2(new_n763), .ZN(new_n771));
  OAI22_X1  g0571(.A1(new_n771), .A2(new_n541), .B1(new_n722), .B2(new_n762), .ZN(new_n772));
  INV_X1    g0572(.A(KEYINPUT99), .ZN(new_n773));
  XNOR2_X1  g0573(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n770), .A2(new_n774), .ZN(G399));
  INV_X1    g0575(.A(new_n215), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(G41), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n655), .A2(G116), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n778), .A2(G1), .A3(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n209), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n780), .B1(new_n781), .B2(new_n778), .ZN(new_n782));
  XNOR2_X1  g0582(.A(new_n782), .B(KEYINPUT28), .ZN(new_n783));
  INV_X1    g0583(.A(KEYINPUT29), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n733), .A2(new_n540), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n646), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(KEYINPUT103), .ZN(new_n787));
  INV_X1    g0587(.A(new_n593), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n787), .B1(new_n788), .B2(new_n532), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n528), .A2(new_n531), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n719), .A2(new_n790), .ZN(new_n791));
  NOR3_X1   g0591(.A1(new_n791), .A2(new_n593), .A3(KEYINPUT103), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n786), .B1(new_n789), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(KEYINPUT104), .ZN(new_n794));
  NAND4_X1  g0594(.A1(new_n692), .A2(new_n734), .A3(new_n696), .A4(new_n697), .ZN(new_n795));
  NAND4_X1  g0595(.A1(new_n709), .A2(new_n713), .A3(new_n642), .A4(new_n641), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n725), .B1(new_n796), .B2(KEYINPUT26), .ZN(new_n797));
  AND3_X1   g0597(.A1(new_n795), .A2(new_n797), .A3(KEYINPUT102), .ZN(new_n798));
  AOI21_X1  g0598(.A(KEYINPUT102), .B1(new_n795), .B2(new_n797), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(KEYINPUT104), .ZN(new_n801));
  OAI211_X1 g0601(.A(new_n786), .B(new_n801), .C1(new_n789), .C2(new_n792), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n794), .A2(new_n800), .A3(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n784), .B1(new_n803), .B2(new_n763), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n737), .A2(new_n763), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n805), .A2(KEYINPUT29), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  OR2_X1    g0607(.A1(new_n686), .A2(new_n640), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n591), .A2(new_n526), .ZN(new_n809));
  INV_X1    g0609(.A(KEYINPUT30), .ZN(new_n810));
  OR3_X1    g0610(.A1(new_n808), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n810), .B1(new_n808), .B2(new_n809), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n628), .A2(new_n523), .ZN(new_n814));
  INV_X1    g0614(.A(KEYINPUT100), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n816), .A2(new_n551), .A3(new_n705), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n292), .B1(new_n814), .B2(new_n815), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  OAI211_X1 g0619(.A(KEYINPUT31), .B(new_n762), .C1(new_n813), .C2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT101), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n820), .B(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n762), .B1(new_n813), .B2(new_n819), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  NAND4_X1  g0624(.A1(new_n594), .A2(new_n648), .A3(new_n699), .A4(new_n763), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n824), .B1(new_n825), .B2(KEYINPUT31), .ZN(new_n826));
  OAI21_X1  g0626(.A(G330), .B1(new_n822), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n807), .A2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n783), .B1(new_n829), .B2(G1), .ZN(G364));
  NAND2_X1  g0630(.A1(new_n754), .A2(G45), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n778), .A2(G1), .A3(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n765), .A2(G330), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n832), .B1(new_n767), .B2(new_n833), .ZN(new_n834));
  AND2_X1   g0634(.A1(KEYINPUT107), .A2(G169), .ZN(new_n835));
  NOR2_X1   g0635(.A1(KEYINPUT107), .A2(G169), .ZN(new_n836));
  NOR3_X1   g0636(.A1(new_n835), .A2(new_n836), .A3(new_n214), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n837), .A2(new_n263), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n214), .A2(new_n445), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n292), .A2(G200), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n389), .B1(new_n842), .B2(G322), .ZN(new_n843));
  INV_X1    g0643(.A(G294), .ZN(new_n844));
  NOR2_X1   g0644(.A1(G179), .A2(G200), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(G190), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(G20), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n292), .A2(new_n537), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n214), .A2(G190), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  XOR2_X1   g0651(.A(KEYINPUT33), .B(G317), .Z(new_n852));
  OAI221_X1 g0652(.A(new_n843), .B1(new_n844), .B2(new_n848), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n537), .A2(G179), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n850), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n850), .A2(new_n845), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  AOI22_X1  g0658(.A1(G283), .A2(new_n856), .B1(new_n858), .B2(G329), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n839), .A2(new_n854), .ZN(new_n860));
  INV_X1    g0660(.A(G311), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n850), .A2(new_n840), .ZN(new_n862));
  OAI221_X1 g0662(.A(new_n859), .B1(new_n546), .B2(new_n860), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n839), .A2(new_n849), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  AOI211_X1 g0665(.A(new_n853), .B(new_n863), .C1(G326), .C2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n860), .ZN(new_n867));
  AOI22_X1  g0667(.A1(G50), .A2(new_n865), .B1(new_n867), .B2(G87), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n868), .B1(new_n430), .B2(new_n855), .ZN(new_n869));
  INV_X1    g0669(.A(G159), .ZN(new_n870));
  OR3_X1    g0670(.A1(new_n857), .A2(KEYINPUT32), .A3(new_n870), .ZN(new_n871));
  OAI21_X1  g0671(.A(KEYINPUT32), .B1(new_n857), .B2(new_n870), .ZN(new_n872));
  OAI211_X1 g0672(.A(new_n871), .B(new_n872), .C1(new_n556), .C2(new_n848), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n862), .A2(new_n202), .ZN(new_n874));
  INV_X1    g0674(.A(G58), .ZN(new_n875));
  OAI221_X1 g0675(.A(new_n389), .B1(new_n841), .B2(new_n875), .C1(new_n226), .C2(new_n851), .ZN(new_n876));
  NOR4_X1   g0676(.A1(new_n869), .A2(new_n873), .A3(new_n874), .A4(new_n876), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n838), .B1(new_n866), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n209), .A2(new_n269), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n347), .A2(new_n215), .ZN(new_n880));
  XNOR2_X1  g0680(.A(new_n880), .B(KEYINPUT105), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n879), .B(new_n881), .C1(new_n269), .C2(new_n244), .ZN(new_n882));
  INV_X1    g0682(.A(G355), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n389), .A2(new_n215), .ZN(new_n884));
  OAI221_X1 g0684(.A(new_n882), .B1(G116), .B2(new_n215), .C1(new_n883), .C2(new_n884), .ZN(new_n885));
  NOR2_X1   g0685(.A1(G13), .A2(G33), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n214), .ZN(new_n887));
  XOR2_X1   g0687(.A(new_n887), .B(KEYINPUT106), .Z(new_n888));
  INV_X1    g0688(.A(new_n838), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n885), .A2(new_n891), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n878), .B(new_n892), .C1(new_n765), .C2(new_n888), .ZN(new_n893));
  INV_X1    g0693(.A(new_n832), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n834), .A2(new_n895), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n896), .B(KEYINPUT108), .ZN(G396));
  INV_X1    g0697(.A(KEYINPUT109), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n763), .A2(new_n427), .ZN(new_n899));
  AND3_X1   g0699(.A1(new_n443), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  AND2_X1   g0700(.A1(new_n443), .A2(new_n448), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n899), .B1(new_n443), .B2(new_n898), .ZN(new_n902));
  NOR3_X1   g0702(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n805), .B(new_n903), .ZN(new_n904));
  XNOR2_X1  g0704(.A(new_n827), .B(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(new_n832), .ZN(new_n906));
  INV_X1    g0706(.A(new_n851), .ZN(new_n907));
  AOI22_X1  g0707(.A1(G143), .A2(new_n842), .B1(new_n907), .B2(G150), .ZN(new_n908));
  INV_X1    g0708(.A(G137), .ZN(new_n909));
  OAI221_X1 g0709(.A(new_n908), .B1(new_n909), .B2(new_n864), .C1(new_n870), .C2(new_n862), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n910), .B(KEYINPUT34), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n855), .A2(new_n226), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n389), .B1(new_n860), .B2(new_n224), .ZN(new_n913));
  AOI211_X1 g0713(.A(new_n912), .B(new_n913), .C1(G58), .C2(new_n847), .ZN(new_n914));
  INV_X1    g0714(.A(G132), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n911), .B(new_n914), .C1(new_n915), .C2(new_n857), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n855), .A2(new_n220), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n917), .B1(G294), .B2(new_n842), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(new_n430), .B2(new_n860), .ZN(new_n919));
  INV_X1    g0719(.A(new_n862), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n919), .B1(G116), .B2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(G283), .ZN(new_n922));
  OAI221_X1 g0722(.A(new_n347), .B1(new_n851), .B2(new_n922), .C1(new_n546), .C2(new_n864), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n923), .B1(G97), .B2(new_n847), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n921), .B(new_n924), .C1(new_n861), .C2(new_n857), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n889), .B1(new_n916), .B2(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n838), .A2(new_n886), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n926), .B1(new_n202), .B2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(new_n886), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n928), .B(new_n894), .C1(new_n903), .C2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n906), .A2(new_n930), .ZN(G384));
  INV_X1    g0731(.A(KEYINPUT38), .ZN(new_n932));
  INV_X1    g0732(.A(new_n760), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n359), .A2(new_n310), .A3(new_n366), .ZN(new_n934));
  AOI21_X1  g0734(.A(KEYINPUT16), .B1(new_n354), .B2(new_n356), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n373), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  AND3_X1   g0736(.A1(new_n386), .A2(new_n933), .A3(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n760), .B1(new_n344), .B2(new_n345), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n374), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT37), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n939), .A2(new_n940), .A3(new_n383), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT112), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND4_X1  g0743(.A1(new_n939), .A2(KEYINPUT112), .A3(new_n940), .A4(new_n383), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n938), .A2(new_n936), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n383), .ZN(new_n946));
  AOI22_X1  g0746(.A1(new_n943), .A2(new_n944), .B1(KEYINPUT37), .B2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n932), .B1(new_n937), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n943), .A2(new_n944), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n946), .A2(KEYINPUT37), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n386), .A2(new_n933), .A3(new_n936), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n951), .A2(KEYINPUT38), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n948), .A2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(new_n903), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n320), .A2(new_n763), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n330), .A2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(new_n956), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n322), .A2(new_n329), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n955), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT113), .ZN(new_n961));
  OR2_X1    g0761(.A1(new_n961), .A2(KEYINPUT40), .ZN(new_n962));
  INV_X1    g0762(.A(new_n820), .ZN(new_n963));
  OAI211_X1 g0763(.A(new_n960), .B(new_n962), .C1(new_n826), .C2(new_n963), .ZN(new_n964));
  AND3_X1   g0764(.A1(new_n322), .A2(new_n329), .A3(new_n958), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n958), .B1(new_n322), .B2(new_n329), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n903), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n825), .A2(KEYINPUT31), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(new_n823), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n967), .B1(new_n969), .B2(new_n820), .ZN(new_n970));
  OAI211_X1 g0770(.A(new_n954), .B(new_n964), .C1(new_n970), .C2(new_n961), .ZN(new_n971));
  AND3_X1   g0771(.A1(new_n386), .A2(new_n374), .A3(new_n933), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n939), .A2(new_n383), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n943), .A2(new_n944), .B1(KEYINPUT37), .B2(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n932), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n953), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n960), .B1(new_n826), .B2(new_n963), .ZN(new_n979));
  OAI21_X1  g0779(.A(KEYINPUT40), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n971), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n480), .B1(new_n826), .B2(new_n963), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n981), .B(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(G330), .ZN(new_n984));
  AND3_X1   g0784(.A1(new_n948), .A2(new_n953), .A3(KEYINPUT39), .ZN(new_n985));
  AOI21_X1  g0785(.A(KEYINPUT39), .B1(new_n975), .B2(new_n953), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n322), .A2(new_n762), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n376), .A2(new_n382), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(new_n760), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n737), .A2(new_n903), .A3(new_n763), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n443), .A2(new_n762), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n992), .A2(new_n994), .B1(new_n957), .B2(new_n959), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(new_n954), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n989), .A2(new_n991), .A3(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n480), .B1(new_n804), .B2(new_n806), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n998), .A2(new_n751), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n997), .B(new_n999), .Z(new_n1000));
  XNOR2_X1  g0800(.A(new_n984), .B(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n213), .B2(new_n754), .ZN(new_n1002));
  OAI211_X1 g0802(.A(G20), .B(new_n210), .C1(new_n636), .C2(KEYINPUT35), .ZN(new_n1003));
  AOI211_X1 g0803(.A(new_n553), .B(new_n1003), .C1(KEYINPUT35), .C2(new_n636), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n1004), .B(KEYINPUT36), .Z(new_n1005));
  OAI211_X1 g0805(.A(new_n209), .B(G77), .C1(new_n875), .C2(new_n226), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT110), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n201), .A2(G68), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n1006), .A2(new_n1007), .B1(KEYINPUT111), .B2(new_n1008), .ZN(new_n1009));
  OR2_X1    g0809(.A1(new_n1008), .A2(KEYINPUT111), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n1009), .B(new_n1010), .C1(new_n1007), .C2(new_n1006), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1011), .A2(G1), .A3(new_n315), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1002), .A2(new_n1005), .A3(new_n1012), .ZN(G367));
  NAND2_X1  g0813(.A1(new_n831), .A2(G1), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n762), .A2(new_n622), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n698), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n735), .A2(new_n762), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n774), .A2(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT44), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n774), .A2(new_n1018), .ZN(new_n1021));
  XOR2_X1   g0821(.A(KEYINPUT115), .B(KEYINPUT45), .Z(new_n1022));
  XNOR2_X1  g0822(.A(new_n1021), .B(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1020), .A2(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(new_n770), .ZN(new_n1025));
  OR2_X1    g0825(.A1(new_n766), .A2(KEYINPUT116), .ZN(new_n1026));
  OR2_X1    g0826(.A1(new_n771), .A2(new_n541), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n771), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1027), .B1(new_n769), .B2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1029), .B1(new_n766), .B2(KEYINPUT116), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n1026), .B(new_n1030), .Z(new_n1031));
  INV_X1    g0831(.A(new_n1031), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1025), .A2(new_n829), .A3(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(new_n829), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n777), .B(KEYINPUT41), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1014), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n1027), .A2(new_n1016), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT42), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n1018), .A2(new_n791), .B1(new_n696), .B2(new_n697), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1038), .B1(new_n762), .B2(new_n1039), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n763), .A2(new_n707), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(new_n725), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n714), .B2(new_n1041), .ZN(new_n1043));
  OR2_X1    g0843(.A1(new_n1043), .A2(KEYINPUT43), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(KEYINPUT43), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1040), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT114), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n1044), .B2(new_n1040), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n767), .A2(new_n769), .A3(new_n1018), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1048), .B(new_n1049), .ZN(new_n1050));
  OR2_X1    g0850(.A1(new_n1036), .A2(new_n1050), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n841), .A2(new_n546), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n347), .B1(new_n851), .B2(new_n844), .ZN(new_n1053));
  AOI211_X1 g0853(.A(new_n1052), .B(new_n1053), .C1(G107), .C2(new_n847), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1054), .B1(new_n556), .B2(new_n855), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n867), .A2(G116), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT46), .ZN(new_n1057));
  INV_X1    g0857(.A(G317), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n1057), .B1(new_n861), .B2(new_n864), .C1(new_n1058), .C2(new_n857), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n1055), .B(new_n1059), .C1(G283), .C2(new_n920), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n347), .B1(new_n842), .B2(G150), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n1061), .B1(new_n875), .B2(new_n860), .C1(new_n226), .C2(new_n848), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(G77), .A2(new_n856), .B1(new_n858), .B2(G137), .ZN(new_n1063));
  INV_X1    g0863(.A(G143), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n1063), .B1(new_n1064), .B2(new_n864), .C1(new_n201), .C2(new_n862), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n1062), .B(new_n1065), .C1(G159), .C2(new_n907), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1060), .A2(new_n1066), .ZN(new_n1067));
  XOR2_X1   g0867(.A(new_n1067), .B(KEYINPUT47), .Z(new_n1068));
  AOI21_X1  g0868(.A(new_n832), .B1(new_n1068), .B2(new_n838), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n881), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n891), .B1(new_n215), .B2(new_n425), .C1(new_n240), .C2(new_n1070), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1069), .B(new_n1071), .C1(new_n888), .C2(new_n1043), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1051), .A2(new_n1072), .ZN(G387));
  NAND2_X1  g0873(.A1(new_n1032), .A2(new_n829), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n778), .B1(new_n1031), .B2(new_n828), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n881), .B1(new_n236), .B2(new_n269), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1077), .B1(new_n779), .B2(new_n884), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n226), .A2(new_n202), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n411), .A2(new_n224), .ZN(new_n1080));
  AOI211_X1 g0880(.A(G116), .B(new_n655), .C1(new_n1080), .C2(KEYINPUT50), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1081), .B(new_n269), .C1(KEYINPUT50), .C2(new_n1080), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1078), .B1(new_n1079), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n776), .A2(new_n430), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n890), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  AND2_X1   g0885(.A1(new_n858), .A2(G326), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(G311), .A2(new_n907), .B1(new_n842), .B2(G317), .ZN(new_n1087));
  INV_X1    g0887(.A(G322), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n1087), .B1(new_n546), .B2(new_n862), .C1(new_n1088), .C2(new_n864), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT48), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n1090), .B1(new_n922), .B2(new_n848), .C1(new_n844), .C2(new_n860), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT49), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n389), .B(new_n1086), .C1(new_n1091), .C2(new_n1092), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n1093), .B1(new_n1092), .B2(new_n1091), .C1(new_n553), .C2(new_n855), .ZN(new_n1094));
  INV_X1    g0894(.A(G150), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n857), .A2(new_n1095), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n864), .A2(new_n870), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n841), .A2(new_n224), .B1(new_n862), .B2(new_n226), .ZN(new_n1098));
  AOI211_X1 g0898(.A(new_n1097), .B(new_n1098), .C1(new_n411), .C2(new_n907), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n660), .A2(new_n847), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n389), .B1(new_n855), .B2(new_n556), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(G77), .B2(new_n867), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1099), .A2(new_n1100), .A3(new_n1102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1094), .B1(new_n1096), .B2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1085), .B1(new_n1104), .B2(new_n838), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n1105), .B(new_n894), .C1(new_n769), .C2(new_n888), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1014), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n1076), .B(new_n1106), .C1(new_n1107), .C2(new_n1031), .ZN(G393));
  INV_X1    g0908(.A(new_n1025), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n778), .B1(new_n1109), .B2(new_n1074), .ZN(new_n1110));
  AND2_X1   g0910(.A1(new_n1110), .A2(new_n1033), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n920), .A2(G294), .B1(new_n847), .B2(G116), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1112), .B1(new_n546), .B2(new_n851), .ZN(new_n1113));
  OR2_X1    g0913(.A1(new_n1113), .A2(KEYINPUT118), .ZN(new_n1114));
  OAI221_X1 g0914(.A(new_n347), .B1(new_n857), .B2(new_n1088), .C1(new_n430), .C2(new_n855), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1115), .B1(new_n1113), .B2(KEYINPUT118), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n867), .A2(G283), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n864), .A2(new_n1058), .B1(new_n841), .B2(new_n861), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(new_n1118), .B(KEYINPUT52), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n1114), .A2(new_n1116), .A3(new_n1117), .A4(new_n1119), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n864), .A2(new_n1095), .B1(new_n841), .B2(new_n870), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(new_n1121), .B(KEYINPUT117), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n1122), .B(KEYINPUT51), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n848), .A2(new_n202), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n201), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(G68), .A2(new_n867), .B1(new_n907), .B2(new_n1125), .ZN(new_n1126));
  OAI221_X1 g0926(.A(new_n1126), .B1(new_n1064), .B2(new_n857), .C1(new_n370), .C2(new_n862), .ZN(new_n1127));
  OR4_X1    g0927(.A1(new_n347), .A2(new_n1123), .A3(new_n1124), .A4(new_n1127), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1120), .B1(new_n1128), .B2(new_n917), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n832), .B1(new_n1129), .B2(new_n838), .ZN(new_n1130));
  OAI221_X1 g0930(.A(new_n891), .B1(new_n556), .B2(new_n215), .C1(new_n1070), .C2(new_n247), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n1130), .B(new_n1131), .C1(new_n888), .C2(new_n1018), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1132), .B1(new_n1109), .B2(new_n1107), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1111), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(G390));
  NAND3_X1  g0935(.A1(new_n803), .A2(new_n763), .A3(new_n903), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n994), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n965), .A2(new_n966), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n976), .A2(new_n977), .B1(new_n322), .B2(new_n762), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n985), .A2(new_n986), .B1(new_n988), .B2(new_n995), .ZN(new_n1144));
  OAI211_X1 g0944(.A(G330), .B(new_n960), .C1(new_n822), .C2(new_n826), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1143), .A2(KEYINPUT119), .A3(new_n1144), .A4(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1138), .B1(new_n1136), .B2(new_n994), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1144), .B(new_n1145), .C1(new_n1147), .C2(new_n1141), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT119), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1144), .B1(new_n1147), .B2(new_n1141), .ZN(new_n1151));
  OAI211_X1 g0951(.A(G330), .B(new_n903), .C1(new_n826), .C2(new_n963), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1151), .A2(new_n1139), .A3(new_n1153), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1146), .A2(new_n1150), .A3(new_n1154), .A4(new_n1014), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n841), .A2(new_n915), .ZN(new_n1156));
  INV_X1    g0956(.A(G128), .ZN(new_n1157));
  OAI221_X1 g0957(.A(new_n389), .B1(new_n851), .B2(new_n909), .C1(new_n1157), .C2(new_n864), .ZN(new_n1158));
  AOI211_X1 g0958(.A(new_n1156), .B(new_n1158), .C1(G159), .C2(new_n847), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n858), .A2(G125), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n860), .A2(new_n1095), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1161), .B(KEYINPUT53), .ZN(new_n1162));
  XOR2_X1   g0962(.A(KEYINPUT54), .B(G143), .Z(new_n1163));
  AOI22_X1  g0963(.A1(new_n1125), .A2(new_n856), .B1(new_n920), .B2(new_n1163), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n1159), .A2(new_n1160), .A3(new_n1162), .A4(new_n1164), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n864), .A2(new_n922), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n851), .A2(new_n430), .B1(new_n857), .B2(new_n844), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n1166), .B(new_n1167), .C1(G97), .C2(new_n920), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n347), .B1(new_n860), .B2(new_n220), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n912), .B(new_n1169), .C1(G116), .C2(new_n842), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1168), .B(new_n1170), .C1(new_n202), .C2(new_n848), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n889), .B1(new_n1165), .B2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(new_n370), .B2(new_n927), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n894), .B(new_n1173), .C1(new_n987), .C2(new_n929), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1155), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  AND2_X1   g0976(.A1(new_n1136), .A2(new_n994), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1152), .A2(new_n1138), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1177), .A2(new_n1145), .A3(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1179), .A2(KEYINPUT120), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT120), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n1177), .A2(new_n1178), .A3(new_n1181), .A4(new_n1145), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1138), .B1(new_n827), .B2(new_n955), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1184), .B1(new_n1138), .B2(new_n1152), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n992), .A2(new_n994), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1183), .A2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(G330), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n751), .B(new_n998), .C1(new_n982), .C2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1188), .A2(new_n1191), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1146), .A2(new_n1154), .A3(new_n1150), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n777), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1193), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1190), .B1(new_n1183), .B2(new_n1187), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1176), .B1(new_n1194), .B2(new_n1197), .ZN(G378));
  AOI22_X1  g0998(.A1(new_n1180), .A2(new_n1182), .B1(new_n1186), .B2(new_n1185), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1191), .B1(new_n1193), .B2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n981), .A2(G330), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n742), .A2(new_n406), .A3(new_n743), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1202), .A2(KEYINPUT55), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT55), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n742), .A2(new_n1204), .A3(new_n406), .A4(new_n743), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n474), .A2(new_n933), .ZN(new_n1206));
  XOR2_X1   g1006(.A(new_n1206), .B(KEYINPUT56), .Z(new_n1207));
  AND3_X1   g1007(.A1(new_n1203), .A2(new_n1205), .A3(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1207), .B1(new_n1203), .B2(new_n1205), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT121), .ZN(new_n1210));
  NOR3_X1   g1010(.A1(new_n1208), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1201), .A2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n997), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1203), .A2(new_n1205), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1207), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1203), .A2(new_n1205), .A3(new_n1207), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1216), .A2(KEYINPUT121), .A3(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1189), .B1(new_n971), .B2(new_n980), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  AND3_X1   g1020(.A1(new_n1212), .A2(new_n1213), .A3(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1213), .B1(new_n1212), .B2(new_n1220), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1200), .B(KEYINPUT57), .C1(new_n1221), .C2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(new_n777), .ZN(new_n1224));
  AND2_X1   g1024(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n997), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1212), .A2(new_n1213), .A3(new_n1220), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(KEYINPUT57), .B1(new_n1229), .B2(new_n1200), .ZN(new_n1230));
  OR2_X1    g1030(.A1(new_n1224), .A2(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1216), .A2(new_n886), .A3(new_n1217), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n848), .A2(new_n1095), .B1(new_n841), .B2(new_n1157), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n867), .A2(new_n1163), .B1(new_n920), .B2(G137), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1234), .B1(new_n915), .B2(new_n851), .ZN(new_n1235));
  AOI211_X1 g1035(.A(new_n1233), .B(new_n1235), .C1(G125), .C2(new_n865), .ZN(new_n1236));
  XNOR2_X1  g1036(.A(new_n1236), .B(KEYINPUT59), .ZN(new_n1237));
  AOI21_X1  g1037(.A(G41), .B1(new_n858), .B2(G124), .ZN(new_n1238));
  AOI21_X1  g1038(.A(G33), .B1(new_n856), .B2(G159), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1237), .A2(new_n1238), .A3(new_n1239), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n224), .B1(new_n253), .B2(G41), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(G107), .A2(new_n842), .B1(new_n858), .B2(G283), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1242), .B1(new_n202), .B2(new_n860), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n848), .A2(new_n226), .ZN(new_n1244));
  NOR4_X1   g1044(.A1(new_n1243), .A2(G41), .A3(new_n389), .A4(new_n1244), .ZN(new_n1245));
  OAI22_X1  g1045(.A1(new_n864), .A2(new_n553), .B1(new_n855), .B2(new_n875), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1246), .B1(new_n660), .B2(new_n920), .ZN(new_n1247));
  OAI211_X1 g1047(.A(new_n1245), .B(new_n1247), .C1(new_n556), .C2(new_n851), .ZN(new_n1248));
  XNOR2_X1  g1048(.A(new_n1248), .B(KEYINPUT58), .ZN(new_n1249));
  AND3_X1   g1049(.A1(new_n1240), .A2(new_n1241), .A3(new_n1249), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n1232), .B(new_n894), .C1(new_n889), .C2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1251), .B1(new_n201), .B2(new_n927), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1252), .B1(new_n1229), .B2(new_n1014), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1231), .A2(new_n1253), .ZN(G375));
  NAND2_X1  g1054(.A1(new_n1199), .A2(new_n1190), .ZN(new_n1255));
  XOR2_X1   g1055(.A(new_n1035), .B(KEYINPUT122), .Z(new_n1256));
  NAND3_X1  g1056(.A1(new_n1192), .A2(new_n1255), .A3(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n347), .B1(new_n856), .B2(G58), .ZN(new_n1258));
  OAI221_X1 g1058(.A(new_n1258), .B1(new_n224), .B2(new_n848), .C1(new_n909), .C2(new_n841), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(G132), .A2(new_n865), .B1(new_n867), .B2(G159), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n907), .A2(new_n1163), .ZN(new_n1261));
  OAI211_X1 g1061(.A(new_n1260), .B(new_n1261), .C1(new_n1095), .C2(new_n862), .ZN(new_n1262));
  AOI211_X1 g1062(.A(new_n1259), .B(new_n1262), .C1(G128), .C2(new_n858), .ZN(new_n1263));
  OAI22_X1  g1063(.A1(new_n864), .A2(new_n844), .B1(new_n841), .B2(new_n922), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1264), .B1(G107), .B2(new_n920), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n867), .A2(G97), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(G116), .A2(new_n907), .B1(new_n858), .B2(G303), .ZN(new_n1267));
  AND4_X1   g1067(.A1(new_n1100), .A2(new_n1265), .A3(new_n1266), .A4(new_n1267), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n347), .B1(new_n855), .B2(new_n202), .ZN(new_n1269));
  XOR2_X1   g1069(.A(new_n1269), .B(KEYINPUT123), .Z(new_n1270));
  AOI21_X1  g1070(.A(new_n1263), .B1(new_n1268), .B2(new_n1270), .ZN(new_n1271));
  XNOR2_X1  g1071(.A(new_n1271), .B(KEYINPUT124), .ZN(new_n1272));
  OAI221_X1 g1072(.A(new_n894), .B1(new_n889), .B2(new_n1272), .C1(new_n1139), .C2(new_n929), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1273), .B1(new_n226), .B2(new_n927), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1274), .B1(new_n1188), .B2(new_n1014), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1257), .A2(new_n1275), .ZN(G381));
  NAND3_X1  g1076(.A1(new_n1051), .A2(new_n1072), .A3(new_n1134), .ZN(new_n1277));
  OR3_X1    g1077(.A1(new_n1277), .A2(G396), .A3(G393), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  NOR4_X1   g1079(.A1(G375), .A2(G384), .A3(G378), .A4(G381), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(G407));
  INV_X1    g1081(.A(new_n1197), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n778), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1175), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n761), .A2(G213), .ZN(new_n1285));
  XOR2_X1   g1085(.A(new_n1285), .B(KEYINPUT125), .Z(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1231), .A2(new_n1284), .A3(new_n1253), .A4(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(G407), .A2(G213), .A3(new_n1288), .ZN(G409));
  XOR2_X1   g1089(.A(G393), .B(G396), .Z(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1277), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1134), .B1(new_n1051), .B2(new_n1072), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1291), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1293), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1295), .A2(new_n1277), .A3(new_n1290), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1294), .A2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT60), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1255), .A2(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1199), .A2(KEYINPUT60), .A3(new_n1190), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1299), .A2(new_n777), .A3(new_n1192), .A4(new_n1300), .ZN(new_n1301));
  AOI21_X1  g1101(.A(G384), .B1(new_n1301), .B2(new_n1275), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1301), .A2(G384), .A3(new_n1275), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT63), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  OAI211_X1 g1107(.A(G378), .B(new_n1253), .C1(new_n1224), .C2(new_n1230), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1229), .A2(new_n1200), .A3(new_n1256), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1253), .A2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1310), .A2(new_n1284), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1287), .B1(new_n1308), .B2(new_n1311), .ZN(new_n1312));
  AOI21_X1  g1112(.A(KEYINPUT61), .B1(new_n1307), .B2(new_n1312), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1286), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1314));
  AND3_X1   g1114(.A1(new_n1301), .A2(G384), .A3(new_n1275), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1315), .A2(new_n1302), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n761), .A2(G213), .A3(G2897), .ZN(new_n1317));
  AOI22_X1  g1117(.A1(new_n1314), .A2(G2897), .B1(new_n1316), .B2(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1308), .A2(new_n1311), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1319), .A2(new_n1285), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1306), .B1(new_n1318), .B2(new_n1320), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1320), .A2(new_n1305), .ZN(new_n1322));
  OAI211_X1 g1122(.A(new_n1297), .B(new_n1313), .C1(new_n1321), .C2(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT61), .ZN(new_n1324));
  OAI211_X1 g1124(.A(G2897), .B(new_n1287), .C1(new_n1315), .C2(new_n1302), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1317), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1325), .B1(new_n1305), .B2(new_n1326), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1324), .B1(new_n1327), .B2(new_n1312), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT62), .ZN(new_n1329));
  NOR3_X1   g1129(.A1(new_n1315), .A2(new_n1302), .A3(new_n1329), .ZN(new_n1330));
  AND4_X1   g1130(.A1(KEYINPUT126), .A2(new_n1319), .A3(new_n1286), .A4(new_n1330), .ZN(new_n1331));
  AOI21_X1  g1131(.A(KEYINPUT126), .B1(new_n1312), .B2(new_n1330), .ZN(new_n1332));
  NOR2_X1   g1132(.A1(new_n1331), .A2(new_n1332), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1329), .B1(new_n1320), .B2(new_n1305), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1328), .B1(new_n1333), .B2(new_n1334), .ZN(new_n1335));
  OAI21_X1  g1135(.A(new_n1323), .B1(new_n1335), .B2(new_n1297), .ZN(G405));
  NAND2_X1  g1136(.A1(new_n1305), .A2(KEYINPUT127), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT127), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1316), .A2(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1337), .A2(new_n1339), .ZN(new_n1340));
  AOI21_X1  g1140(.A(G378), .B1(new_n1231), .B2(new_n1253), .ZN(new_n1341));
  INV_X1    g1141(.A(new_n1341), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1340), .A2(new_n1308), .A3(new_n1342), .ZN(new_n1343));
  INV_X1    g1143(.A(new_n1308), .ZN(new_n1344));
  OAI21_X1  g1144(.A(new_n1337), .B1(new_n1341), .B2(new_n1344), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1343), .A2(new_n1345), .ZN(new_n1346));
  AND2_X1   g1146(.A1(new_n1294), .A2(new_n1296), .ZN(new_n1347));
  XNOR2_X1  g1147(.A(new_n1346), .B(new_n1347), .ZN(G402));
endmodule


